magic
tech gf180mcuD
magscale 1 10
timestamp 1702341631
<< metal1 >>
rect 1344 46282 48608 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 48608 46282
rect 1344 46196 48608 46230
rect 19182 46114 19234 46126
rect 19182 46050 19234 46062
rect 22094 46114 22146 46126
rect 36990 46114 37042 46126
rect 25218 46062 25230 46114
rect 25282 46062 25294 46114
rect 22094 46050 22146 46062
rect 36990 46050 37042 46062
rect 44606 46114 44658 46126
rect 44606 46050 44658 46062
rect 16034 45950 16046 46002
rect 16098 45950 16110 46002
rect 30258 45950 30270 46002
rect 30322 45950 30334 46002
rect 35074 45950 35086 46002
rect 35138 45950 35150 46002
rect 40338 45950 40350 46002
rect 40402 45950 40414 46002
rect 46834 45950 46846 46002
rect 46898 45950 46910 46002
rect 47966 45890 48018 45902
rect 9650 45838 9662 45890
rect 9714 45838 9726 45890
rect 13122 45838 13134 45890
rect 13186 45838 13198 45890
rect 19730 45838 19742 45890
rect 19794 45838 19806 45890
rect 21074 45838 21086 45890
rect 21138 45838 21150 45890
rect 27122 45838 27134 45890
rect 27186 45838 27198 45890
rect 31154 45838 31166 45890
rect 31218 45838 31230 45890
rect 32162 45838 32174 45890
rect 32226 45838 32238 45890
rect 35970 45838 35982 45890
rect 36034 45838 36046 45890
rect 38882 45838 38894 45890
rect 38946 45838 38958 45890
rect 42354 45838 42366 45890
rect 42418 45838 42430 45890
rect 43922 45838 43934 45890
rect 43986 45838 43998 45890
rect 47966 45826 48018 45838
rect 3838 45778 3890 45790
rect 3838 45714 3890 45726
rect 5518 45778 5570 45790
rect 5518 45714 5570 45726
rect 6974 45778 7026 45790
rect 6974 45714 7026 45726
rect 8542 45778 8594 45790
rect 8542 45714 8594 45726
rect 9326 45778 9378 45790
rect 9326 45714 9378 45726
rect 10110 45778 10162 45790
rect 10110 45714 10162 45726
rect 11678 45778 11730 45790
rect 11678 45714 11730 45726
rect 12574 45778 12626 45790
rect 16942 45778 16994 45790
rect 13906 45726 13918 45778
rect 13970 45726 13982 45778
rect 12574 45714 12626 45726
rect 16942 45714 16994 45726
rect 27470 45778 27522 45790
rect 27470 45714 27522 45726
rect 28702 45778 28754 45790
rect 39230 45778 39282 45790
rect 32946 45726 32958 45778
rect 33010 45726 33022 45778
rect 28702 45714 28754 45726
rect 39230 45714 39282 45726
rect 42702 45778 42754 45790
rect 42702 45714 42754 45726
rect 46510 45778 46562 45790
rect 46510 45714 46562 45726
rect 7982 45666 8034 45678
rect 7982 45602 8034 45614
rect 9438 45666 9490 45678
rect 9438 45602 9490 45614
rect 10894 45666 10946 45678
rect 10894 45602 10946 45614
rect 11342 45666 11394 45678
rect 11342 45602 11394 45614
rect 39118 45666 39170 45678
rect 39118 45602 39170 45614
rect 42814 45666 42866 45678
rect 42814 45602 42866 45614
rect 42926 45666 42978 45678
rect 42926 45602 42978 45614
rect 46734 45666 46786 45678
rect 46734 45602 46786 45614
rect 47406 45666 47458 45678
rect 47406 45602 47458 45614
rect 1344 45498 48608 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 48608 45498
rect 1344 45412 48608 45446
rect 13022 45330 13074 45342
rect 13022 45266 13074 45278
rect 24446 45330 24498 45342
rect 24446 45266 24498 45278
rect 26686 45330 26738 45342
rect 26686 45266 26738 45278
rect 30942 45330 30994 45342
rect 30942 45266 30994 45278
rect 39678 45330 39730 45342
rect 39678 45266 39730 45278
rect 2942 45218 2994 45230
rect 8206 45218 8258 45230
rect 5618 45166 5630 45218
rect 5682 45166 5694 45218
rect 2942 45154 2994 45166
rect 8206 45154 8258 45166
rect 25454 45218 25506 45230
rect 25454 45154 25506 45166
rect 44830 45218 44882 45230
rect 47394 45166 47406 45218
rect 47458 45166 47470 45218
rect 44830 45154 44882 45166
rect 3278 45106 3330 45118
rect 3278 45042 3330 45054
rect 3390 45106 3442 45118
rect 12686 45106 12738 45118
rect 4946 45054 4958 45106
rect 5010 45054 5022 45106
rect 9538 45054 9550 45106
rect 9602 45054 9614 45106
rect 3390 45042 3442 45054
rect 12686 45042 12738 45054
rect 13022 45106 13074 45118
rect 13022 45042 13074 45054
rect 13246 45106 13298 45118
rect 17502 45106 17554 45118
rect 24334 45106 24386 45118
rect 14018 45054 14030 45106
rect 14082 45054 14094 45106
rect 17938 45054 17950 45106
rect 18002 45054 18014 45106
rect 21074 45054 21086 45106
rect 21138 45054 21150 45106
rect 13246 45042 13298 45054
rect 17502 45042 17554 45054
rect 24334 45042 24386 45054
rect 24670 45106 24722 45118
rect 24670 45042 24722 45054
rect 25566 45106 25618 45118
rect 32510 45106 32562 45118
rect 39902 45106 39954 45118
rect 44606 45106 44658 45118
rect 26338 45054 26350 45106
rect 26402 45054 26414 45106
rect 29922 45054 29934 45106
rect 29986 45054 29998 45106
rect 33170 45054 33182 45106
rect 33234 45054 33246 45106
rect 36418 45054 36430 45106
rect 36482 45054 36494 45106
rect 40226 45054 40238 45106
rect 40290 45054 40302 45106
rect 41010 45054 41022 45106
rect 41074 45054 41086 45106
rect 44146 45054 44158 45106
rect 44210 45054 44222 45106
rect 25566 45042 25618 45054
rect 32510 45042 32562 45054
rect 39902 45042 39954 45054
rect 44606 45042 44658 45054
rect 44942 45106 44994 45118
rect 48178 45054 48190 45106
rect 48242 45054 48254 45106
rect 44942 45042 44994 45054
rect 3054 44994 3106 45006
rect 8990 44994 9042 45006
rect 26126 44994 26178 45006
rect 30494 44994 30546 45006
rect 7746 44942 7758 44994
rect 7810 44942 7822 44994
rect 10322 44942 10334 44994
rect 10386 44942 10398 44994
rect 12450 44942 12462 44994
rect 12514 44942 12526 44994
rect 14690 44942 14702 44994
rect 14754 44942 14766 44994
rect 16818 44942 16830 44994
rect 16882 44942 16894 44994
rect 18610 44942 18622 44994
rect 18674 44942 18686 44994
rect 20738 44942 20750 44994
rect 20802 44942 20814 44994
rect 21858 44942 21870 44994
rect 21922 44942 21934 44994
rect 23986 44942 23998 44994
rect 24050 44942 24062 44994
rect 27122 44942 27134 44994
rect 27186 44942 27198 44994
rect 29250 44942 29262 44994
rect 29314 44942 29326 44994
rect 3054 44930 3106 44942
rect 8990 44930 9042 44942
rect 26126 44930 26178 44942
rect 30494 44930 30546 44942
rect 31390 44994 31442 45006
rect 31390 44930 31442 44942
rect 31950 44994 32002 45006
rect 39790 44994 39842 45006
rect 33954 44942 33966 44994
rect 34018 44942 34030 44994
rect 36082 44942 36094 44994
rect 36146 44942 36158 44994
rect 37202 44942 37214 44994
rect 37266 44942 37278 44994
rect 39330 44942 39342 44994
rect 39394 44942 39406 44994
rect 41682 44942 41694 44994
rect 41746 44942 41758 44994
rect 43810 44942 43822 44994
rect 43874 44942 43886 44994
rect 45266 44942 45278 44994
rect 45330 44942 45342 44994
rect 31950 44930 32002 44942
rect 39790 44930 39842 44942
rect 8094 44882 8146 44894
rect 8094 44818 8146 44830
rect 8430 44882 8482 44894
rect 8430 44818 8482 44830
rect 25454 44882 25506 44894
rect 25454 44818 25506 44830
rect 26014 44882 26066 44894
rect 44370 44830 44382 44882
rect 44434 44830 44446 44882
rect 26014 44818 26066 44830
rect 1344 44714 48608 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 48608 44714
rect 1344 44628 48608 44662
rect 15374 44546 15426 44558
rect 15374 44482 15426 44494
rect 21310 44546 21362 44558
rect 21310 44482 21362 44494
rect 33742 44546 33794 44558
rect 33742 44482 33794 44494
rect 37214 44546 37266 44558
rect 37214 44482 37266 44494
rect 45838 44546 45890 44558
rect 45838 44482 45890 44494
rect 6190 44434 6242 44446
rect 2594 44382 2606 44434
rect 2658 44382 2670 44434
rect 4722 44382 4734 44434
rect 4786 44382 4798 44434
rect 6190 44370 6242 44382
rect 9102 44434 9154 44446
rect 9102 44370 9154 44382
rect 10222 44434 10274 44446
rect 19618 44382 19630 44434
rect 19682 44382 19694 44434
rect 26002 44382 26014 44434
rect 26066 44382 26078 44434
rect 32386 44382 32398 44434
rect 32450 44382 32462 44434
rect 36306 44382 36318 44434
rect 36370 44382 36382 44434
rect 44258 44382 44270 44434
rect 44322 44382 44334 44434
rect 10222 44370 10274 44382
rect 9662 44322 9714 44334
rect 24558 44322 24610 44334
rect 26910 44322 26962 44334
rect 28366 44322 28418 44334
rect 40014 44322 40066 44334
rect 1922 44270 1934 44322
rect 1986 44270 1998 44322
rect 7746 44270 7758 44322
rect 7810 44270 7822 44322
rect 8642 44270 8654 44322
rect 8706 44270 8718 44322
rect 12226 44270 12238 44322
rect 12290 44270 12302 44322
rect 16034 44270 16046 44322
rect 16098 44270 16110 44322
rect 16818 44270 16830 44322
rect 16882 44270 16894 44322
rect 24210 44270 24222 44322
rect 24274 44270 24286 44322
rect 25442 44270 25454 44322
rect 25506 44270 25518 44322
rect 27122 44270 27134 44322
rect 27186 44270 27198 44322
rect 29586 44270 29598 44322
rect 29650 44270 29662 44322
rect 32722 44270 32734 44322
rect 32786 44270 32798 44322
rect 35970 44270 35982 44322
rect 36034 44270 36046 44322
rect 39106 44270 39118 44322
rect 39170 44270 39182 44322
rect 40338 44270 40350 44322
rect 40402 44270 40414 44322
rect 41346 44270 41358 44322
rect 41410 44270 41422 44322
rect 45042 44270 45054 44322
rect 45106 44270 45118 44322
rect 9662 44258 9714 44270
rect 24558 44258 24610 44270
rect 26910 44258 26962 44270
rect 28366 44258 28418 44270
rect 40014 44258 40066 44270
rect 5742 44210 5794 44222
rect 5742 44146 5794 44158
rect 5854 44210 5906 44222
rect 5854 44146 5906 44158
rect 6302 44210 6354 44222
rect 9550 44210 9602 44222
rect 7410 44158 7422 44210
rect 7474 44158 7486 44210
rect 6302 44146 6354 44158
rect 9550 44146 9602 44158
rect 10334 44210 10386 44222
rect 10334 44146 10386 44158
rect 10670 44210 10722 44222
rect 21422 44210 21474 44222
rect 10882 44158 10894 44210
rect 10946 44158 10958 44210
rect 12562 44158 12574 44210
rect 12626 44158 12638 44210
rect 17490 44158 17502 44210
rect 17554 44158 17566 44210
rect 10670 44146 10722 44158
rect 21422 44146 21474 44158
rect 23326 44210 23378 44222
rect 23326 44146 23378 44158
rect 27806 44210 27858 44222
rect 27806 44146 27858 44158
rect 28254 44210 28306 44222
rect 39902 44210 39954 44222
rect 47742 44210 47794 44222
rect 30258 44158 30270 44210
rect 30322 44158 30334 44210
rect 42130 44158 42142 44210
rect 42194 44158 42206 44210
rect 28254 44146 28306 44158
rect 39902 44146 39954 44158
rect 47742 44146 47794 44158
rect 48078 44210 48130 44222
rect 48078 44146 48130 44158
rect 5518 44098 5570 44110
rect 5518 44034 5570 44046
rect 9326 44098 9378 44110
rect 9326 44034 9378 44046
rect 10110 44098 10162 44110
rect 10110 44034 10162 44046
rect 20078 44098 20130 44110
rect 20078 44034 20130 44046
rect 20526 44098 20578 44110
rect 20526 44034 20578 44046
rect 21870 44098 21922 44110
rect 21870 44034 21922 44046
rect 22318 44098 22370 44110
rect 22318 44034 22370 44046
rect 22990 44098 23042 44110
rect 22990 44034 23042 44046
rect 26462 44098 26514 44110
rect 26462 44034 26514 44046
rect 28030 44098 28082 44110
rect 28030 44034 28082 44046
rect 1344 43930 48608 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 48608 43930
rect 1344 43844 48608 43878
rect 3278 43762 3330 43774
rect 3278 43698 3330 43710
rect 3390 43762 3442 43774
rect 3390 43698 3442 43710
rect 6526 43762 6578 43774
rect 6526 43698 6578 43710
rect 7310 43762 7362 43774
rect 12574 43762 12626 43774
rect 7746 43710 7758 43762
rect 7810 43710 7822 43762
rect 9986 43710 9998 43762
rect 10050 43710 10062 43762
rect 7310 43698 7362 43710
rect 12574 43698 12626 43710
rect 12798 43762 12850 43774
rect 12798 43698 12850 43710
rect 13022 43762 13074 43774
rect 13022 43698 13074 43710
rect 13134 43762 13186 43774
rect 13134 43698 13186 43710
rect 14814 43762 14866 43774
rect 14814 43698 14866 43710
rect 24334 43762 24386 43774
rect 24334 43698 24386 43710
rect 24558 43762 24610 43774
rect 24558 43698 24610 43710
rect 25230 43762 25282 43774
rect 25230 43698 25282 43710
rect 27806 43762 27858 43774
rect 44606 43762 44658 43774
rect 34066 43710 34078 43762
rect 34130 43710 34142 43762
rect 27806 43698 27858 43710
rect 44606 43698 44658 43710
rect 4846 43650 4898 43662
rect 4846 43586 4898 43598
rect 7198 43650 7250 43662
rect 12462 43650 12514 43662
rect 8642 43598 8654 43650
rect 8706 43598 8718 43650
rect 7198 43586 7250 43598
rect 12462 43586 12514 43598
rect 13918 43650 13970 43662
rect 13918 43586 13970 43598
rect 14030 43650 14082 43662
rect 14030 43586 14082 43598
rect 14702 43650 14754 43662
rect 14702 43586 14754 43598
rect 15374 43650 15426 43662
rect 15374 43586 15426 43598
rect 20974 43650 21026 43662
rect 20974 43586 21026 43598
rect 22766 43650 22818 43662
rect 22766 43586 22818 43598
rect 24222 43650 24274 43662
rect 24222 43586 24274 43598
rect 25118 43650 25170 43662
rect 25118 43586 25170 43598
rect 25678 43650 25730 43662
rect 25678 43586 25730 43598
rect 26574 43650 26626 43662
rect 26574 43586 26626 43598
rect 26686 43650 26738 43662
rect 26686 43586 26738 43598
rect 27470 43650 27522 43662
rect 27470 43586 27522 43598
rect 27918 43650 27970 43662
rect 34750 43650 34802 43662
rect 30930 43598 30942 43650
rect 30994 43598 31006 43650
rect 33394 43598 33406 43650
rect 33458 43598 33470 43650
rect 27918 43586 27970 43598
rect 34750 43586 34802 43598
rect 34862 43650 34914 43662
rect 34862 43586 34914 43598
rect 38334 43650 38386 43662
rect 38334 43586 38386 43598
rect 38782 43650 38834 43662
rect 38782 43586 38834 43598
rect 44830 43650 44882 43662
rect 44830 43586 44882 43598
rect 3502 43538 3554 43550
rect 6078 43538 6130 43550
rect 3826 43486 3838 43538
rect 3890 43486 3902 43538
rect 5394 43486 5406 43538
rect 5458 43486 5470 43538
rect 3502 43474 3554 43486
rect 6078 43474 6130 43486
rect 6750 43538 6802 43550
rect 10334 43538 10386 43550
rect 7858 43486 7870 43538
rect 7922 43486 7934 43538
rect 8754 43486 8766 43538
rect 8818 43486 8830 43538
rect 6750 43474 6802 43486
rect 10334 43474 10386 43486
rect 13246 43538 13298 43550
rect 15262 43538 15314 43550
rect 13570 43486 13582 43538
rect 13634 43486 13646 43538
rect 13246 43474 13298 43486
rect 15262 43474 15314 43486
rect 15486 43538 15538 43550
rect 15486 43474 15538 43486
rect 15710 43538 15762 43550
rect 15710 43474 15762 43486
rect 16158 43538 16210 43550
rect 16158 43474 16210 43486
rect 16382 43538 16434 43550
rect 16382 43474 16434 43486
rect 16830 43538 16882 43550
rect 22654 43538 22706 43550
rect 17490 43486 17502 43538
rect 17554 43486 17566 43538
rect 16830 43474 16882 43486
rect 22654 43474 22706 43486
rect 22990 43538 23042 43550
rect 26462 43538 26514 43550
rect 28030 43538 28082 43550
rect 23762 43486 23774 43538
rect 23826 43486 23838 43538
rect 25442 43486 25454 43538
rect 25506 43486 25518 43538
rect 27010 43486 27022 43538
rect 27074 43486 27086 43538
rect 22990 43474 23042 43486
rect 26462 43474 26514 43486
rect 28030 43474 28082 43486
rect 28478 43538 28530 43550
rect 29710 43538 29762 43550
rect 31614 43538 31666 43550
rect 38558 43538 38610 43550
rect 44942 43538 44994 43550
rect 29026 43486 29038 43538
rect 29090 43486 29102 43538
rect 30146 43486 30158 43538
rect 30210 43486 30222 43538
rect 31154 43486 31166 43538
rect 31218 43486 31230 43538
rect 32050 43486 32062 43538
rect 32114 43486 32126 43538
rect 33282 43486 33294 43538
rect 33346 43486 33358 43538
rect 33954 43486 33966 43538
rect 34018 43486 34030 43538
rect 37538 43486 37550 43538
rect 37602 43486 37614 43538
rect 38098 43486 38110 43538
rect 38162 43486 38174 43538
rect 39106 43486 39118 43538
rect 39170 43486 39182 43538
rect 43026 43486 43038 43538
rect 43090 43486 43102 43538
rect 43922 43486 43934 43538
rect 43986 43486 43998 43538
rect 48178 43486 48190 43538
rect 48242 43486 48254 43538
rect 28478 43474 28530 43486
rect 29710 43474 29762 43486
rect 31614 43474 31666 43486
rect 38558 43474 38610 43486
rect 44942 43474 44994 43486
rect 1822 43426 1874 43438
rect 1822 43362 1874 43374
rect 4510 43426 4562 43438
rect 6638 43426 6690 43438
rect 5730 43374 5742 43426
rect 5794 43374 5806 43426
rect 4510 43362 4562 43374
rect 6638 43362 6690 43374
rect 9662 43426 9714 43438
rect 9662 43362 9714 43374
rect 10782 43426 10834 43438
rect 10782 43362 10834 43374
rect 11342 43426 11394 43438
rect 11342 43362 11394 43374
rect 11790 43426 11842 43438
rect 11790 43362 11842 43374
rect 12238 43426 12290 43438
rect 12238 43362 12290 43374
rect 14926 43426 14978 43438
rect 14926 43362 14978 43374
rect 16270 43426 16322 43438
rect 21982 43426 22034 43438
rect 18162 43374 18174 43426
rect 18226 43374 18238 43426
rect 20290 43374 20302 43426
rect 20354 43374 20366 43426
rect 20850 43374 20862 43426
rect 20914 43374 20926 43426
rect 16270 43362 16322 43374
rect 21982 43362 22034 43374
rect 22430 43426 22482 43438
rect 22430 43362 22482 43374
rect 23438 43426 23490 43438
rect 26126 43426 26178 43438
rect 32510 43426 32562 43438
rect 24322 43374 24334 43426
rect 24386 43374 24398 43426
rect 29362 43374 29374 43426
rect 29426 43374 29438 43426
rect 31042 43374 31054 43426
rect 31106 43374 31118 43426
rect 23438 43362 23490 43374
rect 26126 43362 26178 43374
rect 32510 43362 32562 43374
rect 35422 43426 35474 43438
rect 35422 43362 35474 43374
rect 38446 43426 38498 43438
rect 38446 43362 38498 43374
rect 40014 43426 40066 43438
rect 41134 43426 41186 43438
rect 40226 43374 40238 43426
rect 40290 43374 40302 43426
rect 40014 43362 40066 43374
rect 41134 43362 41186 43374
rect 44382 43426 44434 43438
rect 45266 43374 45278 43426
rect 45330 43374 45342 43426
rect 47394 43374 47406 43426
rect 47458 43374 47470 43426
rect 44382 43362 44434 43374
rect 14030 43314 14082 43326
rect 11330 43262 11342 43314
rect 11394 43311 11406 43314
rect 12226 43311 12238 43314
rect 11394 43265 12238 43311
rect 11394 43262 11406 43265
rect 12226 43262 12238 43265
rect 12290 43262 12302 43314
rect 14030 43250 14082 43262
rect 21198 43314 21250 43326
rect 21198 43250 21250 43262
rect 34750 43314 34802 43326
rect 34750 43250 34802 43262
rect 39118 43314 39170 43326
rect 39118 43250 39170 43262
rect 39454 43314 39506 43326
rect 39454 43250 39506 43262
rect 1344 43146 48608 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 48608 43146
rect 1344 43060 48608 43094
rect 6302 42978 6354 42990
rect 6302 42914 6354 42926
rect 18958 42978 19010 42990
rect 18958 42914 19010 42926
rect 22318 42978 22370 42990
rect 22318 42914 22370 42926
rect 37102 42978 37154 42990
rect 37102 42914 37154 42926
rect 39342 42978 39394 42990
rect 39342 42914 39394 42926
rect 45838 42978 45890 42990
rect 45838 42914 45890 42926
rect 3726 42866 3778 42878
rect 23662 42866 23714 42878
rect 3154 42814 3166 42866
rect 3218 42814 3230 42866
rect 4722 42814 4734 42866
rect 4786 42814 4798 42866
rect 7858 42814 7870 42866
rect 7922 42814 7934 42866
rect 9538 42814 9550 42866
rect 9602 42814 9614 42866
rect 14130 42814 14142 42866
rect 14194 42814 14206 42866
rect 22866 42814 22878 42866
rect 22930 42814 22942 42866
rect 3726 42802 3778 42814
rect 23662 42802 23714 42814
rect 29262 42866 29314 42878
rect 30942 42866 30994 42878
rect 36206 42866 36258 42878
rect 43262 42866 43314 42878
rect 29474 42814 29486 42866
rect 29538 42814 29550 42866
rect 30034 42814 30046 42866
rect 30098 42814 30110 42866
rect 34066 42814 34078 42866
rect 34130 42814 34142 42866
rect 35298 42814 35310 42866
rect 35362 42814 35374 42866
rect 39666 42814 39678 42866
rect 39730 42814 39742 42866
rect 29262 42802 29314 42814
rect 30942 42802 30994 42814
rect 36206 42802 36258 42814
rect 43262 42802 43314 42814
rect 43710 42866 43762 42878
rect 43710 42802 43762 42814
rect 2270 42754 2322 42766
rect 5630 42754 5682 42766
rect 1810 42702 1822 42754
rect 1874 42702 1886 42754
rect 4050 42702 4062 42754
rect 4114 42702 4126 42754
rect 4834 42702 4846 42754
rect 4898 42702 4910 42754
rect 2270 42690 2322 42702
rect 5630 42690 5682 42702
rect 5966 42754 6018 42766
rect 5966 42690 6018 42702
rect 6974 42754 7026 42766
rect 6974 42690 7026 42702
rect 13694 42754 13746 42766
rect 21422 42754 21474 42766
rect 14578 42702 14590 42754
rect 14642 42702 14654 42754
rect 15698 42702 15710 42754
rect 15762 42702 15774 42754
rect 17938 42702 17950 42754
rect 18002 42702 18014 42754
rect 13694 42690 13746 42702
rect 21422 42690 21474 42702
rect 21982 42754 22034 42766
rect 26462 42754 26514 42766
rect 22978 42702 22990 42754
rect 23042 42702 23054 42754
rect 21982 42690 22034 42702
rect 26462 42690 26514 42702
rect 27694 42754 27746 42766
rect 27694 42690 27746 42702
rect 27918 42754 27970 42766
rect 27918 42690 27970 42702
rect 28142 42754 28194 42766
rect 31838 42754 31890 42766
rect 43934 42754 43986 42766
rect 30258 42702 30270 42754
rect 30322 42702 30334 42754
rect 31266 42702 31278 42754
rect 31330 42702 31342 42754
rect 33730 42702 33742 42754
rect 33794 42702 33806 42754
rect 34178 42702 34190 42754
rect 34242 42702 34254 42754
rect 35522 42702 35534 42754
rect 35586 42702 35598 42754
rect 38098 42702 38110 42754
rect 38162 42702 38174 42754
rect 38322 42702 38334 42754
rect 38386 42702 38398 42754
rect 42466 42702 42478 42754
rect 42530 42702 42542 42754
rect 45042 42702 45054 42754
rect 45106 42702 45118 42754
rect 28142 42690 28194 42702
rect 31838 42690 31890 42702
rect 43934 42690 43986 42702
rect 2830 42642 2882 42654
rect 2830 42578 2882 42590
rect 3054 42642 3106 42654
rect 3054 42578 3106 42590
rect 5742 42642 5794 42654
rect 5742 42578 5794 42590
rect 6414 42642 6466 42654
rect 6414 42578 6466 42590
rect 7534 42642 7586 42654
rect 7534 42578 7586 42590
rect 7758 42642 7810 42654
rect 7758 42578 7810 42590
rect 8654 42642 8706 42654
rect 8654 42578 8706 42590
rect 8878 42642 8930 42654
rect 11678 42642 11730 42654
rect 9986 42590 9998 42642
rect 10050 42590 10062 42642
rect 11442 42590 11454 42642
rect 11506 42590 11518 42642
rect 8878 42578 8930 42590
rect 11678 42578 11730 42590
rect 12014 42642 12066 42654
rect 17390 42642 17442 42654
rect 12898 42590 12910 42642
rect 12962 42590 12974 42642
rect 16146 42590 16158 42642
rect 16210 42590 16222 42642
rect 12014 42578 12066 42590
rect 17390 42578 17442 42590
rect 21758 42642 21810 42654
rect 21758 42578 21810 42590
rect 24334 42642 24386 42654
rect 24334 42578 24386 42590
rect 25342 42642 25394 42654
rect 25342 42578 25394 42590
rect 25790 42642 25842 42654
rect 25790 42578 25842 42590
rect 26126 42642 26178 42654
rect 26126 42578 26178 42590
rect 26798 42642 26850 42654
rect 26798 42578 26850 42590
rect 37102 42642 37154 42654
rect 37102 42578 37154 42590
rect 37214 42642 37266 42654
rect 37214 42578 37266 42590
rect 38558 42642 38610 42654
rect 38558 42578 38610 42590
rect 39006 42642 39058 42654
rect 43150 42642 43202 42654
rect 41794 42590 41806 42642
rect 41858 42590 41870 42642
rect 39006 42578 39058 42590
rect 43150 42578 43202 42590
rect 43374 42642 43426 42654
rect 43374 42578 43426 42590
rect 48190 42642 48242 42654
rect 48190 42578 48242 42590
rect 6302 42530 6354 42542
rect 6302 42466 6354 42478
rect 7086 42530 7138 42542
rect 7086 42466 7138 42478
rect 7310 42530 7362 42542
rect 7310 42466 7362 42478
rect 8766 42530 8818 42542
rect 8766 42466 8818 42478
rect 12126 42530 12178 42542
rect 12126 42466 12178 42478
rect 12350 42530 12402 42542
rect 12350 42466 12402 42478
rect 12574 42530 12626 42542
rect 12574 42466 12626 42478
rect 13358 42530 13410 42542
rect 13358 42466 13410 42478
rect 13582 42530 13634 42542
rect 13582 42466 13634 42478
rect 16942 42530 16994 42542
rect 16942 42466 16994 42478
rect 17502 42530 17554 42542
rect 17502 42466 17554 42478
rect 17726 42530 17778 42542
rect 17726 42466 17778 42478
rect 21310 42530 21362 42542
rect 21310 42466 21362 42478
rect 24446 42530 24498 42542
rect 24446 42466 24498 42478
rect 24670 42530 24722 42542
rect 24670 42466 24722 42478
rect 25230 42530 25282 42542
rect 25230 42466 25282 42478
rect 26238 42530 26290 42542
rect 26238 42466 26290 42478
rect 26686 42530 26738 42542
rect 26686 42466 26738 42478
rect 26910 42530 26962 42542
rect 26910 42466 26962 42478
rect 27134 42530 27186 42542
rect 27134 42466 27186 42478
rect 27918 42530 27970 42542
rect 27918 42466 27970 42478
rect 29486 42530 29538 42542
rect 29486 42466 29538 42478
rect 39230 42530 39282 42542
rect 47854 42530 47906 42542
rect 44258 42478 44270 42530
rect 44322 42478 44334 42530
rect 39230 42466 39282 42478
rect 47854 42466 47906 42478
rect 1344 42362 48608 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 48608 42362
rect 1344 42276 48608 42310
rect 22318 42194 22370 42206
rect 12114 42142 12126 42194
rect 12178 42142 12190 42194
rect 22318 42130 22370 42142
rect 22542 42194 22594 42206
rect 22542 42130 22594 42142
rect 23102 42194 23154 42206
rect 23102 42130 23154 42142
rect 23326 42194 23378 42206
rect 23326 42130 23378 42142
rect 26462 42194 26514 42206
rect 39778 42142 39790 42194
rect 39842 42142 39854 42194
rect 26462 42130 26514 42142
rect 21198 42082 21250 42094
rect 21870 42082 21922 42094
rect 19618 42030 19630 42082
rect 19682 42030 19694 42082
rect 21522 42030 21534 42082
rect 21586 42030 21598 42082
rect 21198 42018 21250 42030
rect 21870 42018 21922 42030
rect 22206 42082 22258 42094
rect 22206 42018 22258 42030
rect 25230 42082 25282 42094
rect 25230 42018 25282 42030
rect 25342 42082 25394 42094
rect 25342 42018 25394 42030
rect 26126 42082 26178 42094
rect 26126 42018 26178 42030
rect 26238 42082 26290 42094
rect 36430 42082 36482 42094
rect 34626 42030 34638 42082
rect 34690 42030 34702 42082
rect 26238 42018 26290 42030
rect 36430 42018 36482 42030
rect 36990 42082 37042 42094
rect 36990 42018 37042 42030
rect 37662 42082 37714 42094
rect 37662 42018 37714 42030
rect 37998 42082 38050 42094
rect 37998 42018 38050 42030
rect 38222 42082 38274 42094
rect 38882 42030 38894 42082
rect 38946 42030 38958 42082
rect 41458 42030 41470 42082
rect 41522 42030 41534 42082
rect 43362 42030 43374 42082
rect 43426 42030 43438 42082
rect 38222 42018 38274 42030
rect 8318 41970 8370 41982
rect 17950 41970 18002 41982
rect 4610 41918 4622 41970
rect 4674 41918 4686 41970
rect 4946 41918 4958 41970
rect 5010 41918 5022 41970
rect 5730 41918 5742 41970
rect 5794 41918 5806 41970
rect 9426 41918 9438 41970
rect 9490 41918 9502 41970
rect 10210 41918 10222 41970
rect 10274 41918 10286 41970
rect 13122 41918 13134 41970
rect 13186 41918 13198 41970
rect 16818 41918 16830 41970
rect 16882 41918 16894 41970
rect 8318 41906 8370 41918
rect 17950 41906 18002 41918
rect 18398 41970 18450 41982
rect 18398 41906 18450 41918
rect 18622 41970 18674 41982
rect 24670 41970 24722 41982
rect 20514 41918 20526 41970
rect 20578 41918 20590 41970
rect 22754 41918 22766 41970
rect 22818 41918 22830 41970
rect 24210 41918 24222 41970
rect 24274 41918 24286 41970
rect 18622 41906 18674 41918
rect 24670 41906 24722 41918
rect 25566 41970 25618 41982
rect 30046 41970 30098 41982
rect 32398 41970 32450 41982
rect 29474 41918 29486 41970
rect 29538 41918 29550 41970
rect 30706 41918 30718 41970
rect 30770 41918 30782 41970
rect 31938 41918 31950 41970
rect 32002 41918 32014 41970
rect 25566 41906 25618 41918
rect 30046 41906 30098 41918
rect 32398 41906 32450 41918
rect 32510 41970 32562 41982
rect 32510 41906 32562 41918
rect 33070 41970 33122 41982
rect 36766 41970 36818 41982
rect 37774 41970 37826 41982
rect 41134 41970 41186 41982
rect 43822 41970 43874 41982
rect 35858 41918 35870 41970
rect 35922 41918 35934 41970
rect 37314 41918 37326 41970
rect 37378 41918 37390 41970
rect 38770 41918 38782 41970
rect 38834 41918 38846 41970
rect 39666 41918 39678 41970
rect 39730 41918 39742 41970
rect 42130 41918 42142 41970
rect 42194 41918 42206 41970
rect 42690 41918 42702 41970
rect 42754 41918 42766 41970
rect 42914 41918 42926 41970
rect 42978 41918 42990 41970
rect 33070 41906 33122 41918
rect 36766 41906 36818 41918
rect 37774 41906 37826 41918
rect 41134 41906 41186 41918
rect 43822 41906 43874 41918
rect 44830 41970 44882 41982
rect 44830 41906 44882 41918
rect 44942 41970 44994 41982
rect 47394 41918 47406 41970
rect 47458 41918 47470 41970
rect 48066 41918 48078 41970
rect 48130 41918 48142 41970
rect 44942 41906 44994 41918
rect 11566 41858 11618 41870
rect 17502 41858 17554 41870
rect 1698 41806 1710 41858
rect 1762 41806 1774 41858
rect 3826 41806 3838 41858
rect 3890 41806 3902 41858
rect 7858 41806 7870 41858
rect 7922 41806 7934 41858
rect 9762 41806 9774 41858
rect 9826 41806 9838 41858
rect 10098 41806 10110 41858
rect 10162 41806 10174 41858
rect 12674 41806 12686 41858
rect 12738 41806 12750 41858
rect 13906 41806 13918 41858
rect 13970 41806 13982 41858
rect 16034 41806 16046 41858
rect 16098 41806 16110 41858
rect 11566 41794 11618 41806
rect 17502 41794 17554 41806
rect 18174 41858 18226 41870
rect 23214 41858 23266 41870
rect 31166 41858 31218 41870
rect 34414 41858 34466 41870
rect 19058 41806 19070 41858
rect 19122 41806 19134 41858
rect 23762 41806 23774 41858
rect 23826 41806 23838 41858
rect 26674 41806 26686 41858
rect 26738 41806 26750 41858
rect 28802 41806 28814 41858
rect 28866 41806 28878 41858
rect 30594 41806 30606 41858
rect 30658 41806 30670 41858
rect 33506 41806 33518 41858
rect 33570 41806 33582 41858
rect 18174 41794 18226 41806
rect 23214 41794 23266 41806
rect 31166 41794 31218 41806
rect 34414 41794 34466 41806
rect 36878 41858 36930 41870
rect 36878 41794 36930 41806
rect 40238 41858 40290 41870
rect 41794 41806 41806 41858
rect 41858 41806 41870 41858
rect 45266 41806 45278 41858
rect 45330 41806 45342 41858
rect 40238 41794 40290 41806
rect 11790 41746 11842 41758
rect 40350 41746 40402 41758
rect 13458 41694 13470 41746
rect 13522 41694 13534 41746
rect 11790 41682 11842 41694
rect 40350 41682 40402 41694
rect 44046 41746 44098 41758
rect 44370 41694 44382 41746
rect 44434 41694 44446 41746
rect 44046 41682 44098 41694
rect 1344 41578 48608 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 48608 41578
rect 1344 41492 48608 41526
rect 16046 41410 16098 41422
rect 16046 41346 16098 41358
rect 19070 41410 19122 41422
rect 19070 41346 19122 41358
rect 19406 41410 19458 41422
rect 30158 41410 30210 41422
rect 31502 41410 31554 41422
rect 22082 41358 22094 41410
rect 22146 41407 22158 41410
rect 22866 41407 22878 41410
rect 22146 41361 22878 41407
rect 22146 41358 22158 41361
rect 22866 41358 22878 41361
rect 22930 41407 22942 41410
rect 23314 41407 23326 41410
rect 22930 41361 23326 41407
rect 22930 41358 22942 41361
rect 23314 41358 23326 41361
rect 23378 41358 23390 41410
rect 30482 41358 30494 41410
rect 30546 41358 30558 41410
rect 19406 41346 19458 41358
rect 30158 41346 30210 41358
rect 31502 41346 31554 41358
rect 32846 41410 32898 41422
rect 32846 41346 32898 41358
rect 33182 41410 33234 41422
rect 44146 41358 44158 41410
rect 44210 41358 44222 41410
rect 47058 41358 47070 41410
rect 47122 41358 47134 41410
rect 33182 41346 33234 41358
rect 8878 41298 8930 41310
rect 4610 41246 4622 41298
rect 4674 41246 4686 41298
rect 8878 41234 8930 41246
rect 10670 41298 10722 41310
rect 10670 41234 10722 41246
rect 14590 41298 14642 41310
rect 14590 41234 14642 41246
rect 15934 41298 15986 41310
rect 15934 41234 15986 41246
rect 21422 41298 21474 41310
rect 21422 41234 21474 41246
rect 22878 41298 22930 41310
rect 22878 41234 22930 41246
rect 23326 41298 23378 41310
rect 27134 41298 27186 41310
rect 26226 41246 26238 41298
rect 26290 41246 26302 41298
rect 23326 41234 23378 41246
rect 27134 41234 27186 41246
rect 27918 41298 27970 41310
rect 27918 41234 27970 41246
rect 28590 41298 28642 41310
rect 28590 41234 28642 41246
rect 29934 41298 29986 41310
rect 37662 41298 37714 41310
rect 36418 41246 36430 41298
rect 36482 41246 36494 41298
rect 29934 41234 29986 41246
rect 37662 41234 37714 41246
rect 38334 41298 38386 41310
rect 38334 41234 38386 41246
rect 38446 41298 38498 41310
rect 38446 41234 38498 41246
rect 11342 41186 11394 41198
rect 2706 41134 2718 41186
rect 2770 41134 2782 41186
rect 4722 41134 4734 41186
rect 4786 41134 4798 41186
rect 7522 41134 7534 41186
rect 7586 41134 7598 41186
rect 8306 41134 8318 41186
rect 8370 41134 8382 41186
rect 11106 41134 11118 41186
rect 11170 41134 11182 41186
rect 11342 41122 11394 41134
rect 12462 41186 12514 41198
rect 25118 41186 25170 41198
rect 31838 41186 31890 41198
rect 13458 41134 13470 41186
rect 13522 41134 13534 41186
rect 21858 41134 21870 41186
rect 21922 41134 21934 41186
rect 26674 41134 26686 41186
rect 26738 41134 26750 41186
rect 12462 41122 12514 41134
rect 25118 41122 25170 41134
rect 31838 41122 31890 41134
rect 32174 41186 32226 41198
rect 37438 41186 37490 41198
rect 33618 41134 33630 41186
rect 33682 41134 33694 41186
rect 32174 41122 32226 41134
rect 37438 41122 37490 41134
rect 37550 41186 37602 41198
rect 40686 41186 40738 41198
rect 42814 41186 42866 41198
rect 38658 41134 38670 41186
rect 38722 41134 38734 41186
rect 39666 41134 39678 41186
rect 39730 41134 39742 41186
rect 39890 41134 39902 41186
rect 39954 41134 39966 41186
rect 42466 41134 42478 41186
rect 42530 41134 42542 41186
rect 43474 41134 43486 41186
rect 43538 41134 43550 41186
rect 45602 41134 45614 41186
rect 45666 41134 45678 41186
rect 37550 41122 37602 41134
rect 40686 41122 40738 41134
rect 42814 41122 42866 41134
rect 4062 41074 4114 41086
rect 2258 41022 2270 41074
rect 2322 41022 2334 41074
rect 3826 41022 3838 41074
rect 3890 41022 3902 41074
rect 4062 41010 4114 41022
rect 4398 41074 4450 41086
rect 11678 41074 11730 41086
rect 19182 41074 19234 41086
rect 7186 41022 7198 41074
rect 7250 41022 7262 41074
rect 12786 41022 12798 41074
rect 12850 41022 12862 41074
rect 13682 41022 13694 41074
rect 13746 41022 13758 41074
rect 4398 41010 4450 41022
rect 11678 41010 11730 41022
rect 19182 41010 19234 41022
rect 23886 41074 23938 41086
rect 24782 41074 24834 41086
rect 24098 41022 24110 41074
rect 24162 41022 24174 41074
rect 23886 41010 23938 41022
rect 24782 41010 24834 41022
rect 27470 41074 27522 41086
rect 27470 41010 27522 41022
rect 27694 41074 27746 41086
rect 27694 41010 27746 41022
rect 28030 41074 28082 41086
rect 28030 41010 28082 41022
rect 31166 41074 31218 41086
rect 31166 41010 31218 41022
rect 31950 41074 32002 41086
rect 31950 41010 32002 41022
rect 33070 41074 33122 41086
rect 37998 41074 38050 41086
rect 44942 41074 44994 41086
rect 34290 41022 34302 41074
rect 34354 41022 34366 41074
rect 39106 41022 39118 41074
rect 39170 41022 39182 41074
rect 41122 41022 41134 41074
rect 41186 41022 41198 41074
rect 33070 41010 33122 41022
rect 37998 41010 38050 41022
rect 44942 41010 44994 41022
rect 5854 40962 5906 40974
rect 5854 40898 5906 40910
rect 9326 40962 9378 40974
rect 9326 40898 9378 40910
rect 9774 40962 9826 40974
rect 10558 40962 10610 40974
rect 10098 40910 10110 40962
rect 10162 40910 10174 40962
rect 9774 40898 9826 40910
rect 10558 40898 10610 40910
rect 10782 40962 10834 40974
rect 10782 40898 10834 40910
rect 11566 40962 11618 40974
rect 11566 40898 11618 40910
rect 12238 40962 12290 40974
rect 15486 40962 15538 40974
rect 14018 40910 14030 40962
rect 14082 40910 14094 40962
rect 12238 40898 12290 40910
rect 15486 40898 15538 40910
rect 15822 40962 15874 40974
rect 15822 40898 15874 40910
rect 18286 40962 18338 40974
rect 18286 40898 18338 40910
rect 20526 40962 20578 40974
rect 20526 40898 20578 40910
rect 21310 40962 21362 40974
rect 21310 40898 21362 40910
rect 21534 40962 21586 40974
rect 21534 40898 21586 40910
rect 22318 40962 22370 40974
rect 22318 40898 22370 40910
rect 24446 40962 24498 40974
rect 24446 40898 24498 40910
rect 24894 40962 24946 40974
rect 24894 40898 24946 40910
rect 25790 40962 25842 40974
rect 25790 40898 25842 40910
rect 29598 40962 29650 40974
rect 29598 40898 29650 40910
rect 31390 40962 31442 40974
rect 31390 40898 31442 40910
rect 32510 40962 32562 40974
rect 32510 40898 32562 40910
rect 37774 40962 37826 40974
rect 41470 40962 41522 40974
rect 40786 40910 40798 40962
rect 40850 40910 40862 40962
rect 45266 40910 45278 40962
rect 45330 40910 45342 40962
rect 37774 40898 37826 40910
rect 41470 40898 41522 40910
rect 1344 40794 48608 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 48608 40794
rect 1344 40708 48608 40742
rect 2494 40626 2546 40638
rect 2494 40562 2546 40574
rect 3278 40626 3330 40638
rect 5070 40626 5122 40638
rect 11118 40626 11170 40638
rect 4050 40574 4062 40626
rect 4114 40574 4126 40626
rect 7970 40574 7982 40626
rect 8034 40574 8046 40626
rect 10098 40574 10110 40626
rect 10162 40574 10174 40626
rect 3278 40562 3330 40574
rect 5070 40562 5122 40574
rect 11118 40562 11170 40574
rect 11678 40626 11730 40638
rect 11678 40562 11730 40574
rect 16942 40626 16994 40638
rect 16942 40562 16994 40574
rect 17726 40626 17778 40638
rect 25342 40626 25394 40638
rect 21746 40574 21758 40626
rect 21810 40574 21822 40626
rect 17726 40562 17778 40574
rect 25342 40562 25394 40574
rect 25566 40626 25618 40638
rect 27022 40626 27074 40638
rect 26226 40574 26238 40626
rect 26290 40574 26302 40626
rect 25566 40562 25618 40574
rect 27022 40562 27074 40574
rect 27134 40626 27186 40638
rect 27134 40562 27186 40574
rect 27470 40626 27522 40638
rect 27470 40562 27522 40574
rect 35982 40626 36034 40638
rect 35982 40562 36034 40574
rect 37102 40626 37154 40638
rect 37102 40562 37154 40574
rect 38334 40626 38386 40638
rect 38334 40562 38386 40574
rect 38558 40626 38610 40638
rect 38558 40562 38610 40574
rect 38782 40626 38834 40638
rect 38782 40562 38834 40574
rect 39230 40626 39282 40638
rect 39230 40562 39282 40574
rect 40238 40626 40290 40638
rect 40238 40562 40290 40574
rect 46510 40626 46562 40638
rect 46510 40562 46562 40574
rect 46958 40626 47010 40638
rect 46958 40562 47010 40574
rect 47630 40626 47682 40638
rect 47630 40562 47682 40574
rect 2270 40514 2322 40526
rect 2270 40450 2322 40462
rect 2606 40514 2658 40526
rect 2606 40450 2658 40462
rect 2830 40514 2882 40526
rect 2830 40450 2882 40462
rect 3390 40514 3442 40526
rect 3390 40450 3442 40462
rect 6974 40514 7026 40526
rect 6974 40450 7026 40462
rect 9550 40514 9602 40526
rect 10894 40514 10946 40526
rect 10770 40462 10782 40514
rect 10834 40462 10846 40514
rect 9550 40450 9602 40462
rect 10894 40450 10946 40462
rect 11006 40514 11058 40526
rect 11006 40450 11058 40462
rect 12014 40514 12066 40526
rect 12014 40450 12066 40462
rect 12574 40514 12626 40526
rect 12574 40450 12626 40462
rect 13470 40514 13522 40526
rect 13470 40450 13522 40462
rect 16718 40514 16770 40526
rect 16718 40450 16770 40462
rect 17614 40514 17666 40526
rect 25790 40514 25842 40526
rect 23090 40462 23102 40514
rect 23154 40462 23166 40514
rect 24098 40462 24110 40514
rect 24162 40462 24174 40514
rect 17614 40450 17666 40462
rect 25790 40450 25842 40462
rect 25902 40514 25954 40526
rect 33070 40514 33122 40526
rect 29138 40462 29150 40514
rect 29202 40462 29214 40514
rect 30146 40462 30158 40514
rect 30210 40462 30222 40514
rect 32498 40462 32510 40514
rect 32562 40462 32574 40514
rect 25902 40450 25954 40462
rect 33070 40450 33122 40462
rect 35534 40514 35586 40526
rect 35534 40450 35586 40462
rect 35870 40514 35922 40526
rect 35870 40450 35922 40462
rect 36206 40514 36258 40526
rect 36206 40450 36258 40462
rect 36430 40514 36482 40526
rect 36430 40450 36482 40462
rect 36878 40514 36930 40526
rect 36878 40450 36930 40462
rect 39790 40514 39842 40526
rect 39790 40450 39842 40462
rect 40350 40514 40402 40526
rect 47406 40514 47458 40526
rect 41682 40462 41694 40514
rect 41746 40462 41758 40514
rect 44146 40462 44158 40514
rect 44210 40462 44222 40514
rect 46274 40462 46286 40514
rect 46338 40462 46350 40514
rect 40350 40450 40402 40462
rect 47406 40450 47458 40462
rect 47854 40514 47906 40526
rect 47854 40450 47906 40462
rect 3166 40402 3218 40414
rect 6862 40402 6914 40414
rect 3714 40350 3726 40402
rect 3778 40350 3790 40402
rect 3166 40338 3218 40350
rect 6862 40338 6914 40350
rect 7198 40402 7250 40414
rect 7198 40338 7250 40350
rect 7422 40402 7474 40414
rect 7422 40338 7474 40350
rect 8654 40402 8706 40414
rect 8654 40338 8706 40350
rect 9102 40402 9154 40414
rect 9102 40338 9154 40350
rect 11230 40402 11282 40414
rect 11230 40338 11282 40350
rect 11566 40402 11618 40414
rect 11566 40338 11618 40350
rect 11790 40402 11842 40414
rect 11790 40338 11842 40350
rect 13134 40402 13186 40414
rect 13134 40338 13186 40350
rect 15262 40402 15314 40414
rect 15262 40338 15314 40350
rect 15710 40402 15762 40414
rect 15710 40338 15762 40350
rect 16606 40402 16658 40414
rect 16606 40338 16658 40350
rect 17502 40402 17554 40414
rect 17502 40338 17554 40350
rect 18062 40402 18114 40414
rect 24446 40402 24498 40414
rect 27246 40402 27298 40414
rect 33294 40402 33346 40414
rect 36766 40402 36818 40414
rect 18386 40350 18398 40402
rect 18450 40350 18462 40402
rect 21970 40350 21982 40402
rect 22034 40350 22046 40402
rect 22978 40350 22990 40402
rect 23042 40350 23054 40402
rect 26450 40350 26462 40402
rect 26514 40350 26526 40402
rect 27906 40350 27918 40402
rect 27970 40350 27982 40402
rect 28578 40350 28590 40402
rect 28642 40350 28654 40402
rect 30258 40350 30270 40402
rect 30322 40350 30334 40402
rect 31154 40350 31166 40402
rect 31218 40350 31230 40402
rect 33730 40350 33742 40402
rect 33794 40350 33806 40402
rect 35074 40350 35086 40402
rect 35138 40350 35150 40402
rect 18062 40338 18114 40350
rect 24446 40338 24498 40350
rect 27246 40338 27298 40350
rect 33294 40338 33346 40350
rect 36766 40338 36818 40350
rect 37326 40402 37378 40414
rect 37326 40338 37378 40350
rect 38446 40402 38498 40414
rect 38446 40338 38498 40350
rect 40014 40402 40066 40414
rect 47070 40402 47122 40414
rect 41010 40350 41022 40402
rect 41074 40350 41086 40402
rect 44482 40350 44494 40402
rect 44546 40350 44558 40402
rect 44930 40350 44942 40402
rect 44994 40350 45006 40402
rect 45490 40350 45502 40402
rect 45554 40350 45566 40402
rect 45826 40350 45838 40402
rect 45890 40350 45902 40402
rect 40014 40338 40066 40350
rect 47070 40338 47122 40350
rect 47518 40402 47570 40414
rect 47518 40338 47570 40350
rect 4622 40290 4674 40302
rect 4622 40226 4674 40238
rect 13582 40290 13634 40302
rect 13582 40226 13634 40238
rect 14478 40290 14530 40302
rect 14478 40226 14530 40238
rect 16270 40290 16322 40302
rect 29038 40290 29090 40302
rect 19058 40238 19070 40290
rect 19122 40238 19134 40290
rect 21186 40238 21198 40290
rect 21250 40238 21262 40290
rect 35186 40238 35198 40290
rect 35250 40238 35262 40290
rect 37762 40238 37774 40290
rect 37826 40238 37838 40290
rect 43810 40238 43822 40290
rect 43874 40238 43886 40290
rect 16270 40226 16322 40238
rect 29038 40226 29090 40238
rect 4398 40178 4450 40190
rect 4398 40114 4450 40126
rect 7646 40178 7698 40190
rect 7646 40114 7698 40126
rect 9774 40178 9826 40190
rect 9774 40114 9826 40126
rect 1344 40010 48608 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 48608 40010
rect 1344 39924 48608 39958
rect 11790 39842 11842 39854
rect 11790 39778 11842 39790
rect 21422 39842 21474 39854
rect 21422 39778 21474 39790
rect 21758 39842 21810 39854
rect 21758 39778 21810 39790
rect 25006 39842 25058 39854
rect 25006 39778 25058 39790
rect 28254 39842 28306 39854
rect 28254 39778 28306 39790
rect 36318 39842 36370 39854
rect 36318 39778 36370 39790
rect 9662 39730 9714 39742
rect 19966 39730 20018 39742
rect 2482 39678 2494 39730
rect 2546 39678 2558 39730
rect 4610 39678 4622 39730
rect 4674 39678 4686 39730
rect 8530 39678 8542 39730
rect 8594 39678 8606 39730
rect 16930 39678 16942 39730
rect 16994 39678 17006 39730
rect 19394 39678 19406 39730
rect 19458 39678 19470 39730
rect 9662 39666 9714 39678
rect 19966 39666 20018 39678
rect 20638 39730 20690 39742
rect 20638 39666 20690 39678
rect 24558 39730 24610 39742
rect 27358 39730 27410 39742
rect 26002 39678 26014 39730
rect 26066 39678 26078 39730
rect 24558 39666 24610 39678
rect 27358 39666 27410 39678
rect 27806 39730 27858 39742
rect 33406 39730 33458 39742
rect 29250 39678 29262 39730
rect 29314 39678 29326 39730
rect 27806 39666 27858 39678
rect 33406 39666 33458 39678
rect 35086 39730 35138 39742
rect 35086 39666 35138 39678
rect 35982 39730 36034 39742
rect 35982 39666 36034 39678
rect 37550 39730 37602 39742
rect 42478 39730 42530 39742
rect 38210 39678 38222 39730
rect 38274 39678 38286 39730
rect 37550 39666 37602 39678
rect 42478 39666 42530 39678
rect 42702 39730 42754 39742
rect 42702 39666 42754 39678
rect 44382 39730 44434 39742
rect 45266 39678 45278 39730
rect 45330 39678 45342 39730
rect 44382 39666 44434 39678
rect 11118 39618 11170 39630
rect 1810 39566 1822 39618
rect 1874 39566 1886 39618
rect 5618 39566 5630 39618
rect 5682 39566 5694 39618
rect 11118 39554 11170 39566
rect 11678 39618 11730 39630
rect 11678 39554 11730 39566
rect 12350 39618 12402 39630
rect 12350 39554 12402 39566
rect 13022 39618 13074 39630
rect 13022 39554 13074 39566
rect 13806 39618 13858 39630
rect 20750 39618 20802 39630
rect 14130 39566 14142 39618
rect 14194 39566 14206 39618
rect 17938 39566 17950 39618
rect 18002 39566 18014 39618
rect 13806 39554 13858 39566
rect 20750 39554 20802 39566
rect 21982 39618 22034 39630
rect 21982 39554 22034 39566
rect 22318 39618 22370 39630
rect 22318 39554 22370 39566
rect 22878 39618 22930 39630
rect 24446 39618 24498 39630
rect 30158 39618 30210 39630
rect 33182 39618 33234 39630
rect 24098 39566 24110 39618
rect 24162 39566 24174 39618
rect 26114 39566 26126 39618
rect 26178 39566 26190 39618
rect 29474 39566 29486 39618
rect 29538 39566 29550 39618
rect 31154 39566 31166 39618
rect 31218 39566 31230 39618
rect 31826 39566 31838 39618
rect 31890 39566 31902 39618
rect 32498 39566 32510 39618
rect 32562 39566 32574 39618
rect 22878 39554 22930 39566
rect 24446 39554 24498 39566
rect 30158 39554 30210 39566
rect 33182 39554 33234 39566
rect 33742 39618 33794 39630
rect 33742 39554 33794 39566
rect 34414 39618 34466 39630
rect 34414 39554 34466 39566
rect 35534 39618 35586 39630
rect 35534 39554 35586 39566
rect 36430 39618 36482 39630
rect 36430 39554 36482 39566
rect 36990 39618 37042 39630
rect 36990 39554 37042 39566
rect 37214 39618 37266 39630
rect 37214 39554 37266 39566
rect 37438 39618 37490 39630
rect 41582 39618 41634 39630
rect 41122 39566 41134 39618
rect 41186 39566 41198 39618
rect 37438 39554 37490 39566
rect 41582 39554 41634 39566
rect 41694 39618 41746 39630
rect 41694 39554 41746 39566
rect 42030 39618 42082 39630
rect 43374 39618 43426 39630
rect 44046 39618 44098 39630
rect 42242 39566 42254 39618
rect 42306 39566 42318 39618
rect 43026 39566 43038 39618
rect 43090 39566 43102 39618
rect 43810 39566 43822 39618
rect 43874 39566 43886 39618
rect 48066 39566 48078 39618
rect 48130 39566 48142 39618
rect 42030 39554 42082 39566
rect 43374 39554 43426 39566
rect 44046 39554 44098 39566
rect 9998 39506 10050 39518
rect 6402 39454 6414 39506
rect 6466 39454 6478 39506
rect 9998 39442 10050 39454
rect 10334 39506 10386 39518
rect 10334 39442 10386 39454
rect 11230 39506 11282 39518
rect 11230 39442 11282 39454
rect 11790 39506 11842 39518
rect 11790 39442 11842 39454
rect 12574 39506 12626 39518
rect 12574 39442 12626 39454
rect 13470 39506 13522 39518
rect 20526 39506 20578 39518
rect 14802 39454 14814 39506
rect 14866 39454 14878 39506
rect 18834 39454 18846 39506
rect 18898 39454 18910 39506
rect 13470 39442 13522 39454
rect 20526 39442 20578 39454
rect 21534 39506 21586 39518
rect 21534 39442 21586 39454
rect 22206 39506 22258 39518
rect 24894 39506 24946 39518
rect 23202 39454 23214 39506
rect 23266 39454 23278 39506
rect 22206 39442 22258 39454
rect 24894 39442 24946 39454
rect 26798 39506 26850 39518
rect 26798 39442 26850 39454
rect 28142 39506 28194 39518
rect 33630 39506 33682 39518
rect 44830 39506 44882 39518
rect 32162 39454 32174 39506
rect 32226 39454 32238 39506
rect 32722 39454 32734 39506
rect 32786 39454 32798 39506
rect 40338 39454 40350 39506
rect 40402 39454 40414 39506
rect 47394 39454 47406 39506
rect 47458 39454 47470 39506
rect 28142 39442 28194 39454
rect 33630 39442 33682 39454
rect 44830 39442 44882 39454
rect 5070 39394 5122 39406
rect 9214 39394 9266 39406
rect 8866 39342 8878 39394
rect 8930 39342 8942 39394
rect 5070 39330 5122 39342
rect 9214 39330 9266 39342
rect 10894 39394 10946 39406
rect 10894 39330 10946 39342
rect 11454 39394 11506 39406
rect 11454 39330 11506 39342
rect 12798 39394 12850 39406
rect 12798 39330 12850 39342
rect 13582 39394 13634 39406
rect 25006 39394 25058 39406
rect 17378 39342 17390 39394
rect 17442 39342 17454 39394
rect 13582 39330 13634 39342
rect 25006 39330 25058 39342
rect 30606 39394 30658 39406
rect 30606 39330 30658 39342
rect 37662 39394 37714 39406
rect 37662 39330 37714 39342
rect 42478 39394 42530 39406
rect 42478 39330 42530 39342
rect 43262 39394 43314 39406
rect 43262 39330 43314 39342
rect 43822 39394 43874 39406
rect 43822 39330 43874 39342
rect 44942 39394 44994 39406
rect 44942 39330 44994 39342
rect 1344 39226 48608 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 48608 39226
rect 1344 39140 48608 39174
rect 4286 39058 4338 39070
rect 4286 38994 4338 39006
rect 4622 39058 4674 39070
rect 4622 38994 4674 39006
rect 5966 39058 6018 39070
rect 5966 38994 6018 39006
rect 8094 39058 8146 39070
rect 8094 38994 8146 39006
rect 9886 39058 9938 39070
rect 9886 38994 9938 39006
rect 11118 39058 11170 39070
rect 11118 38994 11170 39006
rect 11342 39058 11394 39070
rect 11342 38994 11394 39006
rect 14926 39058 14978 39070
rect 14926 38994 14978 39006
rect 15934 39058 15986 39070
rect 15934 38994 15986 39006
rect 17838 39058 17890 39070
rect 17838 38994 17890 39006
rect 17950 39058 18002 39070
rect 17950 38994 18002 39006
rect 20974 39058 21026 39070
rect 20974 38994 21026 39006
rect 22654 39058 22706 39070
rect 22654 38994 22706 39006
rect 23214 39058 23266 39070
rect 23214 38994 23266 39006
rect 28590 39058 28642 39070
rect 28590 38994 28642 39006
rect 29038 39058 29090 39070
rect 29038 38994 29090 39006
rect 32062 39058 32114 39070
rect 32062 38994 32114 39006
rect 35198 39058 35250 39070
rect 35198 38994 35250 39006
rect 36766 39058 36818 39070
rect 36766 38994 36818 39006
rect 40014 39058 40066 39070
rect 40014 38994 40066 39006
rect 41022 39058 41074 39070
rect 41022 38994 41074 39006
rect 42030 39058 42082 39070
rect 42030 38994 42082 39006
rect 42366 39058 42418 39070
rect 42366 38994 42418 39006
rect 44270 39058 44322 39070
rect 44270 38994 44322 39006
rect 44830 39058 44882 39070
rect 44830 38994 44882 39006
rect 2494 38946 2546 38958
rect 2494 38882 2546 38894
rect 4846 38946 4898 38958
rect 4846 38882 4898 38894
rect 8318 38946 8370 38958
rect 8318 38882 8370 38894
rect 9662 38946 9714 38958
rect 9662 38882 9714 38894
rect 10558 38946 10610 38958
rect 10558 38882 10610 38894
rect 11006 38946 11058 38958
rect 11006 38882 11058 38894
rect 13918 38946 13970 38958
rect 13918 38882 13970 38894
rect 14366 38946 14418 38958
rect 14366 38882 14418 38894
rect 15374 38946 15426 38958
rect 15374 38882 15426 38894
rect 15598 38946 15650 38958
rect 15598 38882 15650 38894
rect 19854 38946 19906 38958
rect 19854 38882 19906 38894
rect 20302 38946 20354 38958
rect 20302 38882 20354 38894
rect 21310 38946 21362 38958
rect 21310 38882 21362 38894
rect 21758 38946 21810 38958
rect 21758 38882 21810 38894
rect 21870 38946 21922 38958
rect 21870 38882 21922 38894
rect 22318 38946 22370 38958
rect 22318 38882 22370 38894
rect 22430 38946 22482 38958
rect 22430 38882 22482 38894
rect 22990 38946 23042 38958
rect 22990 38882 23042 38894
rect 24558 38946 24610 38958
rect 24558 38882 24610 38894
rect 25454 38946 25506 38958
rect 25454 38882 25506 38894
rect 27694 38946 27746 38958
rect 27694 38882 27746 38894
rect 29150 38946 29202 38958
rect 34078 38946 34130 38958
rect 40910 38946 40962 38958
rect 31266 38894 31278 38946
rect 31330 38894 31342 38946
rect 37538 38894 37550 38946
rect 37602 38894 37614 38946
rect 29150 38882 29202 38894
rect 34078 38882 34130 38894
rect 40910 38882 40962 38894
rect 42478 38946 42530 38958
rect 44482 38894 44494 38946
rect 44546 38894 44558 38946
rect 42478 38882 42530 38894
rect 4174 38834 4226 38846
rect 3154 38782 3166 38834
rect 3218 38782 3230 38834
rect 3826 38782 3838 38834
rect 3890 38782 3902 38834
rect 4174 38770 4226 38782
rect 4398 38834 4450 38846
rect 4398 38770 4450 38782
rect 4958 38834 5010 38846
rect 4958 38770 5010 38782
rect 5630 38834 5682 38846
rect 5630 38770 5682 38782
rect 5854 38834 5906 38846
rect 5854 38770 5906 38782
rect 6190 38834 6242 38846
rect 7646 38834 7698 38846
rect 6962 38782 6974 38834
rect 7026 38782 7038 38834
rect 6190 38770 6242 38782
rect 7646 38770 7698 38782
rect 8206 38834 8258 38846
rect 8206 38770 8258 38782
rect 9550 38834 9602 38846
rect 9550 38770 9602 38782
rect 10334 38834 10386 38846
rect 10334 38770 10386 38782
rect 10670 38834 10722 38846
rect 14254 38834 14306 38846
rect 13010 38782 13022 38834
rect 13074 38782 13086 38834
rect 10670 38770 10722 38782
rect 14254 38770 14306 38782
rect 14590 38834 14642 38846
rect 14590 38770 14642 38782
rect 16046 38834 16098 38846
rect 17278 38834 17330 38846
rect 16370 38782 16382 38834
rect 16434 38782 16446 38834
rect 16046 38770 16098 38782
rect 17278 38770 17330 38782
rect 17726 38834 17778 38846
rect 17726 38770 17778 38782
rect 20750 38834 20802 38846
rect 20750 38770 20802 38782
rect 20974 38834 21026 38846
rect 20974 38770 21026 38782
rect 22878 38834 22930 38846
rect 27470 38834 27522 38846
rect 23650 38782 23662 38834
rect 23714 38782 23726 38834
rect 26002 38782 26014 38834
rect 26066 38782 26078 38834
rect 26226 38782 26238 38834
rect 26290 38782 26302 38834
rect 27234 38782 27246 38834
rect 27298 38782 27310 38834
rect 22878 38770 22930 38782
rect 27470 38770 27522 38782
rect 27806 38834 27858 38846
rect 34750 38834 34802 38846
rect 29698 38782 29710 38834
rect 29762 38782 29774 38834
rect 30034 38782 30046 38834
rect 30098 38782 30110 38834
rect 33394 38782 33406 38834
rect 33458 38782 33470 38834
rect 27806 38770 27858 38782
rect 34750 38770 34802 38782
rect 34974 38834 35026 38846
rect 34974 38770 35026 38782
rect 36542 38834 36594 38846
rect 43038 38834 43090 38846
rect 38098 38782 38110 38834
rect 38162 38782 38174 38834
rect 38770 38782 38782 38834
rect 38834 38782 38846 38834
rect 36542 38770 36594 38782
rect 43038 38770 43090 38782
rect 43150 38834 43202 38846
rect 43150 38770 43202 38782
rect 43262 38834 43314 38846
rect 44158 38834 44210 38846
rect 43698 38782 43710 38834
rect 43762 38782 43774 38834
rect 48066 38782 48078 38834
rect 48130 38782 48142 38834
rect 43262 38770 43314 38782
rect 44158 38770 44210 38782
rect 6414 38722 6466 38734
rect 8878 38722 8930 38734
rect 3378 38670 3390 38722
rect 3442 38670 3454 38722
rect 6850 38670 6862 38722
rect 6914 38670 6926 38722
rect 6414 38658 6466 38670
rect 8878 38658 8930 38670
rect 12014 38722 12066 38734
rect 12014 38658 12066 38670
rect 12574 38722 12626 38734
rect 18398 38722 18450 38734
rect 13122 38670 13134 38722
rect 13186 38670 13198 38722
rect 15250 38670 15262 38722
rect 15314 38670 15326 38722
rect 12574 38658 12626 38670
rect 18398 38658 18450 38670
rect 18958 38722 19010 38734
rect 18958 38658 19010 38670
rect 19406 38722 19458 38734
rect 21646 38722 21698 38734
rect 28926 38722 28978 38734
rect 20402 38670 20414 38722
rect 20466 38670 20478 38722
rect 24098 38670 24110 38722
rect 24162 38670 24174 38722
rect 25554 38670 25566 38722
rect 25618 38670 25630 38722
rect 27010 38670 27022 38722
rect 27074 38670 27086 38722
rect 19406 38658 19458 38670
rect 21646 38658 21698 38670
rect 28926 38658 28978 38670
rect 32510 38722 32562 38734
rect 34862 38722 34914 38734
rect 36094 38722 36146 38734
rect 39454 38722 39506 38734
rect 33170 38670 33182 38722
rect 33234 38670 33246 38722
rect 35746 38670 35758 38722
rect 35810 38670 35822 38722
rect 36866 38670 36878 38722
rect 36930 38670 36942 38722
rect 32510 38658 32562 38670
rect 34862 38658 34914 38670
rect 36094 38658 36146 38670
rect 39454 38658 39506 38670
rect 39790 38722 39842 38734
rect 43822 38722 43874 38734
rect 40114 38670 40126 38722
rect 40178 38670 40190 38722
rect 41570 38670 41582 38722
rect 41634 38670 41646 38722
rect 47394 38670 47406 38722
rect 47458 38670 47470 38722
rect 39790 38658 39842 38670
rect 43822 38658 43874 38670
rect 16382 38610 16434 38622
rect 16382 38546 16434 38558
rect 16718 38610 16770 38622
rect 20078 38610 20130 38622
rect 18498 38558 18510 38610
rect 18562 38607 18574 38610
rect 19394 38607 19406 38610
rect 18562 38561 19406 38607
rect 18562 38558 18574 38561
rect 19394 38558 19406 38561
rect 19458 38558 19470 38610
rect 16718 38546 16770 38558
rect 20078 38546 20130 38558
rect 25230 38610 25282 38622
rect 45266 38614 45278 38666
rect 45330 38614 45342 38666
rect 25230 38546 25282 38558
rect 1344 38442 48608 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 48608 38442
rect 1344 38356 48608 38390
rect 3614 38274 3666 38286
rect 31390 38274 31442 38286
rect 5618 38222 5630 38274
rect 5682 38271 5694 38274
rect 6178 38271 6190 38274
rect 5682 38225 6190 38271
rect 5682 38222 5694 38225
rect 6178 38222 6190 38225
rect 6242 38222 6254 38274
rect 3614 38210 3666 38222
rect 31390 38210 31442 38222
rect 3166 38162 3218 38174
rect 3166 38098 3218 38110
rect 5070 38162 5122 38174
rect 5070 38098 5122 38110
rect 8318 38162 8370 38174
rect 23998 38162 24050 38174
rect 35870 38162 35922 38174
rect 15026 38110 15038 38162
rect 15090 38110 15102 38162
rect 15586 38110 15598 38162
rect 15650 38110 15662 38162
rect 16258 38110 16270 38162
rect 16322 38110 16334 38162
rect 20290 38110 20302 38162
rect 20354 38110 20366 38162
rect 25666 38110 25678 38162
rect 25730 38110 25742 38162
rect 29586 38110 29598 38162
rect 29650 38110 29662 38162
rect 34850 38110 34862 38162
rect 34914 38110 34926 38162
rect 8318 38098 8370 38110
rect 23998 38098 24050 38110
rect 35870 38098 35922 38110
rect 37102 38162 37154 38174
rect 44034 38110 44046 38162
rect 44098 38110 44110 38162
rect 44930 38110 44942 38162
rect 44994 38110 45006 38162
rect 37102 38098 37154 38110
rect 3726 38050 3778 38062
rect 3726 37986 3778 37998
rect 4174 38050 4226 38062
rect 4174 37986 4226 37998
rect 4734 38050 4786 38062
rect 4734 37986 4786 37998
rect 6414 38050 6466 38062
rect 6414 37986 6466 37998
rect 6638 38050 6690 38062
rect 6638 37986 6690 37998
rect 7086 38050 7138 38062
rect 7086 37986 7138 37998
rect 10334 38050 10386 38062
rect 10334 37986 10386 37998
rect 11230 38050 11282 38062
rect 23886 38050 23938 38062
rect 12450 37998 12462 38050
rect 12514 37998 12526 38050
rect 13570 37998 13582 38050
rect 13634 37998 13646 38050
rect 13906 37998 13918 38050
rect 13970 37998 13982 38050
rect 15362 37998 15374 38050
rect 15426 37998 15438 38050
rect 16146 37998 16158 38050
rect 16210 37998 16222 38050
rect 17490 37998 17502 38050
rect 17554 37998 17566 38050
rect 21298 37998 21310 38050
rect 21362 37998 21374 38050
rect 23538 37998 23550 38050
rect 23602 37998 23614 38050
rect 11230 37986 11282 37998
rect 23886 37986 23938 37998
rect 24334 38050 24386 38062
rect 30046 38050 30098 38062
rect 47630 38050 47682 38062
rect 28466 37998 28478 38050
rect 28530 37998 28542 38050
rect 30258 37998 30270 38050
rect 30322 37998 30334 38050
rect 31938 37998 31950 38050
rect 32002 37998 32014 38050
rect 41122 37998 41134 38050
rect 41186 37998 41198 38050
rect 24334 37986 24386 37998
rect 30046 37986 30098 37998
rect 47630 37986 47682 37998
rect 10446 37938 10498 37950
rect 8642 37886 8654 37938
rect 8706 37886 8718 37938
rect 9650 37886 9662 37938
rect 9714 37886 9726 37938
rect 10446 37874 10498 37886
rect 10894 37938 10946 37950
rect 21534 37938 21586 37950
rect 18162 37886 18174 37938
rect 18226 37886 18238 37938
rect 10894 37874 10946 37886
rect 21534 37874 21586 37886
rect 21646 37938 21698 37950
rect 27806 37938 27858 37950
rect 22306 37886 22318 37938
rect 22370 37886 22382 37938
rect 24658 37886 24670 37938
rect 24722 37886 24734 37938
rect 26002 37886 26014 37938
rect 26066 37886 26078 37938
rect 27570 37886 27582 37938
rect 27634 37886 27646 37938
rect 21646 37874 21698 37886
rect 27806 37874 27858 37886
rect 28142 37938 28194 37950
rect 28142 37874 28194 37886
rect 29262 37938 29314 37950
rect 29262 37874 29314 37886
rect 30942 37938 30994 37950
rect 30942 37874 30994 37886
rect 31502 37938 31554 37950
rect 36206 37938 36258 37950
rect 32722 37886 32734 37938
rect 32786 37886 32798 37938
rect 31502 37874 31554 37886
rect 36206 37874 36258 37886
rect 36990 37938 37042 37950
rect 36990 37874 37042 37886
rect 37774 37938 37826 37950
rect 37774 37874 37826 37886
rect 40686 37938 40738 37950
rect 40686 37874 40738 37886
rect 40798 37938 40850 37950
rect 41906 37886 41918 37938
rect 41970 37886 41982 37938
rect 45154 37886 45166 37938
rect 45218 37886 45230 37938
rect 46834 37886 46846 37938
rect 46898 37886 46910 37938
rect 40798 37874 40850 37886
rect 2270 37826 2322 37838
rect 2270 37762 2322 37774
rect 3614 37826 3666 37838
rect 3614 37762 3666 37774
rect 4062 37826 4114 37838
rect 4062 37762 4114 37774
rect 4286 37826 4338 37838
rect 4286 37762 4338 37774
rect 5742 37826 5794 37838
rect 5742 37762 5794 37774
rect 6526 37826 6578 37838
rect 6526 37762 6578 37774
rect 7646 37826 7698 37838
rect 7646 37762 7698 37774
rect 8990 37826 9042 37838
rect 8990 37762 9042 37774
rect 9326 37826 9378 37838
rect 9326 37762 9378 37774
rect 10670 37826 10722 37838
rect 10670 37762 10722 37774
rect 11006 37826 11058 37838
rect 11006 37762 11058 37774
rect 11566 37826 11618 37838
rect 11566 37762 11618 37774
rect 11902 37826 11954 37838
rect 11902 37762 11954 37774
rect 12014 37826 12066 37838
rect 12014 37762 12066 37774
rect 12126 37826 12178 37838
rect 12126 37762 12178 37774
rect 13022 37826 13074 37838
rect 13022 37762 13074 37774
rect 20750 37826 20802 37838
rect 20750 37762 20802 37774
rect 22654 37826 22706 37838
rect 22654 37762 22706 37774
rect 25230 37826 25282 37838
rect 25230 37762 25282 37774
rect 28254 37826 28306 37838
rect 28254 37762 28306 37774
rect 29486 37826 29538 37838
rect 29486 37762 29538 37774
rect 31390 37826 31442 37838
rect 31390 37762 31442 37774
rect 35310 37826 35362 37838
rect 35310 37762 35362 37774
rect 36318 37826 36370 37838
rect 36318 37762 36370 37774
rect 36542 37826 36594 37838
rect 36542 37762 36594 37774
rect 37214 37826 37266 37838
rect 37214 37762 37266 37774
rect 37662 37826 37714 37838
rect 37662 37762 37714 37774
rect 38222 37826 38274 37838
rect 38222 37762 38274 37774
rect 38782 37826 38834 37838
rect 38782 37762 38834 37774
rect 39118 37826 39170 37838
rect 39118 37762 39170 37774
rect 39902 37826 39954 37838
rect 39902 37762 39954 37774
rect 40350 37826 40402 37838
rect 48190 37826 48242 37838
rect 46722 37774 46734 37826
rect 46786 37774 46798 37826
rect 40350 37762 40402 37774
rect 48190 37762 48242 37774
rect 1344 37658 48608 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 48608 37658
rect 1344 37572 48608 37606
rect 5406 37490 5458 37502
rect 5406 37426 5458 37438
rect 6638 37490 6690 37502
rect 6638 37426 6690 37438
rect 7646 37490 7698 37502
rect 34414 37490 34466 37502
rect 21634 37438 21646 37490
rect 21698 37438 21710 37490
rect 7646 37426 7698 37438
rect 34414 37426 34466 37438
rect 41022 37490 41074 37502
rect 41022 37426 41074 37438
rect 43486 37490 43538 37502
rect 43486 37426 43538 37438
rect 6862 37378 6914 37390
rect 6862 37314 6914 37326
rect 10670 37378 10722 37390
rect 16494 37378 16546 37390
rect 14690 37326 14702 37378
rect 14754 37326 14766 37378
rect 10670 37314 10722 37326
rect 16494 37314 16546 37326
rect 19182 37378 19234 37390
rect 23774 37378 23826 37390
rect 34302 37378 34354 37390
rect 20290 37326 20302 37378
rect 20354 37326 20366 37378
rect 21522 37326 21534 37378
rect 21586 37326 21598 37378
rect 29250 37326 29262 37378
rect 29314 37326 29326 37378
rect 19182 37314 19234 37326
rect 23774 37314 23826 37326
rect 34302 37314 34354 37326
rect 34862 37378 34914 37390
rect 34862 37314 34914 37326
rect 35198 37378 35250 37390
rect 35198 37314 35250 37326
rect 36990 37378 37042 37390
rect 41122 37326 41134 37378
rect 41186 37326 41198 37378
rect 43026 37326 43038 37378
rect 43090 37326 43102 37378
rect 47058 37326 47070 37378
rect 47122 37326 47134 37378
rect 36990 37314 37042 37326
rect 4846 37266 4898 37278
rect 1810 37214 1822 37266
rect 1874 37214 1886 37266
rect 4846 37202 4898 37214
rect 5294 37266 5346 37278
rect 5294 37202 5346 37214
rect 5518 37266 5570 37278
rect 5518 37202 5570 37214
rect 5742 37266 5794 37278
rect 5742 37202 5794 37214
rect 6190 37266 6242 37278
rect 6190 37202 6242 37214
rect 6302 37266 6354 37278
rect 6302 37202 6354 37214
rect 6974 37266 7026 37278
rect 9774 37266 9826 37278
rect 17502 37266 17554 37278
rect 8418 37214 8430 37266
rect 8482 37214 8494 37266
rect 8754 37214 8766 37266
rect 8818 37214 8830 37266
rect 10210 37214 10222 37266
rect 10274 37214 10286 37266
rect 10994 37214 11006 37266
rect 11058 37214 11070 37266
rect 15922 37214 15934 37266
rect 15986 37214 15998 37266
rect 6974 37202 7026 37214
rect 9774 37202 9826 37214
rect 17502 37202 17554 37214
rect 18734 37266 18786 37278
rect 18734 37202 18786 37214
rect 19070 37266 19122 37278
rect 19070 37202 19122 37214
rect 19406 37266 19458 37278
rect 32510 37266 32562 37278
rect 23202 37214 23214 37266
rect 23266 37214 23278 37266
rect 30034 37214 30046 37266
rect 30098 37214 30110 37266
rect 30818 37214 30830 37266
rect 30882 37214 30894 37266
rect 31042 37214 31054 37266
rect 31106 37214 31118 37266
rect 31714 37214 31726 37266
rect 31778 37214 31790 37266
rect 19406 37202 19458 37214
rect 32510 37202 32562 37214
rect 33518 37266 33570 37278
rect 33518 37202 33570 37214
rect 34638 37266 34690 37278
rect 36766 37266 36818 37278
rect 35410 37214 35422 37266
rect 35474 37214 35486 37266
rect 35858 37214 35870 37266
rect 35922 37214 35934 37266
rect 34638 37202 34690 37214
rect 36766 37202 36818 37214
rect 37102 37266 37154 37278
rect 42702 37266 42754 37278
rect 37426 37214 37438 37266
rect 37490 37214 37502 37266
rect 41682 37214 41694 37266
rect 41746 37214 41758 37266
rect 41906 37214 41918 37266
rect 41970 37214 41982 37266
rect 37102 37202 37154 37214
rect 42702 37202 42754 37214
rect 44494 37266 44546 37278
rect 47730 37214 47742 37266
rect 47794 37214 47806 37266
rect 44494 37202 44546 37214
rect 5966 37154 6018 37166
rect 2482 37102 2494 37154
rect 2546 37102 2558 37154
rect 4610 37102 4622 37154
rect 4674 37102 4686 37154
rect 5966 37090 6018 37102
rect 8990 37154 9042 37166
rect 18398 37154 18450 37166
rect 22318 37154 22370 37166
rect 26350 37154 26402 37166
rect 11778 37102 11790 37154
rect 11842 37102 11854 37154
rect 13906 37102 13918 37154
rect 13970 37102 13982 37154
rect 14354 37102 14366 37154
rect 14418 37102 14430 37154
rect 19730 37102 19742 37154
rect 19794 37102 19806 37154
rect 22978 37102 22990 37154
rect 23042 37102 23054 37154
rect 8990 37090 9042 37102
rect 18398 37090 18450 37102
rect 22318 37090 22370 37102
rect 26350 37090 26402 37102
rect 26798 37154 26850 37166
rect 33966 37154 34018 37166
rect 43934 37154 43986 37166
rect 27122 37102 27134 37154
rect 27186 37102 27198 37154
rect 31826 37102 31838 37154
rect 31890 37102 31902 37154
rect 38210 37102 38222 37154
rect 38274 37102 38286 37154
rect 40338 37102 40350 37154
rect 40402 37102 40414 37154
rect 44930 37102 44942 37154
rect 44994 37102 45006 37154
rect 26798 37090 26850 37102
rect 33966 37090 34018 37102
rect 43934 37090 43986 37102
rect 17390 37042 17442 37054
rect 17390 36978 17442 36990
rect 1344 36874 48608 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 48608 36874
rect 1344 36788 48608 36822
rect 5854 36706 5906 36718
rect 5854 36642 5906 36654
rect 8430 36706 8482 36718
rect 10446 36706 10498 36718
rect 9986 36654 9998 36706
rect 10050 36654 10062 36706
rect 8430 36642 8482 36654
rect 10446 36642 10498 36654
rect 14702 36706 14754 36718
rect 14702 36642 14754 36654
rect 15038 36706 15090 36718
rect 27582 36706 27634 36718
rect 46846 36706 46898 36718
rect 21858 36654 21870 36706
rect 21922 36654 21934 36706
rect 37986 36654 37998 36706
rect 38050 36654 38062 36706
rect 15038 36642 15090 36654
rect 27582 36642 27634 36654
rect 46846 36642 46898 36654
rect 4510 36594 4562 36606
rect 4510 36530 4562 36542
rect 7310 36594 7362 36606
rect 7310 36530 7362 36542
rect 8766 36594 8818 36606
rect 21310 36594 21362 36606
rect 38670 36594 38722 36606
rect 10882 36542 10894 36594
rect 10946 36542 10958 36594
rect 15362 36542 15374 36594
rect 15426 36542 15438 36594
rect 17490 36542 17502 36594
rect 17554 36542 17566 36594
rect 23762 36542 23774 36594
rect 23826 36542 23838 36594
rect 31042 36542 31054 36594
rect 31106 36542 31118 36594
rect 35074 36542 35086 36594
rect 35138 36542 35150 36594
rect 36306 36542 36318 36594
rect 36370 36542 36382 36594
rect 8766 36530 8818 36542
rect 21310 36530 21362 36542
rect 38670 36530 38722 36542
rect 40798 36594 40850 36606
rect 40798 36530 40850 36542
rect 43150 36594 43202 36606
rect 43150 36530 43202 36542
rect 45838 36594 45890 36606
rect 47618 36542 47630 36594
rect 47682 36542 47694 36594
rect 45838 36530 45890 36542
rect 4398 36482 4450 36494
rect 4050 36430 4062 36482
rect 4114 36430 4126 36482
rect 4398 36418 4450 36430
rect 6526 36482 6578 36494
rect 6526 36418 6578 36430
rect 7198 36482 7250 36494
rect 7198 36418 7250 36430
rect 8206 36482 8258 36494
rect 9438 36482 9490 36494
rect 11902 36482 11954 36494
rect 9202 36430 9214 36482
rect 9266 36430 9278 36482
rect 10546 36430 10558 36482
rect 10610 36430 10622 36482
rect 11330 36430 11342 36482
rect 11394 36430 11406 36482
rect 8206 36418 8258 36430
rect 9438 36418 9490 36430
rect 11902 36418 11954 36430
rect 12350 36482 12402 36494
rect 12350 36418 12402 36430
rect 12462 36482 12514 36494
rect 12462 36418 12514 36430
rect 13918 36482 13970 36494
rect 13918 36418 13970 36430
rect 14142 36482 14194 36494
rect 18734 36482 18786 36494
rect 15026 36430 15038 36482
rect 15090 36430 15102 36482
rect 18274 36430 18286 36482
rect 18338 36430 18350 36482
rect 14142 36418 14194 36430
rect 18734 36418 18786 36430
rect 18846 36482 18898 36494
rect 18846 36418 18898 36430
rect 19966 36482 20018 36494
rect 19966 36418 20018 36430
rect 20414 36482 20466 36494
rect 20414 36418 20466 36430
rect 20526 36482 20578 36494
rect 20526 36418 20578 36430
rect 21534 36482 21586 36494
rect 21534 36418 21586 36430
rect 22206 36482 22258 36494
rect 22206 36418 22258 36430
rect 22430 36482 22482 36494
rect 27358 36482 27410 36494
rect 32958 36482 33010 36494
rect 34190 36482 34242 36494
rect 22754 36430 22766 36482
rect 22818 36430 22830 36482
rect 23090 36430 23102 36482
rect 23154 36430 23166 36482
rect 23986 36430 23998 36482
rect 24050 36430 24062 36482
rect 26562 36430 26574 36482
rect 26626 36430 26638 36482
rect 26786 36430 26798 36482
rect 26850 36430 26862 36482
rect 30370 36430 30382 36482
rect 30434 36430 30446 36482
rect 30930 36430 30942 36482
rect 30994 36430 31006 36482
rect 33618 36430 33630 36482
rect 33682 36430 33694 36482
rect 22430 36418 22482 36430
rect 27358 36418 27410 36430
rect 32958 36418 33010 36430
rect 34190 36418 34242 36430
rect 36206 36482 36258 36494
rect 36206 36418 36258 36430
rect 39230 36482 39282 36494
rect 39230 36418 39282 36430
rect 39342 36482 39394 36494
rect 39342 36418 39394 36430
rect 39678 36482 39730 36494
rect 39678 36418 39730 36430
rect 41582 36482 41634 36494
rect 41582 36418 41634 36430
rect 42142 36482 42194 36494
rect 42142 36418 42194 36430
rect 42254 36482 42306 36494
rect 42254 36418 42306 36430
rect 44830 36482 44882 36494
rect 46062 36482 46114 36494
rect 45490 36430 45502 36482
rect 45554 36430 45566 36482
rect 46610 36430 46622 36482
rect 46674 36430 46686 36482
rect 47394 36430 47406 36482
rect 47458 36430 47470 36482
rect 44830 36418 44882 36430
rect 46062 36418 46114 36430
rect 4958 36370 5010 36382
rect 4958 36306 5010 36318
rect 5070 36370 5122 36382
rect 5070 36306 5122 36318
rect 5854 36370 5906 36382
rect 5854 36306 5906 36318
rect 5966 36370 6018 36382
rect 5966 36306 6018 36318
rect 6302 36370 6354 36382
rect 6302 36306 6354 36318
rect 6862 36370 6914 36382
rect 6862 36306 6914 36318
rect 7422 36370 7474 36382
rect 7422 36306 7474 36318
rect 9550 36370 9602 36382
rect 9550 36306 9602 36318
rect 13582 36370 13634 36382
rect 13582 36306 13634 36318
rect 19182 36370 19234 36382
rect 19742 36370 19794 36382
rect 27022 36370 27074 36382
rect 19182 36306 19234 36318
rect 19630 36314 19682 36326
rect 1822 36258 1874 36270
rect 1822 36194 1874 36206
rect 2270 36258 2322 36270
rect 2270 36194 2322 36206
rect 2718 36258 2770 36270
rect 2718 36194 2770 36206
rect 3166 36258 3218 36270
rect 3166 36194 3218 36206
rect 4734 36258 4786 36270
rect 4734 36194 4786 36206
rect 6414 36258 6466 36270
rect 6414 36194 6466 36206
rect 7646 36258 7698 36270
rect 7646 36194 7698 36206
rect 12126 36258 12178 36270
rect 12126 36194 12178 36206
rect 13694 36258 13746 36270
rect 13694 36194 13746 36206
rect 14254 36258 14306 36270
rect 14254 36194 14306 36206
rect 14478 36258 14530 36270
rect 14478 36194 14530 36206
rect 19070 36258 19122 36270
rect 19070 36194 19122 36206
rect 19406 36258 19458 36270
rect 23202 36318 23214 36370
rect 23266 36318 23278 36370
rect 19742 36306 19794 36318
rect 27022 36306 27074 36318
rect 29150 36370 29202 36382
rect 31838 36370 31890 36382
rect 31042 36318 31054 36370
rect 31106 36318 31118 36370
rect 29150 36306 29202 36318
rect 31838 36306 31890 36318
rect 32398 36370 32450 36382
rect 32398 36306 32450 36318
rect 34302 36370 34354 36382
rect 34302 36306 34354 36318
rect 34638 36370 34690 36382
rect 34638 36306 34690 36318
rect 35758 36370 35810 36382
rect 35758 36306 35810 36318
rect 36990 36370 37042 36382
rect 36990 36306 37042 36318
rect 38558 36370 38610 36382
rect 38558 36306 38610 36318
rect 42366 36370 42418 36382
rect 42366 36306 42418 36318
rect 42702 36370 42754 36382
rect 42702 36306 42754 36318
rect 43486 36370 43538 36382
rect 43486 36306 43538 36318
rect 19630 36250 19682 36262
rect 20638 36258 20690 36270
rect 19406 36194 19458 36206
rect 20638 36194 20690 36206
rect 24670 36258 24722 36270
rect 24670 36194 24722 36206
rect 25118 36258 25170 36270
rect 28590 36258 28642 36270
rect 27906 36206 27918 36258
rect 27970 36206 27982 36258
rect 25118 36194 25170 36206
rect 28590 36194 28642 36206
rect 29262 36258 29314 36270
rect 29262 36194 29314 36206
rect 29374 36258 29426 36270
rect 29374 36194 29426 36206
rect 29598 36258 29650 36270
rect 29598 36194 29650 36206
rect 31950 36258 32002 36270
rect 31950 36194 32002 36206
rect 32174 36258 32226 36270
rect 32174 36194 32226 36206
rect 35982 36258 36034 36270
rect 35982 36194 36034 36206
rect 36318 36258 36370 36270
rect 36318 36194 36370 36206
rect 38782 36258 38834 36270
rect 38782 36194 38834 36206
rect 39566 36258 39618 36270
rect 39566 36194 39618 36206
rect 40126 36258 40178 36270
rect 40126 36194 40178 36206
rect 41134 36258 41186 36270
rect 41134 36194 41186 36206
rect 41246 36258 41298 36270
rect 41246 36194 41298 36206
rect 41358 36258 41410 36270
rect 41358 36194 41410 36206
rect 41470 36258 41522 36270
rect 41470 36194 41522 36206
rect 42478 36258 42530 36270
rect 42478 36194 42530 36206
rect 43598 36258 43650 36270
rect 43598 36194 43650 36206
rect 43934 36258 43986 36270
rect 45166 36258 45218 36270
rect 44258 36206 44270 36258
rect 44322 36206 44334 36258
rect 43934 36194 43986 36206
rect 45166 36194 45218 36206
rect 45726 36258 45778 36270
rect 45726 36194 45778 36206
rect 45950 36258 46002 36270
rect 45950 36194 46002 36206
rect 1344 36090 48608 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 48608 36090
rect 1344 36004 48608 36038
rect 5742 35922 5794 35934
rect 5742 35858 5794 35870
rect 7534 35922 7586 35934
rect 7534 35858 7586 35870
rect 7646 35922 7698 35934
rect 9774 35922 9826 35934
rect 8530 35870 8542 35922
rect 8594 35870 8606 35922
rect 7646 35858 7698 35870
rect 9774 35858 9826 35870
rect 10222 35922 10274 35934
rect 10222 35858 10274 35870
rect 12686 35922 12738 35934
rect 15150 35922 15202 35934
rect 13682 35870 13694 35922
rect 13746 35870 13758 35922
rect 12686 35858 12738 35870
rect 15150 35858 15202 35870
rect 23662 35922 23714 35934
rect 39342 35922 39394 35934
rect 28130 35870 28142 35922
rect 28194 35870 28206 35922
rect 34962 35870 34974 35922
rect 35026 35870 35038 35922
rect 23662 35858 23714 35870
rect 39342 35858 39394 35870
rect 43150 35922 43202 35934
rect 43150 35858 43202 35870
rect 44158 35922 44210 35934
rect 44158 35858 44210 35870
rect 44830 35922 44882 35934
rect 44830 35858 44882 35870
rect 7086 35810 7138 35822
rect 2482 35758 2494 35810
rect 2546 35758 2558 35810
rect 7086 35746 7138 35758
rect 7422 35810 7474 35822
rect 7422 35746 7474 35758
rect 9998 35810 10050 35822
rect 9998 35746 10050 35758
rect 11790 35810 11842 35822
rect 15710 35810 15762 35822
rect 14018 35758 14030 35810
rect 14082 35758 14094 35810
rect 11790 35746 11842 35758
rect 15710 35746 15762 35758
rect 16494 35810 16546 35822
rect 16494 35746 16546 35758
rect 16830 35810 16882 35822
rect 23326 35810 23378 35822
rect 18162 35758 18174 35810
rect 18226 35758 18238 35810
rect 16830 35746 16882 35758
rect 23326 35746 23378 35758
rect 26238 35810 26290 35822
rect 26238 35746 26290 35758
rect 27694 35810 27746 35822
rect 30046 35810 30098 35822
rect 29138 35758 29150 35810
rect 29202 35758 29214 35810
rect 27694 35746 27746 35758
rect 30046 35746 30098 35758
rect 30158 35810 30210 35822
rect 30158 35746 30210 35758
rect 32286 35810 32338 35822
rect 38894 35810 38946 35822
rect 33506 35758 33518 35810
rect 33570 35758 33582 35810
rect 32286 35746 32338 35758
rect 38894 35746 38946 35758
rect 39902 35810 39954 35822
rect 39902 35746 39954 35758
rect 42142 35810 42194 35822
rect 42142 35746 42194 35758
rect 44718 35810 44770 35822
rect 46050 35758 46062 35810
rect 46114 35758 46126 35810
rect 44718 35746 44770 35758
rect 6190 35698 6242 35710
rect 8878 35698 8930 35710
rect 1698 35646 1710 35698
rect 1762 35646 1774 35698
rect 6626 35646 6638 35698
rect 6690 35646 6702 35698
rect 7970 35646 7982 35698
rect 8034 35646 8046 35698
rect 6190 35634 6242 35646
rect 8878 35634 8930 35646
rect 9886 35698 9938 35710
rect 9886 35634 9938 35646
rect 10670 35698 10722 35710
rect 10670 35634 10722 35646
rect 11230 35698 11282 35710
rect 11230 35634 11282 35646
rect 12126 35698 12178 35710
rect 12126 35634 12178 35646
rect 12574 35698 12626 35710
rect 12574 35634 12626 35646
rect 12798 35698 12850 35710
rect 12798 35634 12850 35646
rect 13134 35698 13186 35710
rect 13134 35634 13186 35646
rect 14366 35698 14418 35710
rect 14366 35634 14418 35646
rect 16046 35698 16098 35710
rect 20750 35698 20802 35710
rect 23214 35698 23266 35710
rect 17378 35646 17390 35698
rect 17442 35646 17454 35698
rect 21074 35646 21086 35698
rect 21138 35646 21150 35698
rect 22866 35646 22878 35698
rect 22930 35646 22942 35698
rect 16046 35634 16098 35646
rect 20750 35634 20802 35646
rect 23214 35634 23266 35646
rect 23998 35698 24050 35710
rect 23998 35634 24050 35646
rect 26462 35698 26514 35710
rect 26462 35634 26514 35646
rect 27022 35698 27074 35710
rect 27022 35634 27074 35646
rect 27470 35698 27522 35710
rect 30382 35698 30434 35710
rect 31950 35698 32002 35710
rect 39118 35698 39170 35710
rect 41694 35698 41746 35710
rect 28018 35646 28030 35698
rect 28082 35646 28094 35698
rect 28578 35646 28590 35698
rect 28642 35646 28654 35698
rect 31154 35646 31166 35698
rect 31218 35646 31230 35698
rect 34626 35646 34638 35698
rect 34690 35646 34702 35698
rect 38434 35646 38446 35698
rect 38498 35646 38510 35698
rect 41458 35646 41470 35698
rect 41522 35646 41534 35698
rect 27470 35634 27522 35646
rect 30382 35634 30434 35646
rect 31950 35634 32002 35646
rect 39118 35634 39170 35646
rect 41694 35634 41746 35646
rect 41806 35698 41858 35710
rect 41806 35634 41858 35646
rect 42478 35698 42530 35710
rect 42478 35634 42530 35646
rect 43598 35698 43650 35710
rect 45378 35646 45390 35698
rect 45442 35646 45454 35698
rect 43598 35634 43650 35646
rect 5294 35586 5346 35598
rect 15262 35586 15314 35598
rect 20638 35586 20690 35598
rect 4610 35534 4622 35586
rect 4674 35534 4686 35586
rect 11890 35534 11902 35586
rect 11954 35534 11966 35586
rect 20290 35534 20302 35586
rect 20354 35534 20366 35586
rect 5294 35522 5346 35534
rect 15262 35522 15314 35534
rect 20638 35522 20690 35534
rect 24446 35586 24498 35598
rect 24446 35522 24498 35534
rect 25342 35586 25394 35598
rect 25342 35522 25394 35534
rect 25790 35586 25842 35598
rect 25790 35522 25842 35534
rect 26798 35586 26850 35598
rect 26798 35522 26850 35534
rect 27246 35586 27298 35598
rect 27246 35522 27298 35534
rect 29710 35586 29762 35598
rect 31614 35586 31666 35598
rect 39006 35586 39058 35598
rect 30818 35534 30830 35586
rect 30882 35534 30894 35586
rect 33170 35534 33182 35586
rect 33234 35534 33246 35586
rect 35634 35534 35646 35586
rect 35698 35534 35710 35586
rect 37762 35534 37774 35586
rect 37826 35534 37838 35586
rect 29710 35522 29762 35534
rect 31614 35522 31666 35534
rect 39006 35522 39058 35534
rect 40350 35586 40402 35598
rect 40350 35522 40402 35534
rect 41246 35586 41298 35598
rect 41246 35522 41298 35534
rect 42590 35586 42642 35598
rect 42590 35522 42642 35534
rect 42702 35586 42754 35598
rect 48178 35534 48190 35586
rect 48242 35534 48254 35586
rect 42702 35522 42754 35534
rect 11566 35474 11618 35486
rect 11566 35410 11618 35422
rect 13358 35474 13410 35486
rect 13358 35410 13410 35422
rect 15374 35474 15426 35486
rect 15374 35410 15426 35422
rect 1344 35306 48608 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 48608 35306
rect 1344 35220 48608 35254
rect 13358 35138 13410 35150
rect 13358 35074 13410 35086
rect 14814 35138 14866 35150
rect 14814 35074 14866 35086
rect 19518 35138 19570 35150
rect 19518 35074 19570 35086
rect 28478 35138 28530 35150
rect 30494 35138 30546 35150
rect 29698 35086 29710 35138
rect 29762 35086 29774 35138
rect 28478 35074 28530 35086
rect 30494 35074 30546 35086
rect 36990 35138 37042 35150
rect 36990 35074 37042 35086
rect 37326 35138 37378 35150
rect 37326 35074 37378 35086
rect 3726 35026 3778 35038
rect 3726 34962 3778 34974
rect 5742 35026 5794 35038
rect 14254 35026 14306 35038
rect 9874 34974 9886 35026
rect 9938 34974 9950 35026
rect 10882 34974 10894 35026
rect 10946 34974 10958 35026
rect 5742 34962 5794 34974
rect 14254 34962 14306 34974
rect 15150 35026 15202 35038
rect 18734 35026 18786 35038
rect 35982 35026 36034 35038
rect 42478 35026 42530 35038
rect 15922 34974 15934 35026
rect 15986 34974 15998 35026
rect 17826 34974 17838 35026
rect 17890 34974 17902 35026
rect 21298 34974 21310 35026
rect 21362 34974 21374 35026
rect 24322 34974 24334 35026
rect 24386 34974 24398 35026
rect 26450 34974 26462 35026
rect 26514 34974 26526 35026
rect 30930 34974 30942 35026
rect 30994 34974 31006 35026
rect 38658 34974 38670 35026
rect 38722 34974 38734 35026
rect 40786 34974 40798 35026
rect 40850 34974 40862 35026
rect 41234 34974 41246 35026
rect 41298 34974 41310 35026
rect 15150 34962 15202 34974
rect 18734 34962 18786 34974
rect 35982 34962 36034 34974
rect 42478 34962 42530 34974
rect 44158 35026 44210 35038
rect 48178 34974 48190 35026
rect 48242 34974 48254 35026
rect 44158 34962 44210 34974
rect 2606 34914 2658 34926
rect 2606 34850 2658 34862
rect 5630 34914 5682 34926
rect 6414 34914 6466 34926
rect 6178 34862 6190 34914
rect 6242 34862 6254 34914
rect 5630 34850 5682 34862
rect 6414 34850 6466 34862
rect 6750 34914 6802 34926
rect 6750 34850 6802 34862
rect 7646 34914 7698 34926
rect 13806 34914 13858 34926
rect 9650 34862 9662 34914
rect 9714 34862 9726 34914
rect 11666 34862 11678 34914
rect 11730 34862 11742 34914
rect 7646 34850 7698 34862
rect 13806 34850 13858 34862
rect 14030 34914 14082 34926
rect 18174 34914 18226 34926
rect 16258 34862 16270 34914
rect 16322 34862 16334 34914
rect 16594 34862 16606 34914
rect 16658 34862 16670 34914
rect 14030 34850 14082 34862
rect 18174 34850 18226 34862
rect 18622 34914 18674 34926
rect 18622 34850 18674 34862
rect 18846 34914 18898 34926
rect 22318 34914 22370 34926
rect 29150 34914 29202 34926
rect 18846 34850 18898 34862
rect 19406 34858 19458 34870
rect 2942 34802 2994 34814
rect 2942 34738 2994 34750
rect 3166 34802 3218 34814
rect 3166 34738 3218 34750
rect 4174 34802 4226 34814
rect 4174 34738 4226 34750
rect 7310 34802 7362 34814
rect 8766 34802 8818 34814
rect 7858 34750 7870 34802
rect 7922 34750 7934 34802
rect 7310 34738 7362 34750
rect 8766 34738 8818 34750
rect 10334 34802 10386 34814
rect 10334 34738 10386 34750
rect 11006 34802 11058 34814
rect 11006 34738 11058 34750
rect 11230 34802 11282 34814
rect 15374 34802 15426 34814
rect 22866 34862 22878 34914
rect 22930 34862 22942 34914
rect 23538 34862 23550 34914
rect 23602 34862 23614 34914
rect 27346 34862 27358 34914
rect 27410 34862 27422 34914
rect 27570 34862 27582 34914
rect 27634 34862 27646 34914
rect 28242 34862 28254 34914
rect 28306 34862 28318 34914
rect 22318 34850 22370 34862
rect 29150 34850 29202 34862
rect 29374 34914 29426 34926
rect 32734 34914 32786 34926
rect 30370 34862 30382 34914
rect 30434 34862 30446 34914
rect 31378 34862 31390 34914
rect 31442 34862 31454 34914
rect 32386 34862 32398 34914
rect 32450 34862 32462 34914
rect 29374 34850 29426 34862
rect 32734 34850 32786 34862
rect 34302 34914 34354 34926
rect 34302 34850 34354 34862
rect 35198 34914 35250 34926
rect 35198 34850 35250 34862
rect 35310 34914 35362 34926
rect 35310 34850 35362 34862
rect 35870 34914 35922 34926
rect 35870 34850 35922 34862
rect 36206 34914 36258 34926
rect 37986 34862 37998 34914
rect 38050 34862 38062 34914
rect 41794 34862 41806 34914
rect 41858 34862 41870 34914
rect 45266 34862 45278 34914
rect 45330 34862 45342 34914
rect 36206 34850 36258 34862
rect 11890 34750 11902 34802
rect 11954 34750 11966 34802
rect 12562 34750 12574 34802
rect 12626 34750 12638 34802
rect 15698 34750 15710 34802
rect 15762 34750 15774 34802
rect 19406 34794 19458 34806
rect 19966 34802 20018 34814
rect 11230 34738 11282 34750
rect 15374 34738 15426 34750
rect 19966 34738 20018 34750
rect 20078 34802 20130 34814
rect 20078 34738 20130 34750
rect 20526 34802 20578 34814
rect 20526 34738 20578 34750
rect 21422 34802 21474 34814
rect 21422 34738 21474 34750
rect 21646 34802 21698 34814
rect 33406 34802 33458 34814
rect 21970 34750 21982 34802
rect 22034 34750 22046 34802
rect 22642 34750 22654 34802
rect 22706 34750 22718 34802
rect 21646 34738 21698 34750
rect 33406 34738 33458 34750
rect 34414 34802 34466 34814
rect 34414 34738 34466 34750
rect 34974 34802 35026 34814
rect 34974 34738 35026 34750
rect 36318 34802 36370 34814
rect 44046 34802 44098 34814
rect 42914 34750 42926 34802
rect 42978 34750 42990 34802
rect 36318 34738 36370 34750
rect 44046 34738 44098 34750
rect 44270 34802 44322 34814
rect 46050 34750 46062 34802
rect 46114 34750 46126 34802
rect 44270 34738 44322 34750
rect 1822 34690 1874 34702
rect 1822 34626 1874 34638
rect 2382 34690 2434 34702
rect 2382 34626 2434 34638
rect 2718 34690 2770 34702
rect 2718 34626 2770 34638
rect 4622 34690 4674 34702
rect 4622 34626 4674 34638
rect 5182 34690 5234 34702
rect 5182 34626 5234 34638
rect 5854 34690 5906 34702
rect 5854 34626 5906 34638
rect 6638 34690 6690 34702
rect 6638 34626 6690 34638
rect 7422 34690 7474 34702
rect 7422 34626 7474 34638
rect 8206 34690 8258 34702
rect 8206 34626 8258 34638
rect 8878 34690 8930 34702
rect 8878 34626 8930 34638
rect 9102 34690 9154 34702
rect 9102 34626 9154 34638
rect 12238 34690 12290 34702
rect 12238 34626 12290 34638
rect 17390 34690 17442 34702
rect 17390 34626 17442 34638
rect 19518 34690 19570 34702
rect 19518 34626 19570 34638
rect 20302 34690 20354 34702
rect 20302 34626 20354 34638
rect 20638 34690 20690 34702
rect 20638 34626 20690 34638
rect 20862 34690 20914 34702
rect 20862 34626 20914 34638
rect 32846 34690 32898 34702
rect 32846 34626 32898 34638
rect 32958 34690 33010 34702
rect 32958 34626 33010 34638
rect 33854 34690 33906 34702
rect 33854 34626 33906 34638
rect 35422 34690 35474 34702
rect 35422 34626 35474 34638
rect 37214 34690 37266 34702
rect 37214 34626 37266 34638
rect 41246 34690 41298 34702
rect 41246 34626 41298 34638
rect 41358 34690 41410 34702
rect 41358 34626 41410 34638
rect 41582 34690 41634 34702
rect 41582 34626 41634 34638
rect 42590 34690 42642 34702
rect 42590 34626 42642 34638
rect 43262 34690 43314 34702
rect 43262 34626 43314 34638
rect 44942 34690 44994 34702
rect 44942 34626 44994 34638
rect 1344 34522 48608 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 48608 34522
rect 1344 34436 48608 34470
rect 6862 34354 6914 34366
rect 6862 34290 6914 34302
rect 12350 34354 12402 34366
rect 12350 34290 12402 34302
rect 19182 34354 19234 34366
rect 19182 34290 19234 34302
rect 19294 34354 19346 34366
rect 19294 34290 19346 34302
rect 42030 34354 42082 34366
rect 42030 34290 42082 34302
rect 45726 34354 45778 34366
rect 45726 34290 45778 34302
rect 45838 34354 45890 34366
rect 45838 34290 45890 34302
rect 47854 34354 47906 34366
rect 47854 34290 47906 34302
rect 6526 34242 6578 34254
rect 2482 34190 2494 34242
rect 2546 34190 2558 34242
rect 6526 34178 6578 34190
rect 7086 34242 7138 34254
rect 7086 34178 7138 34190
rect 7198 34242 7250 34254
rect 7198 34178 7250 34190
rect 7870 34242 7922 34254
rect 7870 34178 7922 34190
rect 9998 34242 10050 34254
rect 15710 34242 15762 34254
rect 11666 34190 11678 34242
rect 11730 34190 11742 34242
rect 9998 34178 10050 34190
rect 15710 34178 15762 34190
rect 17726 34242 17778 34254
rect 23550 34242 23602 34254
rect 20962 34190 20974 34242
rect 21026 34190 21038 34242
rect 17726 34178 17778 34190
rect 23550 34178 23602 34190
rect 23662 34242 23714 34254
rect 23662 34178 23714 34190
rect 23886 34242 23938 34254
rect 23886 34178 23938 34190
rect 28814 34242 28866 34254
rect 32174 34242 32226 34254
rect 41022 34242 41074 34254
rect 30818 34190 30830 34242
rect 30882 34190 30894 34242
rect 37314 34190 37326 34242
rect 37378 34190 37390 34242
rect 38658 34190 38670 34242
rect 38722 34190 38734 34242
rect 44370 34190 44382 34242
rect 44434 34190 44446 34242
rect 28814 34178 28866 34190
rect 32174 34178 32226 34190
rect 41022 34178 41074 34190
rect 4958 34130 5010 34142
rect 6302 34130 6354 34142
rect 1698 34078 1710 34130
rect 1762 34078 1774 34130
rect 5170 34078 5182 34130
rect 5234 34078 5246 34130
rect 5618 34078 5630 34130
rect 5682 34078 5694 34130
rect 4958 34066 5010 34078
rect 6302 34066 6354 34078
rect 6638 34130 6690 34142
rect 6638 34066 6690 34078
rect 7758 34130 7810 34142
rect 7758 34066 7810 34078
rect 8094 34130 8146 34142
rect 8094 34066 8146 34078
rect 8878 34130 8930 34142
rect 13246 34130 13298 34142
rect 10322 34078 10334 34130
rect 10386 34078 10398 34130
rect 11106 34078 11118 34130
rect 11170 34078 11182 34130
rect 8878 34066 8930 34078
rect 13246 34066 13298 34078
rect 13582 34130 13634 34142
rect 14366 34130 14418 34142
rect 13906 34078 13918 34130
rect 13970 34078 13982 34130
rect 13582 34066 13634 34078
rect 14366 34066 14418 34078
rect 14814 34130 14866 34142
rect 16718 34130 16770 34142
rect 15138 34078 15150 34130
rect 15202 34078 15214 34130
rect 14814 34066 14866 34078
rect 16718 34066 16770 34078
rect 17390 34130 17442 34142
rect 17390 34066 17442 34078
rect 17838 34130 17890 34142
rect 17838 34066 17890 34078
rect 18286 34130 18338 34142
rect 18286 34066 18338 34078
rect 19406 34130 19458 34142
rect 24110 34130 24162 34142
rect 25230 34130 25282 34142
rect 19730 34078 19742 34130
rect 19794 34078 19806 34130
rect 20178 34078 20190 34130
rect 20242 34078 20254 34130
rect 24546 34078 24558 34130
rect 24610 34078 24622 34130
rect 19406 34066 19458 34078
rect 24110 34066 24162 34078
rect 25230 34066 25282 34078
rect 25342 34130 25394 34142
rect 25342 34066 25394 34078
rect 25454 34130 25506 34142
rect 27470 34130 27522 34142
rect 25778 34078 25790 34130
rect 25842 34078 25854 34130
rect 26562 34078 26574 34130
rect 26626 34078 26638 34130
rect 25454 34066 25506 34078
rect 27470 34066 27522 34078
rect 27918 34130 27970 34142
rect 31278 34130 31330 34142
rect 32958 34130 33010 34142
rect 28130 34078 28142 34130
rect 28194 34078 28206 34130
rect 29586 34078 29598 34130
rect 29650 34078 29662 34130
rect 31490 34078 31502 34130
rect 31554 34078 31566 34130
rect 27918 34066 27970 34078
rect 31278 34066 31330 34078
rect 32958 34066 33010 34078
rect 33294 34130 33346 34142
rect 33294 34066 33346 34078
rect 33518 34130 33570 34142
rect 40014 34130 40066 34142
rect 34178 34078 34190 34130
rect 34242 34078 34254 34130
rect 38434 34078 38446 34130
rect 38498 34078 38510 34130
rect 39666 34078 39678 34130
rect 39730 34078 39742 34130
rect 33518 34066 33570 34078
rect 40014 34066 40066 34078
rect 40238 34130 40290 34142
rect 40238 34066 40290 34078
rect 41470 34130 41522 34142
rect 45950 34130 46002 34142
rect 45154 34078 45166 34130
rect 45218 34078 45230 34130
rect 41470 34066 41522 34078
rect 45950 34066 46002 34078
rect 46286 34130 46338 34142
rect 47170 34078 47182 34130
rect 47234 34078 47246 34130
rect 46286 34066 46338 34078
rect 8318 34018 8370 34030
rect 12686 34018 12738 34030
rect 4610 33966 4622 34018
rect 4674 33966 4686 34018
rect 10098 33966 10110 34018
rect 10162 33966 10174 34018
rect 10994 33966 11006 34018
rect 11058 33966 11070 34018
rect 8318 33954 8370 33966
rect 12686 33954 12738 33966
rect 16158 34018 16210 34030
rect 16158 33954 16210 33966
rect 17502 34018 17554 34030
rect 33182 34018 33234 34030
rect 37102 34018 37154 34030
rect 18722 33966 18734 34018
rect 18786 33966 18798 34018
rect 23090 33966 23102 34018
rect 23154 33966 23166 34018
rect 26786 33966 26798 34018
rect 26850 33966 26862 34018
rect 29698 33966 29710 34018
rect 29762 33966 29774 34018
rect 35522 33966 35534 34018
rect 35586 33966 35598 34018
rect 17502 33954 17554 33966
rect 33182 33954 33234 33966
rect 37102 33954 37154 33966
rect 40126 34018 40178 34030
rect 42242 33966 42254 34018
rect 42306 33966 42318 34018
rect 46610 33966 46622 34018
rect 46674 33966 46686 34018
rect 40126 33954 40178 33966
rect 9774 33906 9826 33918
rect 9774 33842 9826 33854
rect 40910 33906 40962 33918
rect 41234 33854 41246 33906
rect 41298 33903 41310 33906
rect 42018 33903 42030 33906
rect 41298 33857 42030 33903
rect 41298 33854 41310 33857
rect 42018 33854 42030 33857
rect 42082 33854 42094 33906
rect 40910 33842 40962 33854
rect 1344 33738 48608 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 48608 33738
rect 1344 33652 48608 33686
rect 4510 33570 4562 33582
rect 4510 33506 4562 33518
rect 6078 33570 6130 33582
rect 6078 33506 6130 33518
rect 7422 33570 7474 33582
rect 7422 33506 7474 33518
rect 12910 33570 12962 33582
rect 12910 33506 12962 33518
rect 28254 33570 28306 33582
rect 36094 33570 36146 33582
rect 31042 33518 31054 33570
rect 31106 33518 31118 33570
rect 28254 33506 28306 33518
rect 36094 33506 36146 33518
rect 46846 33570 46898 33582
rect 46846 33506 46898 33518
rect 3054 33458 3106 33470
rect 3054 33394 3106 33406
rect 4398 33458 4450 33470
rect 27358 33458 27410 33470
rect 7970 33406 7982 33458
rect 8034 33406 8046 33458
rect 10098 33406 10110 33458
rect 10162 33406 10174 33458
rect 14018 33406 14030 33458
rect 14082 33406 14094 33458
rect 15474 33406 15486 33458
rect 15538 33406 15550 33458
rect 17602 33406 17614 33458
rect 17666 33406 17678 33458
rect 18946 33406 18958 33458
rect 19010 33406 19022 33458
rect 4398 33394 4450 33406
rect 27358 33394 27410 33406
rect 27694 33458 27746 33470
rect 27694 33394 27746 33406
rect 29710 33458 29762 33470
rect 35422 33458 35474 33470
rect 30818 33406 30830 33458
rect 30882 33406 30894 33458
rect 32722 33406 32734 33458
rect 32786 33406 32798 33458
rect 34850 33406 34862 33458
rect 34914 33406 34926 33458
rect 29710 33394 29762 33406
rect 35422 33394 35474 33406
rect 37326 33458 37378 33470
rect 44942 33458 44994 33470
rect 40114 33406 40126 33458
rect 40178 33406 40190 33458
rect 42242 33406 42254 33458
rect 42306 33406 42318 33458
rect 37326 33394 37378 33406
rect 44942 33394 44994 33406
rect 3614 33346 3666 33358
rect 11678 33346 11730 33358
rect 19742 33346 19794 33358
rect 27918 33346 27970 33358
rect 7410 33294 7422 33346
rect 7474 33294 7486 33346
rect 10882 33294 10894 33346
rect 10946 33294 10958 33346
rect 12002 33294 12014 33346
rect 12066 33294 12078 33346
rect 12898 33294 12910 33346
rect 12962 33294 12974 33346
rect 14242 33294 14254 33346
rect 14306 33294 14318 33346
rect 18386 33294 18398 33346
rect 18450 33294 18462 33346
rect 19282 33294 19294 33346
rect 19346 33294 19358 33346
rect 22082 33294 22094 33346
rect 22146 33294 22158 33346
rect 22866 33294 22878 33346
rect 22930 33294 22942 33346
rect 24882 33294 24894 33346
rect 24946 33294 24958 33346
rect 25666 33294 25678 33346
rect 25730 33294 25742 33346
rect 3614 33282 3666 33294
rect 11678 33282 11730 33294
rect 19742 33282 19794 33294
rect 27918 33282 27970 33294
rect 29374 33346 29426 33358
rect 38334 33346 38386 33358
rect 30146 33294 30158 33346
rect 30210 33294 30222 33346
rect 30930 33294 30942 33346
rect 30994 33294 31006 33346
rect 32050 33294 32062 33346
rect 32114 33294 32126 33346
rect 36082 33294 36094 33346
rect 36146 33294 36158 33346
rect 37650 33294 37662 33346
rect 37714 33294 37726 33346
rect 29374 33282 29426 33294
rect 38334 33282 38386 33294
rect 38782 33346 38834 33358
rect 43710 33346 43762 33358
rect 47070 33346 47122 33358
rect 39330 33294 39342 33346
rect 39394 33294 39406 33346
rect 45826 33294 45838 33346
rect 45890 33294 45902 33346
rect 38782 33282 38834 33294
rect 43710 33282 43762 33294
rect 47070 33282 47122 33294
rect 47630 33346 47682 33358
rect 47630 33282 47682 33294
rect 47854 33346 47906 33358
rect 47854 33282 47906 33294
rect 1710 33234 1762 33246
rect 1710 33170 1762 33182
rect 1822 33234 1874 33246
rect 1822 33170 1874 33182
rect 2270 33234 2322 33246
rect 2270 33170 2322 33182
rect 3166 33234 3218 33246
rect 3166 33170 3218 33182
rect 4062 33234 4114 33246
rect 4062 33170 4114 33182
rect 5070 33234 5122 33246
rect 7086 33234 7138 33246
rect 5070 33170 5122 33182
rect 6638 33178 6690 33190
rect 2046 33122 2098 33134
rect 2046 33058 2098 33070
rect 2382 33122 2434 33134
rect 2382 33058 2434 33070
rect 2606 33122 2658 33134
rect 2606 33058 2658 33070
rect 2942 33122 2994 33134
rect 2942 33058 2994 33070
rect 3726 33122 3778 33134
rect 3726 33058 3778 33070
rect 3950 33122 4002 33134
rect 3950 33058 4002 33070
rect 4734 33122 4786 33134
rect 4734 33058 4786 33070
rect 4958 33122 5010 33134
rect 4958 33058 5010 33070
rect 5854 33122 5906 33134
rect 5854 33058 5906 33070
rect 5966 33122 6018 33134
rect 5966 33058 6018 33070
rect 6302 33122 6354 33134
rect 6302 33058 6354 33070
rect 6526 33122 6578 33134
rect 7086 33170 7138 33182
rect 12574 33234 12626 33246
rect 12574 33170 12626 33182
rect 14926 33234 14978 33246
rect 26350 33234 26402 33246
rect 23090 33182 23102 33234
rect 23154 33182 23166 33234
rect 24434 33182 24446 33234
rect 24498 33182 24510 33234
rect 14926 33170 14978 33182
rect 26350 33170 26402 33182
rect 29150 33234 29202 33246
rect 29150 33170 29202 33182
rect 35758 33234 35810 33246
rect 35758 33170 35810 33182
rect 36990 33234 37042 33246
rect 36990 33170 37042 33182
rect 37998 33234 38050 33246
rect 37998 33170 38050 33182
rect 43374 33234 43426 33246
rect 43374 33170 43426 33182
rect 43934 33234 43986 33246
rect 43934 33170 43986 33182
rect 44830 33234 44882 33246
rect 44830 33170 44882 33182
rect 46174 33234 46226 33246
rect 46174 33170 46226 33182
rect 47406 33234 47458 33246
rect 47406 33170 47458 33182
rect 47518 33234 47570 33246
rect 47518 33170 47570 33182
rect 6638 33114 6690 33126
rect 11454 33122 11506 33134
rect 6526 33058 6578 33070
rect 11454 33058 11506 33070
rect 11566 33122 11618 33134
rect 11566 33058 11618 33070
rect 13694 33122 13746 33134
rect 13694 33058 13746 33070
rect 20414 33122 20466 33134
rect 26798 33122 26850 33134
rect 20738 33070 20750 33122
rect 20802 33070 20814 33122
rect 21634 33070 21646 33122
rect 21698 33070 21710 33122
rect 20414 33058 20466 33070
rect 26798 33058 26850 33070
rect 37214 33122 37266 33134
rect 37214 33058 37266 33070
rect 37438 33122 37490 33134
rect 37438 33058 37490 33070
rect 38110 33122 38162 33134
rect 38110 33058 38162 33070
rect 38446 33122 38498 33134
rect 38446 33058 38498 33070
rect 38670 33122 38722 33134
rect 38670 33058 38722 33070
rect 43038 33122 43090 33134
rect 43038 33058 43090 33070
rect 43822 33122 43874 33134
rect 43822 33058 43874 33070
rect 45390 33122 45442 33134
rect 45390 33058 45442 33070
rect 46062 33122 46114 33134
rect 46498 33070 46510 33122
rect 46562 33070 46574 33122
rect 46062 33058 46114 33070
rect 1344 32954 48608 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 48608 32954
rect 1344 32868 48608 32902
rect 15374 32786 15426 32798
rect 11890 32734 11902 32786
rect 11954 32734 11966 32786
rect 15374 32722 15426 32734
rect 23214 32786 23266 32798
rect 31502 32786 31554 32798
rect 24098 32734 24110 32786
rect 24162 32734 24174 32786
rect 23214 32722 23266 32734
rect 31502 32722 31554 32734
rect 32510 32786 32562 32798
rect 36318 32786 36370 32798
rect 34962 32734 34974 32786
rect 35026 32734 35038 32786
rect 32510 32722 32562 32734
rect 36318 32722 36370 32734
rect 3054 32674 3106 32686
rect 3054 32610 3106 32622
rect 3838 32674 3890 32686
rect 23438 32674 23490 32686
rect 8194 32622 8206 32674
rect 8258 32622 8270 32674
rect 10098 32622 10110 32674
rect 10162 32622 10174 32674
rect 3838 32610 3890 32622
rect 23438 32610 23490 32622
rect 24446 32674 24498 32686
rect 24446 32610 24498 32622
rect 24558 32674 24610 32686
rect 24558 32610 24610 32622
rect 25230 32674 25282 32686
rect 25230 32610 25282 32622
rect 27022 32674 27074 32686
rect 27022 32610 27074 32622
rect 29598 32674 29650 32686
rect 36430 32674 36482 32686
rect 33506 32622 33518 32674
rect 33570 32622 33582 32674
rect 29598 32610 29650 32622
rect 36430 32610 36482 32622
rect 40910 32674 40962 32686
rect 40910 32610 40962 32622
rect 41470 32674 41522 32686
rect 46050 32622 46062 32674
rect 46114 32622 46126 32674
rect 41470 32610 41522 32622
rect 2046 32562 2098 32574
rect 2046 32498 2098 32510
rect 2270 32562 2322 32574
rect 2270 32498 2322 32510
rect 2494 32562 2546 32574
rect 2494 32498 2546 32510
rect 2830 32562 2882 32574
rect 3614 32562 3666 32574
rect 3378 32510 3390 32562
rect 3442 32510 3454 32562
rect 2830 32498 2882 32510
rect 3614 32498 3666 32510
rect 3950 32562 4002 32574
rect 15262 32562 15314 32574
rect 4946 32510 4958 32562
rect 5010 32510 5022 32562
rect 5730 32510 5742 32562
rect 5794 32510 5806 32562
rect 8978 32510 8990 32562
rect 9042 32510 9054 32562
rect 11330 32510 11342 32562
rect 11394 32510 11406 32562
rect 14466 32510 14478 32562
rect 14530 32510 14542 32562
rect 3950 32498 4002 32510
rect 15262 32498 15314 32510
rect 15598 32562 15650 32574
rect 16830 32562 16882 32574
rect 23774 32562 23826 32574
rect 41134 32562 41186 32574
rect 16370 32510 16382 32562
rect 16434 32510 16446 32562
rect 19730 32510 19742 32562
rect 19794 32510 19806 32562
rect 21298 32510 21310 32562
rect 21362 32510 21374 32562
rect 22418 32510 22430 32562
rect 22482 32510 22494 32562
rect 22642 32510 22654 32562
rect 22706 32510 22718 32562
rect 25666 32510 25678 32562
rect 25730 32510 25742 32562
rect 27234 32510 27246 32562
rect 27298 32510 27310 32562
rect 28690 32510 28702 32562
rect 28754 32510 28766 32562
rect 30594 32510 30606 32562
rect 30658 32510 30670 32562
rect 34850 32510 34862 32562
rect 34914 32510 34926 32562
rect 37090 32510 37102 32562
rect 37154 32510 37166 32562
rect 44706 32510 44718 32562
rect 44770 32510 44782 32562
rect 45378 32510 45390 32562
rect 45442 32510 45454 32562
rect 15598 32498 15650 32510
rect 16830 32498 16882 32510
rect 23774 32498 23826 32510
rect 41134 32498 41186 32510
rect 2382 32450 2434 32462
rect 2382 32386 2434 32398
rect 2942 32450 2994 32462
rect 9998 32450 10050 32462
rect 20638 32450 20690 32462
rect 27806 32450 27858 32462
rect 35982 32450 36034 32462
rect 40238 32450 40290 32462
rect 5058 32398 5070 32450
rect 5122 32398 5134 32450
rect 5618 32398 5630 32450
rect 5682 32398 5694 32450
rect 12562 32398 12574 32450
rect 12626 32398 12638 32450
rect 16034 32398 16046 32450
rect 16098 32398 16110 32450
rect 19170 32398 19182 32450
rect 19234 32398 19246 32450
rect 20850 32398 20862 32450
rect 20914 32398 20926 32450
rect 21634 32398 21646 32450
rect 21698 32398 21710 32450
rect 23090 32398 23102 32450
rect 23154 32398 23166 32450
rect 25554 32398 25566 32450
rect 25618 32398 25630 32450
rect 29250 32398 29262 32450
rect 29314 32398 29326 32450
rect 30706 32398 30718 32450
rect 30770 32398 30782 32450
rect 33170 32398 33182 32450
rect 33234 32398 33246 32450
rect 38210 32398 38222 32450
rect 38274 32398 38286 32450
rect 2942 32386 2994 32398
rect 6066 32342 6078 32394
rect 6130 32342 6142 32394
rect 9998 32386 10050 32398
rect 20638 32386 20690 32398
rect 27806 32386 27858 32398
rect 35982 32386 36034 32398
rect 40238 32386 40290 32398
rect 41358 32450 41410 32462
rect 41906 32398 41918 32450
rect 41970 32398 41982 32450
rect 44034 32398 44046 32450
rect 44098 32398 44110 32450
rect 48178 32398 48190 32450
rect 48242 32398 48254 32450
rect 41358 32386 41410 32398
rect 24558 32338 24610 32350
rect 24558 32274 24610 32286
rect 1344 32170 48608 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 48608 32170
rect 1344 32084 48608 32118
rect 3054 32002 3106 32014
rect 3054 31938 3106 31950
rect 8542 32002 8594 32014
rect 11790 32002 11842 32014
rect 8866 31950 8878 32002
rect 8930 31950 8942 32002
rect 8542 31938 8594 31950
rect 11790 31938 11842 31950
rect 12238 32002 12290 32014
rect 12238 31938 12290 31950
rect 22094 32002 22146 32014
rect 45726 32002 45778 32014
rect 43922 31950 43934 32002
rect 43986 31950 43998 32002
rect 22094 31938 22146 31950
rect 45726 31938 45778 31950
rect 8318 31890 8370 31902
rect 23102 31890 23154 31902
rect 37326 31890 37378 31902
rect 9762 31838 9774 31890
rect 9826 31838 9838 31890
rect 10210 31838 10222 31890
rect 10274 31838 10286 31890
rect 13794 31838 13806 31890
rect 13858 31838 13870 31890
rect 16146 31838 16158 31890
rect 16210 31838 16222 31890
rect 20290 31838 20302 31890
rect 20354 31838 20366 31890
rect 23986 31838 23998 31890
rect 24050 31838 24062 31890
rect 32610 31838 32622 31890
rect 32674 31838 32686 31890
rect 33506 31838 33518 31890
rect 33570 31838 33582 31890
rect 8318 31826 8370 31838
rect 23102 31826 23154 31838
rect 37326 31826 37378 31838
rect 38110 31890 38162 31902
rect 39330 31838 39342 31890
rect 39394 31838 39406 31890
rect 41458 31838 41470 31890
rect 41522 31838 41534 31890
rect 44146 31838 44158 31890
rect 44210 31887 44222 31890
rect 44370 31887 44382 31890
rect 44210 31841 44382 31887
rect 44210 31838 44222 31841
rect 44370 31838 44382 31841
rect 44434 31838 44446 31890
rect 38110 31826 38162 31838
rect 1934 31778 1986 31790
rect 1934 31714 1986 31726
rect 2830 31778 2882 31790
rect 12462 31778 12514 31790
rect 14590 31778 14642 31790
rect 21198 31778 21250 31790
rect 6962 31726 6974 31778
rect 7026 31726 7038 31778
rect 9426 31726 9438 31778
rect 9490 31726 9502 31778
rect 10322 31726 10334 31778
rect 10386 31726 10398 31778
rect 13682 31726 13694 31778
rect 13746 31726 13758 31778
rect 15810 31726 15822 31778
rect 15874 31726 15886 31778
rect 16594 31726 16606 31778
rect 16658 31726 16670 31778
rect 17490 31726 17502 31778
rect 17554 31726 17566 31778
rect 2830 31714 2882 31726
rect 12462 31714 12514 31726
rect 14590 31714 14642 31726
rect 21198 31714 21250 31726
rect 22766 31778 22818 31790
rect 25454 31778 25506 31790
rect 23314 31726 23326 31778
rect 23378 31726 23390 31778
rect 24098 31726 24110 31778
rect 24162 31726 24174 31778
rect 22766 31714 22818 31726
rect 25454 31714 25506 31726
rect 25790 31778 25842 31790
rect 27134 31778 27186 31790
rect 37998 31778 38050 31790
rect 45950 31778 46002 31790
rect 47630 31778 47682 31790
rect 26450 31726 26462 31778
rect 26514 31726 26526 31778
rect 28018 31726 28030 31778
rect 28082 31726 28094 31778
rect 30482 31726 30494 31778
rect 30546 31726 30558 31778
rect 31602 31726 31614 31778
rect 31666 31726 31678 31778
rect 36418 31726 36430 31778
rect 36482 31726 36494 31778
rect 38546 31726 38558 31778
rect 38610 31726 38622 31778
rect 42242 31726 42254 31778
rect 42306 31726 42318 31778
rect 43586 31726 43598 31778
rect 43650 31726 43662 31778
rect 43922 31726 43934 31778
rect 43986 31726 43998 31778
rect 46162 31726 46174 31778
rect 46226 31726 46238 31778
rect 46722 31726 46734 31778
rect 46786 31726 46798 31778
rect 48066 31726 48078 31778
rect 48130 31726 48142 31778
rect 25790 31714 25842 31726
rect 27134 31714 27186 31726
rect 37998 31714 38050 31726
rect 45950 31714 46002 31726
rect 47630 31714 47682 31726
rect 3726 31666 3778 31678
rect 9214 31666 9266 31678
rect 5842 31614 5854 31666
rect 5906 31614 5918 31666
rect 7186 31614 7198 31666
rect 7250 31614 7262 31666
rect 3726 31602 3778 31614
rect 9214 31602 9266 31614
rect 11678 31666 11730 31678
rect 11678 31602 11730 31614
rect 11902 31666 11954 31678
rect 20750 31666 20802 31678
rect 16258 31614 16270 31666
rect 16322 31614 16334 31666
rect 16930 31614 16942 31666
rect 16994 31614 17006 31666
rect 18162 31614 18174 31666
rect 18226 31614 18238 31666
rect 11902 31602 11954 31614
rect 20750 31602 20802 31614
rect 21422 31666 21474 31678
rect 21422 31602 21474 31614
rect 21646 31666 21698 31678
rect 21646 31602 21698 31614
rect 21870 31666 21922 31678
rect 28590 31666 28642 31678
rect 24770 31614 24782 31666
rect 24834 31614 24846 31666
rect 21870 31602 21922 31614
rect 28590 31602 28642 31614
rect 29150 31666 29202 31678
rect 33070 31666 33122 31678
rect 30370 31614 30382 31666
rect 30434 31614 30446 31666
rect 29150 31602 29202 31614
rect 33070 31602 33122 31614
rect 33182 31666 33234 31678
rect 45614 31666 45666 31678
rect 35634 31614 35646 31666
rect 35698 31614 35710 31666
rect 45154 31614 45166 31666
rect 45218 31614 45230 31666
rect 46498 31614 46510 31666
rect 46562 31614 46574 31666
rect 46946 31614 46958 31666
rect 47010 31614 47022 31666
rect 33182 31602 33234 31614
rect 45614 31602 45666 31614
rect 2046 31554 2098 31566
rect 2046 31490 2098 31502
rect 2158 31554 2210 31566
rect 2158 31490 2210 31502
rect 2382 31554 2434 31566
rect 3838 31554 3890 31566
rect 3378 31502 3390 31554
rect 3442 31502 3454 31554
rect 2382 31490 2434 31502
rect 3838 31490 3890 31502
rect 3950 31554 4002 31566
rect 3950 31490 4002 31502
rect 4174 31554 4226 31566
rect 5070 31554 5122 31566
rect 11342 31554 11394 31566
rect 4722 31502 4734 31554
rect 4786 31502 4798 31554
rect 5954 31502 5966 31554
rect 6018 31502 6030 31554
rect 4174 31490 4226 31502
rect 5070 31490 5122 31502
rect 11342 31490 11394 31502
rect 15262 31554 15314 31566
rect 15262 31490 15314 31502
rect 20638 31554 20690 31566
rect 20638 31490 20690 31502
rect 22206 31554 22258 31566
rect 22206 31490 22258 31502
rect 22430 31554 22482 31566
rect 22430 31490 22482 31502
rect 25566 31554 25618 31566
rect 25566 31490 25618 31502
rect 29262 31554 29314 31566
rect 29262 31490 29314 31502
rect 29486 31554 29538 31566
rect 29486 31490 29538 31502
rect 32846 31554 32898 31566
rect 32846 31490 32898 31502
rect 37438 31554 37490 31566
rect 37438 31490 37490 31502
rect 37550 31554 37602 31566
rect 37550 31490 37602 31502
rect 38222 31554 38274 31566
rect 38222 31490 38274 31502
rect 39006 31554 39058 31566
rect 39006 31490 39058 31502
rect 42702 31554 42754 31566
rect 42702 31490 42754 31502
rect 44830 31554 44882 31566
rect 44830 31490 44882 31502
rect 1344 31386 48608 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 48608 31386
rect 1344 31300 48608 31334
rect 7198 31218 7250 31230
rect 6850 31166 6862 31218
rect 6914 31166 6926 31218
rect 7198 31154 7250 31166
rect 8766 31218 8818 31230
rect 8766 31154 8818 31166
rect 17390 31218 17442 31230
rect 17390 31154 17442 31166
rect 22766 31218 22818 31230
rect 28254 31218 28306 31230
rect 33966 31218 34018 31230
rect 25666 31166 25678 31218
rect 25730 31166 25742 31218
rect 30594 31166 30606 31218
rect 30658 31166 30670 31218
rect 22766 31154 22818 31166
rect 28254 31154 28306 31166
rect 33966 31154 34018 31166
rect 34526 31218 34578 31230
rect 34526 31154 34578 31166
rect 34638 31218 34690 31230
rect 34638 31154 34690 31166
rect 44270 31218 44322 31230
rect 44270 31154 44322 31166
rect 46174 31218 46226 31230
rect 46174 31154 46226 31166
rect 48302 31218 48354 31230
rect 48302 31154 48354 31166
rect 16158 31106 16210 31118
rect 2482 31054 2494 31106
rect 2546 31054 2558 31106
rect 7858 31054 7870 31106
rect 7922 31054 7934 31106
rect 8194 31054 8206 31106
rect 8258 31054 8270 31106
rect 16158 31042 16210 31054
rect 22094 31106 22146 31118
rect 28030 31106 28082 31118
rect 33070 31106 33122 31118
rect 22418 31054 22430 31106
rect 22482 31054 22494 31106
rect 30146 31054 30158 31106
rect 30210 31054 30222 31106
rect 31154 31054 31166 31106
rect 31218 31054 31230 31106
rect 22094 31042 22146 31054
rect 28030 31042 28082 31054
rect 33070 31042 33122 31054
rect 33294 31106 33346 31118
rect 33294 31042 33346 31054
rect 34750 31106 34802 31118
rect 38558 31106 38610 31118
rect 37202 31054 37214 31106
rect 37266 31054 37278 31106
rect 34750 31042 34802 31054
rect 38558 31042 38610 31054
rect 40238 31106 40290 31118
rect 40238 31042 40290 31054
rect 44718 31106 44770 31118
rect 44718 31042 44770 31054
rect 45614 31106 45666 31118
rect 45614 31042 45666 31054
rect 45950 31106 46002 31118
rect 45950 31042 46002 31054
rect 46398 31106 46450 31118
rect 46398 31042 46450 31054
rect 47406 31106 47458 31118
rect 47406 31042 47458 31054
rect 6526 30994 6578 31006
rect 15822 30994 15874 31006
rect 17950 30994 18002 31006
rect 26014 30994 26066 31006
rect 27470 30994 27522 31006
rect 1698 30942 1710 30994
rect 1762 30942 1774 30994
rect 5170 30942 5182 30994
rect 5234 30942 5246 30994
rect 6066 30942 6078 30994
rect 6130 30942 6142 30994
rect 9650 30942 9662 30994
rect 9714 30942 9726 30994
rect 15362 30942 15374 30994
rect 15426 30942 15438 30994
rect 16594 30942 16606 30994
rect 16658 30942 16670 30994
rect 17602 30942 17614 30994
rect 17666 30942 17678 30994
rect 18722 30942 18734 30994
rect 18786 30942 18798 30994
rect 21522 30942 21534 30994
rect 21586 30942 21598 30994
rect 24098 30942 24110 30994
rect 24162 30942 24174 30994
rect 26786 30942 26798 30994
rect 26850 30942 26862 30994
rect 6526 30930 6578 30942
rect 15822 30930 15874 30942
rect 17950 30930 18002 30942
rect 26014 30930 26066 30942
rect 27470 30930 27522 30942
rect 28254 30994 28306 31006
rect 28254 30930 28306 30942
rect 28478 30994 28530 31006
rect 33182 30994 33234 31006
rect 29698 30942 29710 30994
rect 29762 30942 29774 30994
rect 30818 30942 30830 30994
rect 30882 30942 30894 30994
rect 31714 30942 31726 30994
rect 31778 30942 31790 30994
rect 32610 30942 32622 30994
rect 32674 30942 32686 30994
rect 28478 30930 28530 30942
rect 33182 30930 33234 30942
rect 33742 30994 33794 31006
rect 38334 30994 38386 31006
rect 39342 30994 39394 31006
rect 44158 30994 44210 31006
rect 45054 30994 45106 31006
rect 37874 30942 37886 30994
rect 37938 30942 37950 30994
rect 38882 30942 38894 30994
rect 38946 30942 38958 30994
rect 39554 30942 39566 30994
rect 39618 30942 39630 30994
rect 41458 30942 41470 30994
rect 41522 30942 41534 30994
rect 44370 30942 44382 30994
rect 44434 30942 44446 30994
rect 33742 30930 33794 30942
rect 38334 30930 38386 30942
rect 39342 30930 39394 30942
rect 44158 30930 44210 30942
rect 45054 30930 45106 30942
rect 45278 30994 45330 31006
rect 45278 30930 45330 30942
rect 46510 30994 46562 31006
rect 46510 30930 46562 30942
rect 23214 30882 23266 30894
rect 25342 30882 25394 30894
rect 29486 30882 29538 30894
rect 33854 30882 33906 30894
rect 38446 30882 38498 30894
rect 44830 30882 44882 30894
rect 4610 30830 4622 30882
rect 4674 30830 4686 30882
rect 5282 30830 5294 30882
rect 5346 30830 5358 30882
rect 10322 30830 10334 30882
rect 10386 30830 10398 30882
rect 12450 30830 12462 30882
rect 12514 30830 12526 30882
rect 13234 30830 13246 30882
rect 13298 30830 13310 30882
rect 20066 30830 20078 30882
rect 20130 30830 20142 30882
rect 21186 30830 21198 30882
rect 21250 30830 21262 30882
rect 23762 30830 23774 30882
rect 23826 30830 23838 30882
rect 26674 30830 26686 30882
rect 26738 30830 26750 30882
rect 31826 30830 31838 30882
rect 31890 30830 31902 30882
rect 35074 30830 35086 30882
rect 35138 30830 35150 30882
rect 42354 30830 42366 30882
rect 42418 30830 42430 30882
rect 23214 30818 23266 30830
rect 25342 30818 25394 30830
rect 29486 30818 29538 30830
rect 33854 30818 33906 30830
rect 38446 30818 38498 30830
rect 44830 30818 44882 30830
rect 46958 30882 47010 30894
rect 46958 30818 47010 30830
rect 8430 30770 8482 30782
rect 8430 30706 8482 30718
rect 17278 30770 17330 30782
rect 43934 30770 43986 30782
rect 24322 30718 24334 30770
rect 24386 30718 24398 30770
rect 17278 30706 17330 30718
rect 43934 30706 43986 30718
rect 1344 30602 48608 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 48608 30602
rect 1344 30516 48608 30550
rect 7646 30434 7698 30446
rect 7646 30370 7698 30382
rect 7982 30434 8034 30446
rect 20414 30434 20466 30446
rect 17154 30382 17166 30434
rect 17218 30382 17230 30434
rect 7982 30370 8034 30382
rect 20414 30370 20466 30382
rect 20750 30434 20802 30446
rect 24446 30434 24498 30446
rect 46062 30434 46114 30446
rect 22082 30382 22094 30434
rect 22146 30431 22158 30434
rect 22306 30431 22318 30434
rect 22146 30385 22318 30431
rect 22146 30382 22158 30385
rect 22306 30382 22318 30385
rect 22370 30382 22382 30434
rect 25218 30382 25230 30434
rect 25282 30382 25294 30434
rect 43250 30382 43262 30434
rect 43314 30382 43326 30434
rect 20750 30370 20802 30382
rect 24446 30370 24498 30382
rect 46062 30370 46114 30382
rect 46398 30434 46450 30446
rect 46398 30370 46450 30382
rect 1934 30322 1986 30334
rect 3390 30322 3442 30334
rect 13582 30322 13634 30334
rect 19854 30322 19906 30334
rect 3042 30270 3054 30322
rect 3106 30270 3118 30322
rect 4946 30270 4958 30322
rect 5010 30270 5022 30322
rect 12338 30270 12350 30322
rect 12402 30270 12414 30322
rect 16594 30270 16606 30322
rect 16658 30270 16670 30322
rect 1934 30258 1986 30270
rect 3390 30258 3442 30270
rect 13582 30258 13634 30270
rect 19854 30258 19906 30270
rect 20302 30322 20354 30334
rect 20302 30258 20354 30270
rect 21422 30322 21474 30334
rect 21422 30258 21474 30270
rect 24782 30322 24834 30334
rect 24782 30258 24834 30270
rect 28030 30322 28082 30334
rect 31378 30270 31390 30322
rect 31442 30270 31454 30322
rect 31938 30270 31950 30322
rect 32002 30270 32014 30322
rect 39890 30270 39902 30322
rect 39954 30270 39966 30322
rect 42242 30270 42254 30322
rect 42306 30270 42318 30322
rect 45266 30270 45278 30322
rect 45330 30270 45342 30322
rect 28030 30258 28082 30270
rect 7086 30210 7138 30222
rect 2930 30158 2942 30210
rect 2994 30158 3006 30210
rect 7086 30146 7138 30158
rect 7310 30210 7362 30222
rect 9214 30210 9266 30222
rect 8642 30158 8654 30210
rect 8706 30158 8718 30210
rect 7310 30146 7362 30158
rect 9214 30146 9266 30158
rect 9662 30210 9714 30222
rect 9662 30146 9714 30158
rect 9886 30210 9938 30222
rect 9886 30146 9938 30158
rect 10334 30210 10386 30222
rect 10334 30146 10386 30158
rect 10782 30210 10834 30222
rect 18062 30210 18114 30222
rect 12114 30158 12126 30210
rect 12178 30158 12190 30210
rect 12898 30158 12910 30210
rect 12962 30158 12974 30210
rect 14466 30158 14478 30210
rect 14530 30158 14542 30210
rect 15922 30158 15934 30210
rect 15986 30158 15998 30210
rect 16482 30158 16494 30210
rect 16546 30158 16558 30210
rect 17826 30158 17838 30210
rect 17890 30158 17902 30210
rect 10782 30146 10834 30158
rect 18062 30146 18114 30158
rect 20638 30210 20690 30222
rect 20638 30146 20690 30158
rect 21310 30210 21362 30222
rect 21310 30146 21362 30158
rect 21534 30210 21586 30222
rect 21534 30146 21586 30158
rect 21982 30210 22034 30222
rect 25566 30210 25618 30222
rect 23202 30158 23214 30210
rect 23266 30158 23278 30210
rect 23538 30158 23550 30210
rect 23602 30158 23614 30210
rect 21982 30146 22034 30158
rect 25566 30146 25618 30158
rect 25790 30210 25842 30222
rect 25790 30146 25842 30158
rect 26014 30210 26066 30222
rect 26014 30146 26066 30158
rect 27134 30210 27186 30222
rect 33294 30210 33346 30222
rect 27458 30158 27470 30210
rect 27522 30158 27534 30210
rect 30370 30158 30382 30210
rect 30434 30158 30446 30210
rect 30930 30158 30942 30210
rect 30994 30158 31006 30210
rect 32050 30158 32062 30210
rect 32114 30158 32126 30210
rect 32722 30158 32734 30210
rect 32786 30158 32798 30210
rect 27134 30146 27186 30158
rect 33294 30146 33346 30158
rect 34750 30210 34802 30222
rect 34750 30146 34802 30158
rect 34974 30210 35026 30222
rect 34974 30146 35026 30158
rect 35758 30210 35810 30222
rect 43486 30210 43538 30222
rect 37090 30158 37102 30210
rect 37154 30158 37166 30210
rect 40786 30158 40798 30210
rect 40850 30158 40862 30210
rect 35758 30146 35810 30158
rect 43486 30146 43538 30158
rect 43934 30210 43986 30222
rect 45614 30210 45666 30222
rect 45154 30158 45166 30210
rect 45218 30158 45230 30210
rect 43934 30146 43986 30158
rect 45614 30146 45666 30158
rect 46286 30210 46338 30222
rect 47070 30210 47122 30222
rect 46834 30158 46846 30210
rect 46898 30158 46910 30210
rect 47618 30158 47630 30210
rect 47682 30158 47694 30210
rect 46286 30146 46338 30158
rect 47070 30146 47122 30158
rect 1822 30098 1874 30110
rect 1822 30034 1874 30046
rect 2046 30098 2098 30110
rect 2046 30034 2098 30046
rect 3838 30098 3890 30110
rect 3838 30034 3890 30046
rect 4062 30098 4114 30110
rect 10222 30098 10274 30110
rect 6402 30046 6414 30098
rect 6466 30046 6478 30098
rect 6962 30046 6974 30098
rect 7026 30046 7038 30098
rect 8754 30046 8766 30098
rect 8818 30046 8830 30098
rect 4062 30034 4114 30046
rect 10222 30034 10274 30046
rect 10670 30098 10722 30110
rect 15710 30098 15762 30110
rect 11890 30046 11902 30098
rect 11954 30046 11966 30098
rect 14914 30046 14926 30098
rect 14978 30046 14990 30098
rect 10670 30034 10722 30046
rect 15710 30034 15762 30046
rect 17726 30098 17778 30110
rect 17726 30034 17778 30046
rect 18846 30098 18898 30110
rect 18846 30034 18898 30046
rect 19406 30098 19458 30110
rect 24558 30098 24610 30110
rect 22754 30046 22766 30098
rect 22818 30046 22830 30098
rect 19406 30034 19458 30046
rect 24558 30034 24610 30046
rect 26350 30098 26402 30110
rect 26350 30034 26402 30046
rect 29934 30098 29986 30110
rect 45950 30098 46002 30110
rect 31042 30046 31054 30098
rect 31106 30046 31118 30098
rect 31938 30046 31950 30098
rect 32002 30046 32014 30098
rect 37762 30046 37774 30098
rect 37826 30046 37838 30098
rect 45042 30046 45054 30098
rect 45106 30046 45118 30098
rect 29934 30034 29986 30046
rect 45950 30034 46002 30046
rect 47182 30098 47234 30110
rect 47182 30034 47234 30046
rect 3950 29986 4002 29998
rect 3950 29922 4002 29934
rect 4510 29986 4562 29998
rect 4510 29922 4562 29934
rect 5854 29986 5906 29998
rect 5854 29922 5906 29934
rect 9550 29986 9602 29998
rect 14142 29986 14194 29998
rect 22430 29986 22482 29998
rect 26238 29986 26290 29998
rect 11218 29934 11230 29986
rect 11282 29934 11294 29986
rect 15586 29934 15598 29986
rect 15650 29934 15662 29986
rect 23762 29934 23774 29986
rect 23826 29934 23838 29986
rect 23986 29934 23998 29986
rect 24050 29934 24062 29986
rect 9550 29922 9602 29934
rect 14142 29922 14194 29934
rect 22430 29922 22482 29934
rect 26238 29922 26290 29934
rect 28590 29986 28642 29998
rect 28590 29922 28642 29934
rect 29374 29986 29426 29998
rect 29374 29922 29426 29934
rect 29598 29986 29650 29998
rect 29598 29922 29650 29934
rect 29822 29986 29874 29998
rect 29822 29922 29874 29934
rect 33630 29986 33682 29998
rect 36542 29986 36594 29998
rect 35298 29934 35310 29986
rect 35362 29934 35374 29986
rect 33630 29922 33682 29934
rect 36542 29922 36594 29934
rect 45390 29986 45442 29998
rect 45390 29922 45442 29934
rect 48078 29986 48130 29998
rect 48078 29922 48130 29934
rect 1344 29818 48608 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 48608 29818
rect 1344 29732 48608 29766
rect 6526 29650 6578 29662
rect 6526 29586 6578 29598
rect 11790 29650 11842 29662
rect 18062 29650 18114 29662
rect 16594 29598 16606 29650
rect 16658 29598 16670 29650
rect 11790 29586 11842 29598
rect 18062 29586 18114 29598
rect 20862 29650 20914 29662
rect 20862 29586 20914 29598
rect 23326 29650 23378 29662
rect 23326 29586 23378 29598
rect 23438 29650 23490 29662
rect 23438 29586 23490 29598
rect 24110 29650 24162 29662
rect 24110 29586 24162 29598
rect 24222 29650 24274 29662
rect 24222 29586 24274 29598
rect 24334 29650 24386 29662
rect 24334 29586 24386 29598
rect 25790 29650 25842 29662
rect 25790 29586 25842 29598
rect 27134 29650 27186 29662
rect 32286 29650 32338 29662
rect 37438 29650 37490 29662
rect 28466 29598 28478 29650
rect 28530 29598 28542 29650
rect 35858 29598 35870 29650
rect 35922 29598 35934 29650
rect 27134 29586 27186 29598
rect 32286 29586 32338 29598
rect 37438 29586 37490 29598
rect 46846 29650 46898 29662
rect 46846 29586 46898 29598
rect 2494 29538 2546 29550
rect 4846 29538 4898 29550
rect 4162 29486 4174 29538
rect 4226 29486 4238 29538
rect 2494 29474 2546 29486
rect 4846 29474 4898 29486
rect 5070 29538 5122 29550
rect 5070 29474 5122 29486
rect 5294 29538 5346 29550
rect 5294 29474 5346 29486
rect 6974 29538 7026 29550
rect 6974 29474 7026 29486
rect 8430 29538 8482 29550
rect 10222 29538 10274 29550
rect 17950 29538 18002 29550
rect 9874 29486 9886 29538
rect 9938 29486 9950 29538
rect 13570 29486 13582 29538
rect 13634 29486 13646 29538
rect 8430 29474 8482 29486
rect 10222 29474 10274 29486
rect 17950 29474 18002 29486
rect 18846 29538 18898 29550
rect 29150 29538 29202 29550
rect 34078 29538 34130 29550
rect 37774 29538 37826 29550
rect 42814 29538 42866 29550
rect 21186 29486 21198 29538
rect 21250 29486 21262 29538
rect 30146 29486 30158 29538
rect 30210 29486 30222 29538
rect 31602 29486 31614 29538
rect 31666 29486 31678 29538
rect 36754 29486 36766 29538
rect 36818 29486 36830 29538
rect 40002 29486 40014 29538
rect 40066 29486 40078 29538
rect 41122 29486 41134 29538
rect 41186 29486 41198 29538
rect 44146 29486 44158 29538
rect 44210 29486 44222 29538
rect 18846 29474 18898 29486
rect 29150 29474 29202 29486
rect 34078 29474 34130 29486
rect 37774 29474 37826 29486
rect 42814 29474 42866 29486
rect 2046 29426 2098 29438
rect 2046 29362 2098 29374
rect 2158 29426 2210 29438
rect 6078 29426 6130 29438
rect 2818 29374 2830 29426
rect 2882 29374 2894 29426
rect 3602 29374 3614 29426
rect 3666 29374 3678 29426
rect 2158 29362 2210 29374
rect 6078 29362 6130 29374
rect 6302 29426 6354 29438
rect 6302 29362 6354 29374
rect 6750 29426 6802 29438
rect 8878 29426 8930 29438
rect 7970 29374 7982 29426
rect 8034 29374 8046 29426
rect 6750 29362 6802 29374
rect 8878 29362 8930 29374
rect 9550 29426 9602 29438
rect 9550 29362 9602 29374
rect 10558 29426 10610 29438
rect 15374 29426 15426 29438
rect 17390 29426 17442 29438
rect 12338 29374 12350 29426
rect 12402 29374 12414 29426
rect 12674 29374 12686 29426
rect 12738 29374 12750 29426
rect 14354 29374 14366 29426
rect 14418 29374 14430 29426
rect 16370 29374 16382 29426
rect 16434 29374 16446 29426
rect 10558 29362 10610 29374
rect 15374 29362 15426 29374
rect 17390 29362 17442 29374
rect 17838 29426 17890 29438
rect 17838 29362 17890 29374
rect 18958 29426 19010 29438
rect 18958 29362 19010 29374
rect 19070 29426 19122 29438
rect 23214 29426 23266 29438
rect 24782 29426 24834 29438
rect 19842 29374 19854 29426
rect 19906 29374 19918 29426
rect 20178 29374 20190 29426
rect 20242 29374 20254 29426
rect 21298 29374 21310 29426
rect 21362 29374 21374 29426
rect 22306 29374 22318 29426
rect 22370 29374 22382 29426
rect 23762 29374 23774 29426
rect 23826 29374 23838 29426
rect 19070 29362 19122 29374
rect 23214 29362 23266 29374
rect 24782 29362 24834 29374
rect 25678 29426 25730 29438
rect 25678 29362 25730 29374
rect 25902 29426 25954 29438
rect 27918 29426 27970 29438
rect 26226 29374 26238 29426
rect 26290 29374 26302 29426
rect 25902 29362 25954 29374
rect 27918 29362 27970 29374
rect 28814 29426 28866 29438
rect 28814 29362 28866 29374
rect 33182 29426 33234 29438
rect 34526 29426 34578 29438
rect 37214 29426 37266 29438
rect 33618 29374 33630 29426
rect 33682 29374 33694 29426
rect 34738 29374 34750 29426
rect 34802 29374 34814 29426
rect 35746 29374 35758 29426
rect 35810 29374 35822 29426
rect 36306 29374 36318 29426
rect 36370 29374 36382 29426
rect 33182 29362 33234 29374
rect 34526 29362 34578 29374
rect 37214 29362 37266 29374
rect 37438 29426 37490 29438
rect 46622 29426 46674 29438
rect 38770 29374 38782 29426
rect 38834 29374 38846 29426
rect 41234 29374 41246 29426
rect 41298 29374 41310 29426
rect 41906 29374 41918 29426
rect 41970 29374 41982 29426
rect 43362 29374 43374 29426
rect 43426 29374 43438 29426
rect 37438 29362 37490 29374
rect 46622 29362 46674 29374
rect 47070 29426 47122 29438
rect 47070 29362 47122 29374
rect 47294 29426 47346 29438
rect 47294 29362 47346 29374
rect 2382 29314 2434 29326
rect 21758 29314 21810 29326
rect 3714 29262 3726 29314
rect 3778 29262 3790 29314
rect 20402 29262 20414 29314
rect 20466 29262 20478 29314
rect 2382 29250 2434 29262
rect 21758 29250 21810 29262
rect 21870 29314 21922 29326
rect 21870 29250 21922 29262
rect 25342 29314 25394 29326
rect 25342 29250 25394 29262
rect 26574 29314 26626 29326
rect 26574 29250 26626 29262
rect 27582 29314 27634 29326
rect 27582 29250 27634 29262
rect 28142 29314 28194 29326
rect 31838 29314 31890 29326
rect 29698 29262 29710 29314
rect 29762 29262 29774 29314
rect 28142 29250 28194 29262
rect 31838 29250 31890 29262
rect 35422 29314 35474 29326
rect 35422 29250 35474 29262
rect 38110 29314 38162 29326
rect 42702 29314 42754 29326
rect 47854 29314 47906 29326
rect 40226 29262 40238 29314
rect 40290 29262 40302 29314
rect 41682 29262 41694 29314
rect 41746 29262 41758 29314
rect 46274 29262 46286 29314
rect 46338 29262 46350 29314
rect 38110 29250 38162 29262
rect 42702 29250 42754 29262
rect 47854 29250 47906 29262
rect 48190 29314 48242 29326
rect 48190 29250 48242 29262
rect 42590 29202 42642 29214
rect 5618 29150 5630 29202
rect 5682 29150 5694 29202
rect 7186 29150 7198 29202
rect 7250 29150 7262 29202
rect 18386 29150 18398 29202
rect 18450 29150 18462 29202
rect 47394 29150 47406 29202
rect 47458 29199 47470 29202
rect 48066 29199 48078 29202
rect 47458 29153 48078 29199
rect 47458 29150 47470 29153
rect 48066 29150 48078 29153
rect 48130 29150 48142 29202
rect 42590 29138 42642 29150
rect 1344 29034 48608 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 48608 29034
rect 1344 28948 48608 28982
rect 4846 28866 4898 28878
rect 4498 28814 4510 28866
rect 4562 28814 4574 28866
rect 4846 28802 4898 28814
rect 9438 28866 9490 28878
rect 9438 28802 9490 28814
rect 12910 28866 12962 28878
rect 12910 28802 12962 28814
rect 20862 28866 20914 28878
rect 20862 28802 20914 28814
rect 21982 28866 22034 28878
rect 30830 28866 30882 28878
rect 22306 28814 22318 28866
rect 22370 28814 22382 28866
rect 29362 28814 29374 28866
rect 29426 28814 29438 28866
rect 21982 28802 22034 28814
rect 30830 28802 30882 28814
rect 34750 28866 34802 28878
rect 34750 28802 34802 28814
rect 8430 28754 8482 28766
rect 13582 28754 13634 28766
rect 19966 28754 20018 28766
rect 1810 28702 1822 28754
rect 1874 28702 1886 28754
rect 10098 28702 10110 28754
rect 10162 28702 10174 28754
rect 16258 28702 16270 28754
rect 16322 28702 16334 28754
rect 18050 28702 18062 28754
rect 18114 28702 18126 28754
rect 8430 28690 8482 28702
rect 13582 28690 13634 28702
rect 19966 28690 20018 28702
rect 21422 28754 21474 28766
rect 33742 28754 33794 28766
rect 26226 28702 26238 28754
rect 26290 28702 26302 28754
rect 28466 28702 28478 28754
rect 28530 28702 28542 28754
rect 29474 28702 29486 28754
rect 29538 28702 29550 28754
rect 31602 28702 31614 28754
rect 31666 28702 31678 28754
rect 32834 28702 32846 28754
rect 32898 28702 32910 28754
rect 21422 28690 21474 28702
rect 33742 28690 33794 28702
rect 34190 28754 34242 28766
rect 34190 28690 34242 28702
rect 34414 28754 34466 28766
rect 34414 28690 34466 28702
rect 36430 28754 36482 28766
rect 36430 28690 36482 28702
rect 38110 28754 38162 28766
rect 43934 28754 43986 28766
rect 41346 28702 41358 28754
rect 41410 28702 41422 28754
rect 46050 28702 46062 28754
rect 46114 28702 46126 28754
rect 48178 28702 48190 28754
rect 48242 28702 48254 28754
rect 38110 28690 38162 28702
rect 43934 28690 43986 28702
rect 5070 28642 5122 28654
rect 3490 28590 3502 28642
rect 3554 28590 3566 28642
rect 5070 28578 5122 28590
rect 5854 28642 5906 28654
rect 21758 28642 21810 28654
rect 6066 28590 6078 28642
rect 6130 28590 6142 28642
rect 6962 28590 6974 28642
rect 7026 28590 7038 28642
rect 8530 28590 8542 28642
rect 8594 28590 8606 28642
rect 9202 28590 9214 28642
rect 9266 28590 9278 28642
rect 11666 28590 11678 28642
rect 11730 28590 11742 28642
rect 13906 28590 13918 28642
rect 13970 28590 13982 28642
rect 14354 28590 14366 28642
rect 14418 28590 14430 28642
rect 17378 28590 17390 28642
rect 17442 28590 17454 28642
rect 18386 28590 18398 28642
rect 18450 28590 18462 28642
rect 5854 28578 5906 28590
rect 21758 28578 21810 28590
rect 22654 28642 22706 28654
rect 26462 28642 26514 28654
rect 23426 28590 23438 28642
rect 23490 28590 23502 28642
rect 24098 28590 24110 28642
rect 24162 28590 24174 28642
rect 22654 28578 22706 28590
rect 26462 28578 26514 28590
rect 26686 28642 26738 28654
rect 26686 28578 26738 28590
rect 27022 28642 27074 28654
rect 27022 28578 27074 28590
rect 27806 28642 27858 28654
rect 27806 28578 27858 28590
rect 28142 28642 28194 28654
rect 28142 28578 28194 28590
rect 31054 28642 31106 28654
rect 32398 28642 32450 28654
rect 35310 28642 35362 28654
rect 31490 28590 31502 28642
rect 31554 28590 31566 28642
rect 33058 28590 33070 28642
rect 33122 28590 33134 28642
rect 31054 28578 31106 28590
rect 32398 28578 32450 28590
rect 35310 28578 35362 28590
rect 35646 28642 35698 28654
rect 35646 28578 35698 28590
rect 35870 28642 35922 28654
rect 35870 28578 35922 28590
rect 37102 28642 37154 28654
rect 37102 28578 37154 28590
rect 37662 28642 37714 28654
rect 41694 28642 41746 28654
rect 38434 28590 38446 28642
rect 38498 28590 38510 28642
rect 37662 28578 37714 28590
rect 41694 28578 41746 28590
rect 43262 28642 43314 28654
rect 43262 28578 43314 28590
rect 44046 28642 44098 28654
rect 44046 28578 44098 28590
rect 44942 28642 44994 28654
rect 45378 28590 45390 28642
rect 45442 28590 45454 28642
rect 44942 28578 44994 28590
rect 19406 28530 19458 28542
rect 2370 28478 2382 28530
rect 2434 28478 2446 28530
rect 7074 28478 7086 28530
rect 7138 28478 7150 28530
rect 10658 28478 10670 28530
rect 10722 28478 10734 28530
rect 17042 28478 17054 28530
rect 17106 28478 17118 28530
rect 19406 28466 19458 28478
rect 20302 28530 20354 28542
rect 26910 28530 26962 28542
rect 22978 28478 22990 28530
rect 23042 28478 23054 28530
rect 20302 28466 20354 28478
rect 26910 28466 26962 28478
rect 29150 28530 29202 28542
rect 29150 28466 29202 28478
rect 36990 28530 37042 28542
rect 41918 28530 41970 28542
rect 39218 28478 39230 28530
rect 39282 28478 39294 28530
rect 36990 28466 37042 28478
rect 41918 28466 41970 28478
rect 42030 28530 42082 28542
rect 42030 28466 42082 28478
rect 42702 28530 42754 28542
rect 42702 28466 42754 28478
rect 42926 28530 42978 28542
rect 43586 28478 43598 28530
rect 43650 28478 43662 28530
rect 42926 28466 42978 28478
rect 19070 28418 19122 28430
rect 3826 28366 3838 28418
rect 3890 28366 3902 28418
rect 6178 28366 6190 28418
rect 6242 28366 6254 28418
rect 6962 28366 6974 28418
rect 7026 28366 7038 28418
rect 19070 28354 19122 28366
rect 20526 28418 20578 28430
rect 20526 28354 20578 28366
rect 20750 28418 20802 28430
rect 20750 28354 20802 28366
rect 28366 28418 28418 28430
rect 28366 28354 28418 28366
rect 35534 28418 35586 28430
rect 35534 28354 35586 28366
rect 37214 28418 37266 28430
rect 37214 28354 37266 28366
rect 42814 28418 42866 28430
rect 42814 28354 42866 28366
rect 1344 28250 48608 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 48608 28250
rect 1344 28164 48608 28198
rect 5294 28082 5346 28094
rect 9886 28082 9938 28094
rect 13806 28082 13858 28094
rect 5954 28030 5966 28082
rect 6018 28030 6030 28082
rect 10210 28030 10222 28082
rect 10274 28030 10286 28082
rect 11218 28030 11230 28082
rect 11282 28030 11294 28082
rect 5294 28018 5346 28030
rect 9886 28018 9938 28030
rect 13806 28018 13858 28030
rect 18286 28082 18338 28094
rect 18286 28018 18338 28030
rect 18510 28082 18562 28094
rect 24558 28082 24610 28094
rect 20514 28030 20526 28082
rect 20578 28030 20590 28082
rect 18510 28018 18562 28030
rect 24558 28018 24610 28030
rect 24782 28082 24834 28094
rect 24782 28018 24834 28030
rect 37998 28082 38050 28094
rect 37998 28018 38050 28030
rect 38558 28082 38610 28094
rect 38558 28018 38610 28030
rect 39118 28082 39170 28094
rect 39118 28018 39170 28030
rect 39566 28082 39618 28094
rect 39566 28018 39618 28030
rect 39790 28082 39842 28094
rect 39790 28018 39842 28030
rect 40350 28082 40402 28094
rect 40350 28018 40402 28030
rect 41022 28082 41074 28094
rect 41022 28018 41074 28030
rect 41470 28082 41522 28094
rect 41470 28018 41522 28030
rect 47518 28082 47570 28094
rect 47518 28018 47570 28030
rect 5182 27970 5234 27982
rect 9662 27970 9714 27982
rect 14254 27970 14306 27982
rect 21422 27970 21474 27982
rect 26350 27970 26402 27982
rect 3826 27918 3838 27970
rect 3890 27918 3902 27970
rect 6066 27918 6078 27970
rect 6130 27918 6142 27970
rect 6738 27918 6750 27970
rect 6802 27918 6814 27970
rect 8642 27918 8654 27970
rect 8706 27918 8718 27970
rect 11330 27918 11342 27970
rect 11394 27918 11406 27970
rect 17714 27918 17726 27970
rect 17778 27918 17790 27970
rect 24098 27918 24110 27970
rect 24162 27918 24174 27970
rect 5182 27906 5234 27918
rect 9662 27906 9714 27918
rect 14254 27906 14306 27918
rect 21422 27906 21474 27918
rect 26350 27906 26402 27918
rect 27246 27970 27298 27982
rect 34078 27970 34130 27982
rect 28690 27918 28702 27970
rect 28754 27918 28766 27970
rect 29698 27918 29710 27970
rect 29762 27918 29774 27970
rect 32050 27918 32062 27970
rect 32114 27918 32126 27970
rect 27246 27906 27298 27918
rect 34078 27906 34130 27918
rect 34190 27970 34242 27982
rect 39006 27970 39058 27982
rect 36754 27918 36766 27970
rect 36818 27918 36830 27970
rect 34190 27906 34242 27918
rect 39006 27906 39058 27918
rect 39902 27970 39954 27982
rect 39902 27906 39954 27918
rect 47854 27970 47906 27982
rect 47854 27906 47906 27918
rect 9550 27858 9602 27870
rect 15150 27858 15202 27870
rect 18622 27858 18674 27870
rect 4498 27806 4510 27858
rect 4562 27806 4574 27858
rect 6850 27806 6862 27858
rect 6914 27806 6926 27858
rect 7522 27806 7534 27858
rect 7586 27806 7598 27858
rect 8530 27806 8542 27858
rect 8594 27806 8606 27858
rect 8866 27806 8878 27858
rect 8930 27806 8942 27858
rect 10098 27806 10110 27858
rect 10162 27806 10174 27858
rect 10994 27806 11006 27858
rect 11058 27806 11070 27858
rect 12002 27806 12014 27858
rect 12066 27806 12078 27858
rect 12562 27806 12574 27858
rect 12626 27806 12638 27858
rect 12898 27806 12910 27858
rect 12962 27806 12974 27858
rect 17490 27806 17502 27858
rect 17554 27806 17566 27858
rect 9550 27794 9602 27806
rect 15150 27794 15202 27806
rect 18622 27794 18674 27806
rect 19518 27858 19570 27870
rect 24446 27858 24498 27870
rect 26798 27858 26850 27870
rect 22418 27806 22430 27858
rect 22482 27806 22494 27858
rect 22754 27806 22766 27858
rect 22818 27806 22830 27858
rect 23538 27806 23550 27858
rect 23602 27806 23614 27858
rect 25890 27806 25902 27858
rect 25954 27806 25966 27858
rect 19518 27794 19570 27806
rect 24446 27794 24498 27806
rect 26798 27794 26850 27806
rect 27358 27858 27410 27870
rect 27358 27794 27410 27806
rect 27582 27858 27634 27870
rect 33182 27858 33234 27870
rect 27794 27806 27806 27858
rect 27858 27806 27870 27858
rect 28130 27806 28142 27858
rect 28194 27806 28206 27858
rect 29810 27806 29822 27858
rect 29874 27806 29886 27858
rect 31826 27806 31838 27858
rect 31890 27806 31902 27858
rect 27582 27794 27634 27806
rect 33182 27794 33234 27806
rect 33406 27858 33458 27870
rect 33406 27794 33458 27806
rect 33630 27858 33682 27870
rect 33630 27794 33682 27806
rect 33854 27858 33906 27870
rect 38110 27858 38162 27870
rect 45838 27858 45890 27870
rect 37426 27806 37438 27858
rect 37490 27806 37502 27858
rect 39330 27806 39342 27858
rect 39394 27806 39406 27858
rect 41794 27806 41806 27858
rect 41858 27806 41870 27858
rect 33854 27794 33906 27806
rect 38110 27794 38162 27806
rect 45838 27794 45890 27806
rect 46398 27858 46450 27870
rect 46398 27794 46450 27806
rect 46510 27858 46562 27870
rect 46510 27794 46562 27806
rect 46622 27858 46674 27870
rect 46622 27794 46674 27806
rect 48190 27858 48242 27870
rect 48190 27794 48242 27806
rect 7422 27746 7474 27758
rect 15486 27746 15538 27758
rect 1698 27694 1710 27746
rect 1762 27694 1774 27746
rect 13122 27694 13134 27746
rect 13186 27694 13198 27746
rect 7422 27682 7474 27694
rect 15486 27682 15538 27694
rect 16830 27746 16882 27758
rect 20638 27746 20690 27758
rect 33518 27746 33570 27758
rect 17938 27694 17950 27746
rect 18002 27694 18014 27746
rect 19058 27694 19070 27746
rect 19122 27694 19134 27746
rect 23314 27694 23326 27746
rect 23378 27694 23390 27746
rect 25554 27694 25566 27746
rect 25618 27694 25630 27746
rect 27234 27694 27246 27746
rect 27298 27694 27310 27746
rect 31042 27694 31054 27746
rect 31106 27694 31118 27746
rect 34626 27694 34638 27746
rect 34690 27694 34702 27746
rect 42578 27694 42590 27746
rect 42642 27694 42654 27746
rect 44706 27694 44718 27746
rect 44770 27694 44782 27746
rect 16830 27682 16882 27694
rect 20638 27682 20690 27694
rect 33518 27682 33570 27694
rect 5406 27634 5458 27646
rect 37998 27634 38050 27646
rect 26562 27582 26574 27634
rect 26626 27631 26638 27634
rect 26898 27631 26910 27634
rect 26626 27585 26910 27631
rect 26626 27582 26638 27585
rect 26898 27582 26910 27585
rect 26962 27582 26974 27634
rect 5406 27570 5458 27582
rect 37998 27570 38050 27582
rect 45502 27634 45554 27646
rect 45502 27570 45554 27582
rect 45614 27634 45666 27646
rect 45614 27570 45666 27582
rect 45950 27634 46002 27646
rect 47058 27582 47070 27634
rect 47122 27582 47134 27634
rect 45950 27570 46002 27582
rect 1344 27466 48608 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 48608 27466
rect 1344 27380 48608 27414
rect 29374 27298 29426 27310
rect 20402 27246 20414 27298
rect 20466 27246 20478 27298
rect 30370 27246 30382 27298
rect 30434 27246 30446 27298
rect 29374 27234 29426 27246
rect 18398 27186 18450 27198
rect 23326 27186 23378 27198
rect 2034 27134 2046 27186
rect 2098 27134 2110 27186
rect 6514 27134 6526 27186
rect 6578 27134 6590 27186
rect 8306 27134 8318 27186
rect 8370 27134 8382 27186
rect 13570 27134 13582 27186
rect 13634 27134 13646 27186
rect 19954 27134 19966 27186
rect 20018 27134 20030 27186
rect 18398 27122 18450 27134
rect 23326 27122 23378 27134
rect 25118 27186 25170 27198
rect 25118 27122 25170 27134
rect 26462 27186 26514 27198
rect 28030 27186 28082 27198
rect 27458 27134 27470 27186
rect 27522 27134 27534 27186
rect 26462 27122 26514 27134
rect 28030 27122 28082 27134
rect 29150 27186 29202 27198
rect 30930 27134 30942 27186
rect 30994 27134 31006 27186
rect 32162 27134 32174 27186
rect 32226 27134 32238 27186
rect 34290 27134 34302 27186
rect 34354 27134 34366 27186
rect 40002 27134 40014 27186
rect 40066 27134 40078 27186
rect 40450 27134 40462 27186
rect 40514 27134 40526 27186
rect 42130 27134 42142 27186
rect 42194 27134 42206 27186
rect 44258 27134 44270 27186
rect 44322 27134 44334 27186
rect 46050 27134 46062 27186
rect 46114 27134 46126 27186
rect 48178 27134 48190 27186
rect 48242 27134 48254 27186
rect 29150 27122 29202 27134
rect 5070 27074 5122 27086
rect 12350 27074 12402 27086
rect 3602 27022 3614 27074
rect 3666 27022 3678 27074
rect 5842 27022 5854 27074
rect 5906 27022 5918 27074
rect 6962 27022 6974 27074
rect 7026 27022 7038 27074
rect 7522 27022 7534 27074
rect 7586 27022 7598 27074
rect 10434 27022 10446 27074
rect 10498 27022 10510 27074
rect 10882 27022 10894 27074
rect 10946 27022 10958 27074
rect 11778 27022 11790 27074
rect 11842 27022 11854 27074
rect 5070 27010 5122 27022
rect 12350 27010 12402 27022
rect 12686 27074 12738 27086
rect 12686 27010 12738 27022
rect 13022 27074 13074 27086
rect 19182 27074 19234 27086
rect 22094 27074 22146 27086
rect 23214 27074 23266 27086
rect 26350 27074 26402 27086
rect 13682 27022 13694 27074
rect 13746 27022 13758 27074
rect 15810 27022 15822 27074
rect 15874 27022 15886 27074
rect 16482 27022 16494 27074
rect 16546 27022 16558 27074
rect 17154 27022 17166 27074
rect 17218 27022 17230 27074
rect 18050 27022 18062 27074
rect 18114 27022 18126 27074
rect 18946 27022 18958 27074
rect 19010 27022 19022 27074
rect 19842 27022 19854 27074
rect 19906 27022 19918 27074
rect 20066 27022 20078 27074
rect 20130 27022 20142 27074
rect 22530 27022 22542 27074
rect 22594 27022 22606 27074
rect 25330 27022 25342 27074
rect 25394 27022 25406 27074
rect 13022 27010 13074 27022
rect 19182 27010 19234 27022
rect 22094 27010 22146 27022
rect 23214 27010 23266 27022
rect 26350 27010 26402 27022
rect 26574 27074 26626 27086
rect 26574 27010 26626 27022
rect 28254 27074 28306 27086
rect 30594 27022 30606 27074
rect 30658 27022 30670 27074
rect 35074 27022 35086 27074
rect 35138 27022 35150 27074
rect 37202 27022 37214 27074
rect 37266 27022 37278 27074
rect 40786 27022 40798 27074
rect 40850 27022 40862 27074
rect 41458 27022 41470 27074
rect 41522 27022 41534 27074
rect 45378 27022 45390 27074
rect 45442 27022 45454 27074
rect 28254 27010 28306 27022
rect 12014 26962 12066 26974
rect 3154 26910 3166 26962
rect 3218 26910 3230 26962
rect 4162 26910 4174 26962
rect 4226 26910 4238 26962
rect 4834 26910 4846 26962
rect 4898 26910 4910 26962
rect 5954 26910 5966 26962
rect 6018 26910 6030 26962
rect 7634 26910 7646 26962
rect 7698 26910 7710 26962
rect 12014 26898 12066 26910
rect 12798 26962 12850 26974
rect 26798 26962 26850 26974
rect 15138 26910 15150 26962
rect 15202 26910 15214 26962
rect 15586 26910 15598 26962
rect 15650 26910 15662 26962
rect 17826 26910 17838 26962
rect 17890 26910 17902 26962
rect 12798 26898 12850 26910
rect 26798 26898 26850 26910
rect 27246 26962 27298 26974
rect 44942 26962 44994 26974
rect 37874 26910 37886 26962
rect 37938 26910 37950 26962
rect 27246 26898 27298 26910
rect 44942 26898 44994 26910
rect 2494 26850 2546 26862
rect 21534 26850 21586 26862
rect 4498 26798 4510 26850
rect 4562 26798 4574 26850
rect 16370 26798 16382 26850
rect 16434 26798 16446 26850
rect 17042 26798 17054 26850
rect 17106 26798 17118 26850
rect 2494 26786 2546 26798
rect 21534 26786 21586 26798
rect 27470 26850 27522 26862
rect 31838 26850 31890 26862
rect 28578 26798 28590 26850
rect 28642 26798 28654 26850
rect 29698 26798 29710 26850
rect 29762 26798 29774 26850
rect 27470 26786 27522 26798
rect 31838 26786 31890 26798
rect 1344 26682 48608 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 48608 26682
rect 1344 26596 48608 26630
rect 4734 26514 4786 26526
rect 4734 26450 4786 26462
rect 11118 26514 11170 26526
rect 26686 26514 26738 26526
rect 24322 26462 24334 26514
rect 24386 26462 24398 26514
rect 11118 26450 11170 26462
rect 26686 26450 26738 26462
rect 33406 26514 33458 26526
rect 33406 26450 33458 26462
rect 37662 26514 37714 26526
rect 37662 26450 37714 26462
rect 38670 26514 38722 26526
rect 46722 26462 46734 26514
rect 46786 26462 46798 26514
rect 38670 26450 38722 26462
rect 6302 26402 6354 26414
rect 14254 26402 14306 26414
rect 17278 26402 17330 26414
rect 10210 26350 10222 26402
rect 10274 26350 10286 26402
rect 10546 26350 10558 26402
rect 10610 26350 10622 26402
rect 16370 26350 16382 26402
rect 16434 26350 16446 26402
rect 6302 26338 6354 26350
rect 14254 26338 14306 26350
rect 17278 26338 17330 26350
rect 19518 26402 19570 26414
rect 19518 26338 19570 26350
rect 26238 26402 26290 26414
rect 26238 26338 26290 26350
rect 31390 26402 31442 26414
rect 37550 26402 37602 26414
rect 35746 26350 35758 26402
rect 35810 26350 35822 26402
rect 31390 26338 31442 26350
rect 37550 26338 37602 26350
rect 37774 26402 37826 26414
rect 37774 26338 37826 26350
rect 38222 26402 38274 26414
rect 38222 26338 38274 26350
rect 38894 26402 38946 26414
rect 38894 26338 38946 26350
rect 39566 26402 39618 26414
rect 39566 26338 39618 26350
rect 42366 26402 42418 26414
rect 42366 26338 42418 26350
rect 42814 26402 42866 26414
rect 42814 26338 42866 26350
rect 45614 26402 45666 26414
rect 45614 26338 45666 26350
rect 47070 26402 47122 26414
rect 47070 26338 47122 26350
rect 4622 26290 4674 26302
rect 6414 26290 6466 26302
rect 2258 26238 2270 26290
rect 2322 26238 2334 26290
rect 3042 26238 3054 26290
rect 3106 26238 3118 26290
rect 4162 26238 4174 26290
rect 4226 26238 4238 26290
rect 6066 26238 6078 26290
rect 6130 26238 6142 26290
rect 4622 26226 4674 26238
rect 6414 26226 6466 26238
rect 8206 26290 8258 26302
rect 12126 26290 12178 26302
rect 19070 26290 19122 26302
rect 8978 26238 8990 26290
rect 9042 26238 9054 26290
rect 11554 26238 11566 26290
rect 11618 26238 11630 26290
rect 15138 26238 15150 26290
rect 15202 26238 15214 26290
rect 15698 26238 15710 26290
rect 15762 26238 15774 26290
rect 16034 26238 16046 26290
rect 16098 26238 16110 26290
rect 17602 26238 17614 26290
rect 17666 26238 17678 26290
rect 8206 26226 8258 26238
rect 12126 26226 12178 26238
rect 19070 26226 19122 26238
rect 19406 26290 19458 26302
rect 19406 26226 19458 26238
rect 19742 26290 19794 26302
rect 19742 26226 19794 26238
rect 20302 26290 20354 26302
rect 20302 26226 20354 26238
rect 20526 26290 20578 26302
rect 20526 26226 20578 26238
rect 20638 26290 20690 26302
rect 22318 26290 22370 26302
rect 23998 26290 24050 26302
rect 21522 26238 21534 26290
rect 21586 26238 21598 26290
rect 22754 26238 22766 26290
rect 22818 26238 22830 26290
rect 23202 26238 23214 26290
rect 23266 26238 23278 26290
rect 20638 26226 20690 26238
rect 22318 26226 22370 26238
rect 23998 26226 24050 26238
rect 26574 26290 26626 26302
rect 26574 26226 26626 26238
rect 26798 26290 26850 26302
rect 26798 26226 26850 26238
rect 27246 26290 27298 26302
rect 30270 26290 30322 26302
rect 27458 26238 27470 26290
rect 27522 26238 27534 26290
rect 28578 26238 28590 26290
rect 28642 26238 28654 26290
rect 27246 26226 27298 26238
rect 30270 26226 30322 26238
rect 30606 26290 30658 26302
rect 32958 26290 33010 26302
rect 31826 26238 31838 26290
rect 31890 26238 31902 26290
rect 30606 26226 30658 26238
rect 32958 26226 33010 26238
rect 33518 26290 33570 26302
rect 33518 26226 33570 26238
rect 33630 26290 33682 26302
rect 35422 26290 35474 26302
rect 38446 26290 38498 26302
rect 34962 26238 34974 26290
rect 35026 26238 35038 26290
rect 35858 26238 35870 26290
rect 35922 26238 35934 26290
rect 36418 26238 36430 26290
rect 36482 26238 36494 26290
rect 37202 26238 37214 26290
rect 37266 26238 37278 26290
rect 33630 26226 33682 26238
rect 35422 26226 35474 26238
rect 38446 26226 38498 26238
rect 39006 26290 39058 26302
rect 43250 26238 43262 26290
rect 43314 26238 43326 26290
rect 46162 26238 46174 26290
rect 46226 26238 46238 26290
rect 48178 26238 48190 26290
rect 48242 26238 48254 26290
rect 39006 26226 39058 26238
rect 12462 26178 12514 26190
rect 23774 26178 23826 26190
rect 2930 26126 2942 26178
rect 2994 26126 3006 26178
rect 16482 26126 16494 26178
rect 16546 26126 16558 26178
rect 21410 26126 21422 26178
rect 21474 26126 21486 26178
rect 12462 26114 12514 26126
rect 23774 26114 23826 26126
rect 25454 26178 25506 26190
rect 34078 26178 34130 26190
rect 39454 26178 39506 26190
rect 25778 26126 25790 26178
rect 25842 26126 25854 26178
rect 27570 26126 27582 26178
rect 27634 26126 27646 26178
rect 32162 26126 32174 26178
rect 32226 26126 32238 26178
rect 34514 26126 34526 26178
rect 34578 26126 34590 26178
rect 38098 26126 38110 26178
rect 38162 26126 38174 26178
rect 25454 26114 25506 26126
rect 34078 26114 34130 26126
rect 39454 26114 39506 26126
rect 40014 26178 40066 26190
rect 40014 26114 40066 26126
rect 41918 26178 41970 26190
rect 41918 26114 41970 26126
rect 42142 26178 42194 26190
rect 42466 26126 42478 26178
rect 42530 26126 42542 26178
rect 43698 26126 43710 26178
rect 43762 26126 43774 26178
rect 42142 26114 42194 26126
rect 4734 26066 4786 26078
rect 4734 26002 4786 26014
rect 10782 26066 10834 26078
rect 10782 26002 10834 26014
rect 20078 26066 20130 26078
rect 20078 26002 20130 26014
rect 20862 26066 20914 26078
rect 22866 26014 22878 26066
rect 22930 26014 22942 26066
rect 20862 26002 20914 26014
rect 1344 25898 48608 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 48608 25898
rect 1344 25812 48608 25846
rect 12798 25730 12850 25742
rect 6962 25678 6974 25730
rect 7026 25678 7038 25730
rect 12798 25666 12850 25678
rect 13918 25730 13970 25742
rect 13918 25666 13970 25678
rect 17726 25730 17778 25742
rect 26238 25730 26290 25742
rect 47630 25730 47682 25742
rect 23202 25678 23214 25730
rect 23266 25678 23278 25730
rect 29474 25678 29486 25730
rect 29538 25678 29550 25730
rect 17726 25666 17778 25678
rect 26238 25666 26290 25678
rect 47630 25666 47682 25678
rect 14254 25618 14306 25630
rect 24558 25618 24610 25630
rect 35982 25618 36034 25630
rect 2482 25566 2494 25618
rect 2546 25566 2558 25618
rect 4610 25566 4622 25618
rect 4674 25566 4686 25618
rect 8642 25566 8654 25618
rect 8706 25566 8718 25618
rect 21858 25566 21870 25618
rect 21922 25566 21934 25618
rect 27570 25566 27582 25618
rect 27634 25566 27646 25618
rect 29586 25566 29598 25618
rect 29650 25566 29662 25618
rect 31154 25566 31166 25618
rect 31218 25566 31230 25618
rect 14254 25554 14306 25566
rect 24558 25554 24610 25566
rect 35982 25554 36034 25566
rect 39230 25618 39282 25630
rect 39230 25554 39282 25566
rect 43486 25618 43538 25630
rect 43486 25554 43538 25566
rect 43934 25618 43986 25630
rect 43934 25554 43986 25566
rect 44382 25618 44434 25630
rect 44382 25554 44434 25566
rect 46398 25618 46450 25630
rect 46398 25554 46450 25566
rect 47294 25618 47346 25630
rect 47294 25554 47346 25566
rect 48190 25618 48242 25630
rect 48190 25554 48242 25566
rect 6302 25506 6354 25518
rect 14702 25506 14754 25518
rect 19966 25506 20018 25518
rect 24670 25506 24722 25518
rect 26014 25506 26066 25518
rect 1810 25454 1822 25506
rect 1874 25454 1886 25506
rect 5730 25454 5742 25506
rect 5794 25454 5806 25506
rect 6626 25454 6638 25506
rect 6690 25454 6702 25506
rect 7746 25454 7758 25506
rect 7810 25454 7822 25506
rect 8530 25454 8542 25506
rect 8594 25454 8606 25506
rect 11106 25454 11118 25506
rect 11170 25454 11182 25506
rect 12898 25454 12910 25506
rect 12962 25454 12974 25506
rect 17490 25454 17502 25506
rect 17554 25454 17566 25506
rect 18162 25454 18174 25506
rect 18226 25454 18238 25506
rect 21746 25454 21758 25506
rect 21810 25454 21822 25506
rect 23426 25454 23438 25506
rect 23490 25454 23502 25506
rect 24994 25454 25006 25506
rect 25058 25454 25070 25506
rect 6302 25442 6354 25454
rect 14702 25442 14754 25454
rect 19966 25442 20018 25454
rect 24670 25442 24722 25454
rect 26014 25442 26066 25454
rect 26686 25506 26738 25518
rect 30718 25506 30770 25518
rect 34974 25506 35026 25518
rect 29474 25454 29486 25506
rect 29538 25454 29550 25506
rect 30482 25454 30494 25506
rect 30546 25454 30558 25506
rect 32274 25454 32286 25506
rect 32338 25454 32350 25506
rect 34514 25454 34526 25506
rect 34578 25454 34590 25506
rect 26686 25442 26738 25454
rect 30718 25442 30770 25454
rect 34974 25442 35026 25454
rect 36990 25506 37042 25518
rect 45054 25506 45106 25518
rect 40226 25454 40238 25506
rect 40290 25454 40302 25506
rect 40898 25454 40910 25506
rect 40962 25454 40974 25506
rect 36990 25442 37042 25454
rect 45054 25442 45106 25454
rect 45166 25506 45218 25518
rect 46510 25506 46562 25518
rect 45602 25454 45614 25506
rect 45666 25454 45678 25506
rect 45166 25442 45218 25454
rect 46510 25442 46562 25454
rect 46846 25506 46898 25518
rect 46846 25442 46898 25454
rect 47406 25506 47458 25518
rect 47406 25442 47458 25454
rect 5966 25394 6018 25406
rect 13694 25394 13746 25406
rect 19182 25394 19234 25406
rect 9426 25342 9438 25394
rect 9490 25342 9502 25394
rect 12226 25342 12238 25394
rect 12290 25342 12302 25394
rect 16258 25342 16270 25394
rect 16322 25342 16334 25394
rect 16930 25342 16942 25394
rect 16994 25342 17006 25394
rect 5966 25330 6018 25342
rect 13694 25330 13746 25342
rect 19182 25330 19234 25342
rect 27918 25394 27970 25406
rect 27918 25330 27970 25342
rect 28590 25394 28642 25406
rect 28590 25330 28642 25342
rect 31278 25394 31330 25406
rect 35422 25394 35474 25406
rect 32162 25342 32174 25394
rect 32226 25342 32238 25394
rect 33618 25342 33630 25394
rect 33682 25342 33694 25394
rect 31278 25330 31330 25342
rect 35422 25330 35474 25342
rect 35534 25394 35586 25406
rect 35534 25330 35586 25342
rect 41918 25394 41970 25406
rect 41918 25330 41970 25342
rect 44942 25394 44994 25406
rect 46286 25394 46338 25406
rect 45826 25342 45838 25394
rect 45890 25342 45902 25394
rect 44942 25330 44994 25342
rect 46286 25330 46338 25342
rect 5070 25282 5122 25294
rect 5070 25218 5122 25230
rect 18286 25282 18338 25294
rect 31054 25282 31106 25294
rect 35198 25282 35250 25294
rect 28242 25230 28254 25282
rect 28306 25230 28318 25282
rect 33506 25230 33518 25282
rect 33570 25230 33582 25282
rect 18286 25218 18338 25230
rect 31054 25218 31106 25230
rect 35198 25218 35250 25230
rect 36542 25282 36594 25294
rect 36542 25218 36594 25230
rect 37102 25282 37154 25294
rect 37102 25218 37154 25230
rect 37214 25282 37266 25294
rect 37214 25218 37266 25230
rect 37438 25282 37490 25294
rect 37438 25218 37490 25230
rect 39790 25282 39842 25294
rect 41582 25282 41634 25294
rect 40450 25230 40462 25282
rect 40514 25230 40526 25282
rect 41122 25230 41134 25282
rect 41186 25230 41198 25282
rect 39790 25218 39842 25230
rect 41582 25218 41634 25230
rect 47294 25282 47346 25294
rect 47294 25218 47346 25230
rect 1344 25114 48608 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 48608 25114
rect 1344 25028 48608 25062
rect 2158 24946 2210 24958
rect 2158 24882 2210 24894
rect 2606 24946 2658 24958
rect 2606 24882 2658 24894
rect 5630 24946 5682 24958
rect 5630 24882 5682 24894
rect 6526 24946 6578 24958
rect 6526 24882 6578 24894
rect 9774 24946 9826 24958
rect 9774 24882 9826 24894
rect 13022 24946 13074 24958
rect 13022 24882 13074 24894
rect 16830 24946 16882 24958
rect 19518 24946 19570 24958
rect 34862 24946 34914 24958
rect 17490 24894 17502 24946
rect 17554 24894 17566 24946
rect 31826 24894 31838 24946
rect 31890 24894 31902 24946
rect 46946 24894 46958 24946
rect 47010 24894 47022 24946
rect 16830 24882 16882 24894
rect 19518 24882 19570 24894
rect 34862 24882 34914 24894
rect 2942 24834 2994 24846
rect 2942 24770 2994 24782
rect 3838 24834 3890 24846
rect 3838 24770 3890 24782
rect 6974 24834 7026 24846
rect 6974 24770 7026 24782
rect 12574 24834 12626 24846
rect 12574 24770 12626 24782
rect 16494 24834 16546 24846
rect 18958 24834 19010 24846
rect 17602 24782 17614 24834
rect 17666 24782 17678 24834
rect 18274 24782 18286 24834
rect 18338 24782 18350 24834
rect 16494 24770 16546 24782
rect 18958 24770 19010 24782
rect 19966 24834 20018 24846
rect 23650 24782 23662 24834
rect 23714 24782 23726 24834
rect 28802 24782 28814 24834
rect 28866 24782 28878 24834
rect 31154 24782 31166 24834
rect 31218 24782 31230 24834
rect 31490 24782 31502 24834
rect 31554 24782 31566 24834
rect 33730 24782 33742 24834
rect 33794 24782 33806 24834
rect 40338 24782 40350 24834
rect 40402 24782 40414 24834
rect 19966 24770 20018 24782
rect 2270 24722 2322 24734
rect 2270 24658 2322 24670
rect 2718 24722 2770 24734
rect 2718 24658 2770 24670
rect 3390 24722 3442 24734
rect 3390 24658 3442 24670
rect 5070 24722 5122 24734
rect 5070 24658 5122 24670
rect 6526 24722 6578 24734
rect 6526 24658 6578 24670
rect 8206 24722 8258 24734
rect 8206 24658 8258 24670
rect 9438 24722 9490 24734
rect 9438 24658 9490 24670
rect 9886 24722 9938 24734
rect 9886 24658 9938 24670
rect 10110 24722 10162 24734
rect 17502 24722 17554 24734
rect 13122 24670 13134 24722
rect 13186 24670 13198 24722
rect 14018 24670 14030 24722
rect 14082 24670 14094 24722
rect 15922 24670 15934 24722
rect 15986 24670 15998 24722
rect 10110 24658 10162 24670
rect 17502 24658 17554 24670
rect 19070 24722 19122 24734
rect 19070 24658 19122 24670
rect 20862 24722 20914 24734
rect 20862 24658 20914 24670
rect 22654 24722 22706 24734
rect 35086 24722 35138 24734
rect 39118 24722 39170 24734
rect 23090 24670 23102 24722
rect 23154 24670 23166 24722
rect 23538 24670 23550 24722
rect 23602 24670 23614 24722
rect 24434 24670 24446 24722
rect 24498 24670 24510 24722
rect 25218 24670 25230 24722
rect 25282 24670 25294 24722
rect 30930 24670 30942 24722
rect 30994 24670 31006 24722
rect 33618 24670 33630 24722
rect 33682 24670 33694 24722
rect 34290 24670 34302 24722
rect 34354 24670 34366 24722
rect 38770 24670 38782 24722
rect 38834 24670 38846 24722
rect 22654 24658 22706 24670
rect 35086 24658 35138 24670
rect 39118 24658 39170 24670
rect 39678 24722 39730 24734
rect 39678 24658 39730 24670
rect 40014 24722 40066 24734
rect 40014 24658 40066 24670
rect 40910 24722 40962 24734
rect 40910 24658 40962 24670
rect 41470 24722 41522 24734
rect 47294 24722 47346 24734
rect 42242 24670 42254 24722
rect 42306 24670 42318 24722
rect 45938 24670 45950 24722
rect 46002 24670 46014 24722
rect 41470 24658 41522 24670
rect 47294 24658 47346 24670
rect 47518 24722 47570 24734
rect 47518 24658 47570 24670
rect 47966 24722 48018 24734
rect 47966 24658 48018 24670
rect 11342 24610 11394 24622
rect 21198 24610 21250 24622
rect 32510 24610 32562 24622
rect 14130 24558 14142 24610
rect 14194 24558 14206 24610
rect 15586 24558 15598 24610
rect 15650 24558 15662 24610
rect 23874 24558 23886 24610
rect 23938 24558 23950 24610
rect 33842 24558 33854 24610
rect 33906 24558 33918 24610
rect 34738 24558 34750 24610
rect 34802 24558 34814 24610
rect 35858 24558 35870 24610
rect 35922 24558 35934 24610
rect 37986 24558 37998 24610
rect 38050 24558 38062 24610
rect 43026 24558 43038 24610
rect 43090 24558 43102 24610
rect 45154 24558 45166 24610
rect 45218 24558 45230 24610
rect 46386 24558 46398 24610
rect 46450 24558 46462 24610
rect 11342 24546 11394 24558
rect 21198 24546 21250 24558
rect 32510 24546 32562 24558
rect 18958 24498 19010 24510
rect 47854 24498 47906 24510
rect 45602 24446 45614 24498
rect 45666 24446 45678 24498
rect 18958 24434 19010 24446
rect 47854 24434 47906 24446
rect 1344 24330 48608 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 48608 24330
rect 1344 24244 48608 24278
rect 6190 24162 6242 24174
rect 29934 24162 29986 24174
rect 2370 24110 2382 24162
rect 2434 24110 2446 24162
rect 8978 24110 8990 24162
rect 9042 24110 9054 24162
rect 11554 24110 11566 24162
rect 11618 24110 11630 24162
rect 19618 24110 19630 24162
rect 19682 24110 19694 24162
rect 6190 24098 6242 24110
rect 29934 24098 29986 24110
rect 37214 24162 37266 24174
rect 37214 24098 37266 24110
rect 37886 24162 37938 24174
rect 37886 24098 37938 24110
rect 43150 24162 43202 24174
rect 43150 24098 43202 24110
rect 43486 24162 43538 24174
rect 43486 24098 43538 24110
rect 14142 24050 14194 24062
rect 24446 24050 24498 24062
rect 4946 23998 4958 24050
rect 5010 23998 5022 24050
rect 8082 23998 8094 24050
rect 8146 23998 8158 24050
rect 12002 23998 12014 24050
rect 12066 23998 12078 24050
rect 18834 23998 18846 24050
rect 18898 23998 18910 24050
rect 20178 23998 20190 24050
rect 20242 23998 20254 24050
rect 14142 23986 14194 23998
rect 24446 23986 24498 23998
rect 24558 24050 24610 24062
rect 24558 23986 24610 23998
rect 29150 24050 29202 24062
rect 29150 23986 29202 23998
rect 30942 24050 30994 24062
rect 30942 23986 30994 23998
rect 31390 24050 31442 24062
rect 31390 23986 31442 23998
rect 32286 24050 32338 24062
rect 32286 23986 32338 23998
rect 32734 24050 32786 24062
rect 36990 24050 37042 24062
rect 33058 23998 33070 24050
rect 33122 23998 33134 24050
rect 32734 23986 32786 23998
rect 36990 23986 37042 23998
rect 37998 24050 38050 24062
rect 42142 24050 42194 24062
rect 40562 23998 40574 24050
rect 40626 23998 40638 24050
rect 37998 23986 38050 23998
rect 42142 23986 42194 23998
rect 45054 24050 45106 24062
rect 46050 23998 46062 24050
rect 46114 23998 46126 24050
rect 48178 23998 48190 24050
rect 48242 23998 48254 24050
rect 45054 23986 45106 23998
rect 4510 23938 4562 23950
rect 10558 23938 10610 23950
rect 19742 23938 19794 23950
rect 23102 23938 23154 23950
rect 26798 23938 26850 23950
rect 4274 23886 4286 23938
rect 4338 23886 4350 23938
rect 7746 23886 7758 23938
rect 7810 23886 7822 23938
rect 9650 23886 9662 23938
rect 9714 23886 9726 23938
rect 11666 23886 11678 23938
rect 11730 23886 11742 23938
rect 12450 23886 12462 23938
rect 12514 23886 12526 23938
rect 13458 23886 13470 23938
rect 13522 23886 13534 23938
rect 14690 23886 14702 23938
rect 14754 23886 14766 23938
rect 15026 23886 15038 23938
rect 15090 23886 15102 23938
rect 16034 23886 16046 23938
rect 16098 23886 16110 23938
rect 20066 23886 20078 23938
rect 20130 23886 20142 23938
rect 21410 23886 21422 23938
rect 21474 23886 21486 23938
rect 21858 23886 21870 23938
rect 21922 23886 21934 23938
rect 22642 23886 22654 23938
rect 22706 23886 22718 23938
rect 23762 23886 23774 23938
rect 23826 23886 23838 23938
rect 24994 23886 25006 23938
rect 25058 23886 25070 23938
rect 4510 23874 4562 23886
rect 10558 23874 10610 23886
rect 19742 23874 19794 23886
rect 23102 23874 23154 23886
rect 26798 23874 26850 23886
rect 27134 23938 27186 23950
rect 30606 23938 30658 23950
rect 30258 23886 30270 23938
rect 30322 23886 30334 23938
rect 27134 23874 27186 23886
rect 30606 23874 30658 23886
rect 31726 23938 31778 23950
rect 41582 23938 41634 23950
rect 35858 23886 35870 23938
rect 35922 23886 35934 23938
rect 38210 23886 38222 23938
rect 38274 23886 38286 23938
rect 42690 23886 42702 23938
rect 42754 23886 42766 23938
rect 43138 23886 43150 23938
rect 43202 23886 43214 23938
rect 45378 23886 45390 23938
rect 45442 23886 45454 23938
rect 31726 23874 31778 23886
rect 41582 23874 41634 23886
rect 15374 23826 15426 23838
rect 5618 23774 5630 23826
rect 5682 23774 5694 23826
rect 10882 23774 10894 23826
rect 10946 23774 10958 23826
rect 13570 23774 13582 23826
rect 13634 23774 13646 23826
rect 15374 23762 15426 23774
rect 15486 23826 15538 23838
rect 23438 23826 23490 23838
rect 27582 23826 27634 23838
rect 16706 23774 16718 23826
rect 16770 23774 16782 23826
rect 21298 23774 21310 23826
rect 21362 23774 21374 23826
rect 24210 23774 24222 23826
rect 24274 23774 24286 23826
rect 30818 23774 30830 23826
rect 30882 23774 30894 23826
rect 35186 23774 35198 23826
rect 35250 23774 35262 23826
rect 37538 23774 37550 23826
rect 37602 23774 37614 23826
rect 15486 23762 15538 23774
rect 23438 23762 23490 23774
rect 27582 23762 27634 23774
rect 4846 23714 4898 23726
rect 4846 23650 4898 23662
rect 5070 23714 5122 23726
rect 5070 23650 5122 23662
rect 15710 23714 15762 23726
rect 15710 23650 15762 23662
rect 23326 23714 23378 23726
rect 23326 23650 23378 23662
rect 27022 23714 27074 23726
rect 27022 23650 27074 23662
rect 29710 23714 29762 23726
rect 29710 23650 29762 23662
rect 40126 23714 40178 23726
rect 40126 23650 40178 23662
rect 41134 23714 41186 23726
rect 41134 23650 41186 23662
rect 42478 23714 42530 23726
rect 42478 23650 42530 23662
rect 1344 23546 48608 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 48608 23546
rect 1344 23460 48608 23494
rect 12350 23378 12402 23390
rect 8306 23326 8318 23378
rect 8370 23326 8382 23378
rect 12350 23314 12402 23326
rect 22766 23378 22818 23390
rect 35758 23378 35810 23390
rect 23202 23326 23214 23378
rect 23266 23326 23278 23378
rect 22766 23314 22818 23326
rect 35758 23314 35810 23326
rect 44382 23378 44434 23390
rect 44382 23314 44434 23326
rect 46062 23378 46114 23390
rect 46062 23314 46114 23326
rect 7422 23266 7474 23278
rect 12798 23266 12850 23278
rect 9538 23214 9550 23266
rect 9602 23214 9614 23266
rect 7422 23202 7474 23214
rect 12798 23202 12850 23214
rect 18398 23266 18450 23278
rect 18398 23202 18450 23214
rect 22430 23266 22482 23278
rect 22430 23202 22482 23214
rect 22878 23266 22930 23278
rect 22878 23202 22930 23214
rect 24670 23266 24722 23278
rect 24670 23202 24722 23214
rect 26014 23266 26066 23278
rect 38110 23266 38162 23278
rect 26562 23214 26574 23266
rect 26626 23214 26638 23266
rect 28466 23214 28478 23266
rect 28530 23214 28542 23266
rect 30034 23214 30046 23266
rect 30098 23214 30110 23266
rect 31266 23214 31278 23266
rect 31330 23214 31342 23266
rect 31714 23214 31726 23266
rect 31778 23214 31790 23266
rect 26014 23202 26066 23214
rect 38110 23202 38162 23214
rect 44942 23266 44994 23278
rect 44942 23202 44994 23214
rect 45838 23266 45890 23278
rect 47966 23266 48018 23278
rect 47170 23214 47182 23266
rect 47234 23214 47246 23266
rect 45838 23202 45890 23214
rect 47966 23202 48018 23214
rect 6190 23154 6242 23166
rect 22654 23154 22706 23166
rect 24334 23154 24386 23166
rect 30942 23154 30994 23166
rect 1810 23102 1822 23154
rect 1874 23102 1886 23154
rect 7970 23102 7982 23154
rect 8034 23102 8046 23154
rect 12226 23102 12238 23154
rect 12290 23102 12302 23154
rect 14130 23102 14142 23154
rect 14194 23102 14206 23154
rect 16594 23102 16606 23154
rect 16658 23102 16670 23154
rect 17826 23102 17838 23154
rect 17890 23102 17902 23154
rect 18834 23102 18846 23154
rect 18898 23102 18910 23154
rect 24098 23102 24110 23154
rect 24162 23102 24174 23154
rect 25554 23102 25566 23154
rect 25618 23102 25630 23154
rect 25890 23102 25902 23154
rect 25954 23102 25966 23154
rect 27122 23102 27134 23154
rect 27186 23102 27198 23154
rect 28242 23102 28254 23154
rect 28306 23102 28318 23154
rect 30258 23102 30270 23154
rect 30322 23102 30334 23154
rect 6190 23090 6242 23102
rect 22654 23090 22706 23102
rect 24334 23090 24386 23102
rect 30942 23090 30994 23102
rect 32510 23154 32562 23166
rect 32510 23090 32562 23102
rect 32958 23154 33010 23166
rect 32958 23090 33010 23102
rect 33406 23154 33458 23166
rect 33406 23090 33458 23102
rect 33630 23154 33682 23166
rect 45166 23154 45218 23166
rect 34402 23102 34414 23154
rect 34466 23102 34478 23154
rect 38322 23102 38334 23154
rect 38386 23102 38398 23154
rect 38546 23102 38558 23154
rect 38610 23102 38622 23154
rect 38882 23102 38894 23154
rect 38946 23102 38958 23154
rect 41010 23102 41022 23154
rect 41074 23102 41086 23154
rect 33630 23090 33682 23102
rect 45166 23090 45218 23102
rect 45502 23154 45554 23166
rect 45502 23090 45554 23102
rect 46398 23154 46450 23166
rect 46722 23102 46734 23154
rect 46786 23102 46798 23154
rect 47618 23102 47630 23154
rect 47682 23102 47694 23154
rect 46398 23090 46450 23102
rect 8206 23042 8258 23054
rect 2482 22990 2494 23042
rect 2546 22990 2558 23042
rect 4722 22990 4734 23042
rect 4786 22990 4798 23042
rect 8206 22978 8258 22990
rect 12014 23042 12066 23054
rect 23774 23042 23826 23054
rect 14466 22990 14478 23042
rect 14530 22990 14542 23042
rect 16370 22990 16382 23042
rect 16434 22990 16446 23042
rect 17938 22990 17950 23042
rect 18002 22990 18014 23042
rect 19506 22990 19518 23042
rect 19570 22990 19582 23042
rect 21634 22990 21646 23042
rect 21698 22990 21710 23042
rect 12014 22978 12066 22990
rect 23774 22978 23826 22990
rect 30830 23042 30882 23054
rect 30830 22978 30882 22990
rect 33518 23042 33570 23054
rect 33518 22978 33570 22990
rect 33966 23042 34018 23054
rect 36206 23042 36258 23054
rect 35298 22990 35310 23042
rect 35362 22990 35374 23042
rect 35970 22990 35982 23042
rect 36034 22990 36046 23042
rect 33966 22978 34018 22990
rect 10110 22930 10162 22942
rect 10110 22866 10162 22878
rect 23550 22930 23602 22942
rect 23550 22866 23602 22878
rect 24558 22930 24610 22942
rect 35985 22927 36031 22990
rect 36206 22978 36258 22990
rect 36654 23042 36706 23054
rect 36654 22978 36706 22990
rect 37102 23042 37154 23054
rect 37102 22978 37154 22990
rect 38446 23042 38498 23054
rect 38446 22978 38498 22990
rect 39118 23042 39170 23054
rect 44270 23042 44322 23054
rect 41682 22990 41694 23042
rect 41746 22990 41758 23042
rect 43810 22990 43822 23042
rect 43874 22990 43886 23042
rect 39118 22978 39170 22990
rect 44270 22978 44322 22990
rect 45054 23042 45106 23054
rect 47394 22990 47406 23042
rect 47458 22990 47470 23042
rect 45054 22978 45106 22990
rect 39230 22930 39282 22942
rect 36642 22927 36654 22930
rect 35985 22881 36654 22927
rect 36642 22878 36654 22881
rect 36706 22878 36718 22930
rect 24558 22866 24610 22878
rect 39230 22866 39282 22878
rect 44158 22930 44210 22942
rect 44158 22866 44210 22878
rect 45726 22930 45778 22942
rect 45726 22866 45778 22878
rect 1344 22762 48608 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 48608 22762
rect 1344 22676 48608 22710
rect 15150 22594 15202 22606
rect 34974 22594 35026 22606
rect 3378 22542 3390 22594
rect 3442 22542 3454 22594
rect 11106 22542 11118 22594
rect 11170 22542 11182 22594
rect 29586 22542 29598 22594
rect 29650 22542 29662 22594
rect 15150 22530 15202 22542
rect 34974 22530 35026 22542
rect 40574 22594 40626 22606
rect 40574 22530 40626 22542
rect 45950 22594 46002 22606
rect 45950 22530 46002 22542
rect 46622 22594 46674 22606
rect 46622 22530 46674 22542
rect 1822 22482 1874 22494
rect 12910 22482 12962 22494
rect 2818 22430 2830 22482
rect 2882 22430 2894 22482
rect 3938 22430 3950 22482
rect 4002 22430 4014 22482
rect 6066 22430 6078 22482
rect 6130 22430 6142 22482
rect 7746 22430 7758 22482
rect 7810 22430 7822 22482
rect 9986 22430 9998 22482
rect 10050 22430 10062 22482
rect 1822 22418 1874 22430
rect 12910 22418 12962 22430
rect 15262 22482 15314 22494
rect 19966 22482 20018 22494
rect 18722 22430 18734 22482
rect 18786 22430 18798 22482
rect 15262 22418 15314 22430
rect 19966 22418 20018 22430
rect 24446 22482 24498 22494
rect 24446 22418 24498 22430
rect 31390 22482 31442 22494
rect 35086 22482 35138 22494
rect 41134 22482 41186 22494
rect 31714 22430 31726 22482
rect 31778 22430 31790 22482
rect 37202 22430 37214 22482
rect 37266 22430 37278 22482
rect 39330 22430 39342 22482
rect 39394 22430 39406 22482
rect 31390 22418 31442 22430
rect 35086 22418 35138 22430
rect 41134 22418 41186 22430
rect 42254 22482 42306 22494
rect 42254 22418 42306 22430
rect 43598 22482 43650 22494
rect 46946 22430 46958 22482
rect 47010 22430 47022 22482
rect 43598 22418 43650 22430
rect 2382 22370 2434 22382
rect 4846 22370 4898 22382
rect 2930 22318 2942 22370
rect 2994 22318 3006 22370
rect 4498 22318 4510 22370
rect 4562 22318 4574 22370
rect 2382 22306 2434 22318
rect 4846 22306 4898 22318
rect 5630 22370 5682 22382
rect 19742 22370 19794 22382
rect 10658 22318 10670 22370
rect 10722 22318 10734 22370
rect 11666 22318 11678 22370
rect 11730 22318 11742 22370
rect 13458 22318 13470 22370
rect 13522 22318 13534 22370
rect 15922 22318 15934 22370
rect 15986 22318 15998 22370
rect 5630 22306 5682 22318
rect 19742 22306 19794 22318
rect 20078 22370 20130 22382
rect 20078 22306 20130 22318
rect 20414 22370 20466 22382
rect 26350 22370 26402 22382
rect 30830 22370 30882 22382
rect 35758 22370 35810 22382
rect 43934 22370 43986 22382
rect 21522 22318 21534 22370
rect 21586 22318 21598 22370
rect 28130 22318 28142 22370
rect 28194 22318 28206 22370
rect 29250 22318 29262 22370
rect 29314 22318 29326 22370
rect 29698 22318 29710 22370
rect 29762 22318 29774 22370
rect 30594 22318 30606 22370
rect 30658 22318 30670 22370
rect 34514 22318 34526 22370
rect 34578 22318 34590 22370
rect 35298 22318 35310 22370
rect 35362 22318 35374 22370
rect 40114 22318 40126 22370
rect 40178 22318 40190 22370
rect 43138 22318 43150 22370
rect 43202 22318 43214 22370
rect 43362 22318 43374 22370
rect 43426 22318 43438 22370
rect 20414 22306 20466 22318
rect 26350 22306 26402 22318
rect 30830 22306 30882 22318
rect 35758 22306 35810 22318
rect 43934 22306 43986 22318
rect 45502 22370 45554 22382
rect 45502 22306 45554 22318
rect 45726 22370 45778 22382
rect 45726 22306 45778 22318
rect 47182 22370 47234 22382
rect 47182 22306 47234 22318
rect 47518 22370 47570 22382
rect 47518 22306 47570 22318
rect 47742 22370 47794 22382
rect 47742 22306 47794 22318
rect 25230 22258 25282 22270
rect 14242 22206 14254 22258
rect 14306 22206 14318 22258
rect 16594 22206 16606 22258
rect 16658 22206 16670 22258
rect 19058 22206 19070 22258
rect 19122 22206 19134 22258
rect 22306 22206 22318 22258
rect 22370 22206 22382 22258
rect 25230 22194 25282 22206
rect 27582 22258 27634 22270
rect 40462 22258 40514 22270
rect 33842 22206 33854 22258
rect 33906 22206 33918 22258
rect 27582 22194 27634 22206
rect 40462 22194 40514 22206
rect 40574 22258 40626 22270
rect 40574 22194 40626 22206
rect 44270 22258 44322 22270
rect 44270 22194 44322 22206
rect 44830 22258 44882 22270
rect 44830 22194 44882 22206
rect 45054 22258 45106 22270
rect 45054 22194 45106 22206
rect 46846 22258 46898 22270
rect 46846 22194 46898 22206
rect 12350 22146 12402 22158
rect 3826 22094 3838 22146
rect 3890 22094 3902 22146
rect 12350 22082 12402 22094
rect 15374 22146 15426 22158
rect 15374 22082 15426 22094
rect 19406 22146 19458 22158
rect 19406 22082 19458 22094
rect 24894 22146 24946 22158
rect 24894 22082 24946 22094
rect 25118 22146 25170 22158
rect 25118 22082 25170 22094
rect 26686 22146 26738 22158
rect 26686 22082 26738 22094
rect 28702 22146 28754 22158
rect 28702 22082 28754 22094
rect 36206 22146 36258 22158
rect 36206 22082 36258 22094
rect 36318 22146 36370 22158
rect 36318 22082 36370 22094
rect 36430 22146 36482 22158
rect 36430 22082 36482 22094
rect 44046 22146 44098 22158
rect 44046 22082 44098 22094
rect 44942 22146 44994 22158
rect 44942 22082 44994 22094
rect 46398 22146 46450 22158
rect 46398 22082 46450 22094
rect 47518 22146 47570 22158
rect 47518 22082 47570 22094
rect 1344 21978 48608 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 48608 21978
rect 1344 21892 48608 21926
rect 9774 21810 9826 21822
rect 8306 21758 8318 21810
rect 8370 21758 8382 21810
rect 9774 21746 9826 21758
rect 10782 21810 10834 21822
rect 10782 21746 10834 21758
rect 17390 21810 17442 21822
rect 17390 21746 17442 21758
rect 17502 21810 17554 21822
rect 17502 21746 17554 21758
rect 18398 21810 18450 21822
rect 18398 21746 18450 21758
rect 18734 21810 18786 21822
rect 25342 21810 25394 21822
rect 24322 21758 24334 21810
rect 24386 21758 24398 21810
rect 18734 21746 18786 21758
rect 25342 21746 25394 21758
rect 27358 21810 27410 21822
rect 27358 21746 27410 21758
rect 30382 21810 30434 21822
rect 30382 21746 30434 21758
rect 32174 21810 32226 21822
rect 32174 21746 32226 21758
rect 33518 21810 33570 21822
rect 33518 21746 33570 21758
rect 42254 21810 42306 21822
rect 42254 21746 42306 21758
rect 46622 21810 46674 21822
rect 46622 21746 46674 21758
rect 6974 21698 7026 21710
rect 6974 21634 7026 21646
rect 11118 21698 11170 21710
rect 11118 21634 11170 21646
rect 17614 21698 17666 21710
rect 17614 21634 17666 21646
rect 17726 21698 17778 21710
rect 17726 21634 17778 21646
rect 18510 21698 18562 21710
rect 18510 21634 18562 21646
rect 19406 21698 19458 21710
rect 19406 21634 19458 21646
rect 19518 21698 19570 21710
rect 21646 21698 21698 21710
rect 20514 21646 20526 21698
rect 20578 21646 20590 21698
rect 21186 21646 21198 21698
rect 21250 21646 21262 21698
rect 19518 21634 19570 21646
rect 21646 21634 21698 21646
rect 22094 21698 22146 21710
rect 22094 21634 22146 21646
rect 22206 21698 22258 21710
rect 25118 21698 25170 21710
rect 30494 21698 30546 21710
rect 23650 21646 23662 21698
rect 23714 21646 23726 21698
rect 23986 21646 23998 21698
rect 24050 21646 24062 21698
rect 26674 21646 26686 21698
rect 26738 21646 26750 21698
rect 29026 21646 29038 21698
rect 29090 21646 29102 21698
rect 22206 21634 22258 21646
rect 25118 21634 25170 21646
rect 30494 21634 30546 21646
rect 32398 21698 32450 21710
rect 32398 21634 32450 21646
rect 37326 21698 37378 21710
rect 37326 21634 37378 21646
rect 37886 21698 37938 21710
rect 37886 21634 37938 21646
rect 41134 21698 41186 21710
rect 47518 21698 47570 21710
rect 44034 21646 44046 21698
rect 44098 21646 44110 21698
rect 41134 21634 41186 21646
rect 47518 21634 47570 21646
rect 47854 21698 47906 21710
rect 47854 21634 47906 21646
rect 5294 21586 5346 21598
rect 4722 21534 4734 21586
rect 4786 21534 4798 21586
rect 5294 21522 5346 21534
rect 5518 21586 5570 21598
rect 5518 21522 5570 21534
rect 7870 21586 7922 21598
rect 7870 21522 7922 21534
rect 8206 21586 8258 21598
rect 8206 21522 8258 21534
rect 9662 21586 9714 21598
rect 9662 21522 9714 21534
rect 9886 21586 9938 21598
rect 11678 21586 11730 21598
rect 19294 21586 19346 21598
rect 21422 21586 21474 21598
rect 10210 21534 10222 21586
rect 10274 21534 10286 21586
rect 12002 21534 12014 21586
rect 12066 21534 12078 21586
rect 15698 21534 15710 21586
rect 15762 21534 15774 21586
rect 18050 21534 18062 21586
rect 18114 21534 18126 21586
rect 18946 21534 18958 21586
rect 19010 21534 19022 21586
rect 19730 21534 19742 21586
rect 19794 21534 19806 21586
rect 20066 21534 20078 21586
rect 20130 21534 20142 21586
rect 9886 21522 9938 21534
rect 11678 21522 11730 21534
rect 19294 21522 19346 21534
rect 21422 21522 21474 21534
rect 21870 21586 21922 21598
rect 25454 21586 25506 21598
rect 31054 21586 31106 21598
rect 32510 21586 32562 21598
rect 22530 21534 22542 21586
rect 22594 21534 22606 21586
rect 23874 21534 23886 21586
rect 23938 21534 23950 21586
rect 24546 21534 24558 21586
rect 24610 21534 24622 21586
rect 26002 21534 26014 21586
rect 26066 21534 26078 21586
rect 27570 21534 27582 21586
rect 27634 21534 27646 21586
rect 29586 21534 29598 21586
rect 29650 21534 29662 21586
rect 30706 21534 30718 21586
rect 30770 21534 30782 21586
rect 31826 21534 31838 21586
rect 31890 21534 31902 21586
rect 21870 21522 21922 21534
rect 25454 21522 25506 21534
rect 31054 21522 31106 21534
rect 32510 21522 32562 21534
rect 33182 21586 33234 21598
rect 33182 21522 33234 21534
rect 33294 21586 33346 21598
rect 33294 21522 33346 21534
rect 33742 21586 33794 21598
rect 37662 21586 37714 21598
rect 46958 21586 47010 21598
rect 34178 21534 34190 21586
rect 34242 21534 34254 21586
rect 39218 21534 39230 21586
rect 39282 21534 39294 21586
rect 43250 21534 43262 21586
rect 43314 21534 43326 21586
rect 33742 21522 33794 21534
rect 37662 21522 37714 21534
rect 46958 21522 47010 21534
rect 47182 21586 47234 21598
rect 48066 21534 48078 21586
rect 48130 21534 48142 21586
rect 47182 21522 47234 21534
rect 14926 21474 14978 21486
rect 37774 21474 37826 21486
rect 39790 21474 39842 21486
rect 1922 21422 1934 21474
rect 1986 21422 1998 21474
rect 4050 21422 4062 21474
rect 4114 21422 4126 21474
rect 12786 21422 12798 21474
rect 12850 21422 12862 21474
rect 22194 21422 22206 21474
rect 22258 21422 22270 21474
rect 31490 21422 31502 21474
rect 31554 21422 31566 21474
rect 34850 21422 34862 21474
rect 34914 21422 34926 21474
rect 36978 21422 36990 21474
rect 37042 21422 37054 21474
rect 38994 21422 39006 21474
rect 39058 21422 39070 21474
rect 14926 21410 14978 21422
rect 37774 21410 37826 21422
rect 39790 21410 39842 21422
rect 40910 21474 40962 21486
rect 40910 21410 40962 21422
rect 41694 21474 41746 21486
rect 47070 21474 47122 21486
rect 46162 21422 46174 21474
rect 46226 21422 46238 21474
rect 41694 21410 41746 21422
rect 47070 21410 47122 21422
rect 5854 21362 5906 21374
rect 5854 21298 5906 21310
rect 16494 21362 16546 21374
rect 16494 21298 16546 21310
rect 41246 21362 41298 21374
rect 41246 21298 41298 21310
rect 41806 21362 41858 21374
rect 41806 21298 41858 21310
rect 1344 21194 48608 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 48608 21194
rect 1344 21108 48608 21142
rect 42814 21026 42866 21038
rect 6290 20974 6302 21026
rect 6354 20974 6366 21026
rect 10322 20974 10334 21026
rect 10386 20974 10398 21026
rect 20514 20974 20526 21026
rect 20578 20974 20590 21026
rect 42814 20962 42866 20974
rect 13022 20914 13074 20926
rect 22766 20914 22818 20926
rect 27694 20914 27746 20926
rect 33182 20914 33234 20926
rect 4834 20862 4846 20914
rect 4898 20862 4910 20914
rect 10210 20862 10222 20914
rect 10274 20862 10286 20914
rect 15698 20862 15710 20914
rect 15762 20862 15774 20914
rect 21746 20862 21758 20914
rect 21810 20862 21822 20914
rect 23314 20862 23326 20914
rect 23378 20862 23390 20914
rect 30146 20862 30158 20914
rect 30210 20862 30222 20914
rect 32050 20862 32062 20914
rect 32114 20862 32126 20914
rect 13022 20850 13074 20862
rect 22766 20850 22818 20862
rect 27694 20850 27746 20862
rect 33182 20850 33234 20862
rect 38334 20914 38386 20926
rect 44382 20914 44434 20926
rect 39218 20862 39230 20914
rect 39282 20862 39294 20914
rect 41346 20862 41358 20914
rect 41410 20862 41422 20914
rect 42466 20862 42478 20914
rect 42530 20862 42542 20914
rect 38334 20850 38386 20862
rect 44382 20850 44434 20862
rect 45054 20914 45106 20926
rect 48178 20862 48190 20914
rect 48242 20862 48254 20914
rect 45054 20850 45106 20862
rect 6078 20802 6130 20814
rect 12910 20802 12962 20814
rect 22206 20802 22258 20814
rect 2034 20750 2046 20802
rect 2098 20750 2110 20802
rect 6290 20750 6302 20802
rect 6354 20750 6366 20802
rect 6738 20750 6750 20802
rect 6802 20750 6814 20802
rect 7746 20750 7758 20802
rect 7810 20750 7822 20802
rect 8642 20750 8654 20802
rect 8706 20750 8718 20802
rect 9762 20750 9774 20802
rect 9826 20750 9838 20802
rect 18610 20750 18622 20802
rect 18674 20750 18686 20802
rect 18946 20750 18958 20802
rect 19010 20750 19022 20802
rect 20178 20750 20190 20802
rect 20242 20750 20254 20802
rect 21522 20750 21534 20802
rect 21586 20750 21598 20802
rect 6078 20738 6130 20750
rect 12910 20738 12962 20750
rect 22206 20738 22258 20750
rect 23774 20802 23826 20814
rect 23774 20738 23826 20750
rect 25342 20802 25394 20814
rect 28030 20802 28082 20814
rect 25554 20750 25566 20802
rect 25618 20750 25630 20802
rect 25342 20738 25394 20750
rect 28030 20738 28082 20750
rect 28478 20802 28530 20814
rect 32622 20802 32674 20814
rect 36990 20802 37042 20814
rect 29362 20750 29374 20802
rect 29426 20750 29438 20802
rect 31602 20750 31614 20802
rect 31666 20750 31678 20802
rect 32274 20750 32286 20802
rect 32338 20750 32350 20802
rect 33618 20750 33630 20802
rect 33682 20750 33694 20802
rect 33954 20750 33966 20802
rect 34018 20750 34030 20802
rect 35410 20750 35422 20802
rect 35474 20750 35486 20802
rect 36306 20750 36318 20802
rect 36370 20750 36382 20802
rect 28478 20738 28530 20750
rect 32622 20738 32674 20750
rect 36990 20738 37042 20750
rect 38110 20802 38162 20814
rect 38110 20738 38162 20750
rect 38446 20802 38498 20814
rect 42018 20750 42030 20802
rect 42082 20750 42094 20802
rect 45378 20750 45390 20802
rect 45442 20750 45454 20802
rect 38446 20738 38498 20750
rect 24110 20690 24162 20702
rect 2706 20638 2718 20690
rect 2770 20638 2782 20690
rect 11890 20638 11902 20690
rect 11954 20638 11966 20690
rect 12338 20638 12350 20690
rect 12402 20638 12414 20690
rect 13458 20638 13470 20690
rect 13522 20638 13534 20690
rect 15362 20638 15374 20690
rect 15426 20638 15438 20690
rect 17826 20638 17838 20690
rect 17890 20638 17902 20690
rect 19058 20638 19070 20690
rect 19122 20638 19134 20690
rect 24110 20626 24162 20638
rect 24222 20690 24274 20702
rect 24222 20626 24274 20638
rect 26126 20690 26178 20702
rect 31166 20690 31218 20702
rect 34638 20690 34690 20702
rect 37886 20690 37938 20702
rect 30594 20638 30606 20690
rect 30658 20638 30670 20690
rect 34178 20638 34190 20690
rect 34242 20638 34254 20690
rect 37314 20638 37326 20690
rect 37378 20638 37390 20690
rect 26126 20626 26178 20638
rect 31166 20626 31218 20638
rect 34638 20626 34690 20638
rect 37886 20626 37938 20638
rect 42590 20690 42642 20702
rect 46050 20638 46062 20690
rect 46114 20638 46126 20690
rect 42590 20626 42642 20638
rect 14030 20578 14082 20590
rect 14030 20514 14082 20526
rect 15038 20578 15090 20590
rect 27022 20578 27074 20590
rect 19506 20526 19518 20578
rect 19570 20526 19582 20578
rect 15038 20514 15090 20526
rect 27022 20514 27074 20526
rect 32062 20578 32114 20590
rect 32062 20514 32114 20526
rect 1344 20410 48608 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 48608 20410
rect 1344 20324 48608 20358
rect 2494 20242 2546 20254
rect 2494 20178 2546 20190
rect 3278 20242 3330 20254
rect 3278 20178 3330 20190
rect 7758 20242 7810 20254
rect 7758 20178 7810 20190
rect 9886 20242 9938 20254
rect 20302 20242 20354 20254
rect 30494 20242 30546 20254
rect 15698 20190 15710 20242
rect 15762 20190 15774 20242
rect 9886 20178 9938 20190
rect 19294 20186 19346 20198
rect 6862 20130 6914 20142
rect 6862 20066 6914 20078
rect 11118 20130 11170 20142
rect 11118 20066 11170 20078
rect 11566 20130 11618 20142
rect 11566 20066 11618 20078
rect 11902 20130 11954 20142
rect 11902 20066 11954 20078
rect 17950 20130 18002 20142
rect 17950 20066 18002 20078
rect 18622 20130 18674 20142
rect 18622 20066 18674 20078
rect 18734 20130 18786 20142
rect 18734 20066 18786 20078
rect 19182 20130 19234 20142
rect 26226 20190 26238 20242
rect 26290 20190 26302 20242
rect 20302 20178 20354 20190
rect 30494 20178 30546 20190
rect 46398 20242 46450 20254
rect 46398 20178 46450 20190
rect 47294 20242 47346 20254
rect 47294 20178 47346 20190
rect 19294 20122 19346 20134
rect 19406 20130 19458 20142
rect 19182 20066 19234 20078
rect 19406 20066 19458 20078
rect 24110 20130 24162 20142
rect 25230 20130 25282 20142
rect 24434 20078 24446 20130
rect 24498 20078 24510 20130
rect 24110 20066 24162 20078
rect 25230 20066 25282 20078
rect 25342 20130 25394 20142
rect 25342 20066 25394 20078
rect 31838 20130 31890 20142
rect 31838 20066 31890 20078
rect 34078 20130 34130 20142
rect 34078 20066 34130 20078
rect 34414 20130 34466 20142
rect 34414 20066 34466 20078
rect 34526 20130 34578 20142
rect 34526 20066 34578 20078
rect 34638 20130 34690 20142
rect 34638 20066 34690 20078
rect 35310 20130 35362 20142
rect 35310 20066 35362 20078
rect 36094 20130 36146 20142
rect 46734 20130 46786 20142
rect 38434 20078 38446 20130
rect 38498 20078 38510 20130
rect 38770 20078 38782 20130
rect 38834 20078 38846 20130
rect 42466 20078 42478 20130
rect 42530 20078 42542 20130
rect 36094 20066 36146 20078
rect 46734 20066 46786 20078
rect 47182 20130 47234 20142
rect 47182 20066 47234 20078
rect 47518 20130 47570 20142
rect 47518 20066 47570 20078
rect 47854 20130 47906 20142
rect 47854 20066 47906 20078
rect 4398 20018 4450 20030
rect 10894 20018 10946 20030
rect 16270 20018 16322 20030
rect 5730 19966 5742 20018
rect 5794 19966 5806 20018
rect 7858 19966 7870 20018
rect 7922 19966 7934 20018
rect 9874 19966 9886 20018
rect 9938 19966 9950 20018
rect 10546 19966 10558 20018
rect 10610 19966 10622 20018
rect 12114 19966 12126 20018
rect 12178 19966 12190 20018
rect 4398 19954 4450 19966
rect 10894 19954 10946 19966
rect 16270 19954 16322 19966
rect 16830 20018 16882 20030
rect 18174 20018 18226 20030
rect 17378 19966 17390 20018
rect 17442 19966 17454 20018
rect 17714 19966 17726 20018
rect 17778 19966 17790 20018
rect 16830 19954 16882 19966
rect 18174 19954 18226 19966
rect 18398 20018 18450 20030
rect 18398 19954 18450 19966
rect 19070 20018 19122 20030
rect 20190 20018 20242 20030
rect 23886 20018 23938 20030
rect 27470 20018 27522 20030
rect 31390 20018 31442 20030
rect 19842 19966 19854 20018
rect 19906 19966 19918 20018
rect 20738 19966 20750 20018
rect 20802 19966 20814 20018
rect 24322 19966 24334 20018
rect 24386 19966 24398 20018
rect 26450 19966 26462 20018
rect 26514 19966 26526 20018
rect 26786 19966 26798 20018
rect 26850 19966 26862 20018
rect 27682 19966 27694 20018
rect 27746 19966 27758 20018
rect 30146 19966 30158 20018
rect 30210 19966 30222 20018
rect 19070 19954 19122 19966
rect 20190 19954 20242 19966
rect 23886 19954 23938 19966
rect 27470 19954 27522 19966
rect 31390 19954 31442 19966
rect 32062 20018 32114 20030
rect 32062 19954 32114 19966
rect 33518 20018 33570 20030
rect 45278 20018 45330 20030
rect 37202 19966 37214 20018
rect 37266 19966 37278 20018
rect 38994 19966 39006 20018
rect 39058 19966 39070 20018
rect 41794 19966 41806 20018
rect 41858 19966 41870 20018
rect 45042 19966 45054 20018
rect 45106 19966 45118 20018
rect 33518 19954 33570 19966
rect 45278 19954 45330 19966
rect 46510 20018 46562 20030
rect 46510 19954 46562 19966
rect 46846 20018 46898 20030
rect 46846 19954 46898 19966
rect 47742 20018 47794 20030
rect 47742 19954 47794 19966
rect 2158 19906 2210 19918
rect 8094 19906 8146 19918
rect 31054 19906 31106 19918
rect 3826 19854 3838 19906
rect 3890 19854 3902 19906
rect 5282 19854 5294 19906
rect 5346 19854 5358 19906
rect 13010 19854 13022 19906
rect 13074 19854 13086 19906
rect 17826 19854 17838 19906
rect 17890 19854 17902 19906
rect 21410 19854 21422 19906
rect 21474 19854 21486 19906
rect 23538 19854 23550 19906
rect 23602 19854 23614 19906
rect 24658 19854 24670 19906
rect 24722 19854 24734 19906
rect 26898 19854 26910 19906
rect 26962 19854 26974 19906
rect 28578 19854 28590 19906
rect 28642 19903 28654 19906
rect 28914 19903 28926 19906
rect 28642 19857 28926 19903
rect 28642 19854 28654 19857
rect 28914 19854 28926 19857
rect 28978 19854 28990 19906
rect 2158 19842 2210 19854
rect 8094 19842 8146 19854
rect 31054 19842 31106 19854
rect 31950 19906 32002 19918
rect 31950 19842 32002 19854
rect 32510 19906 32562 19918
rect 32510 19842 32562 19854
rect 33182 19906 33234 19918
rect 33182 19842 33234 19854
rect 35646 19906 35698 19918
rect 35646 19842 35698 19854
rect 36542 19906 36594 19918
rect 36542 19842 36594 19854
rect 37438 19906 37490 19918
rect 37438 19842 37490 19854
rect 37886 19906 37938 19918
rect 37886 19842 37938 19854
rect 39566 19906 39618 19918
rect 39566 19842 39618 19854
rect 40014 19906 40066 19918
rect 40014 19842 40066 19854
rect 41022 19906 41074 19918
rect 44594 19854 44606 19906
rect 44658 19854 44670 19906
rect 41022 19842 41074 19854
rect 25342 19794 25394 19806
rect 32398 19794 32450 19806
rect 28018 19742 28030 19794
rect 28082 19742 28094 19794
rect 25342 19730 25394 19742
rect 32398 19730 32450 19742
rect 37550 19794 37602 19806
rect 37550 19730 37602 19742
rect 38110 19794 38162 19806
rect 47854 19794 47906 19806
rect 45042 19742 45054 19794
rect 45106 19742 45118 19794
rect 38110 19730 38162 19742
rect 47854 19730 47906 19742
rect 1344 19626 48608 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 48608 19626
rect 1344 19540 48608 19574
rect 15934 19458 15986 19470
rect 29150 19458 29202 19470
rect 27346 19406 27358 19458
rect 27410 19406 27422 19458
rect 15934 19394 15986 19406
rect 29150 19394 29202 19406
rect 43934 19458 43986 19470
rect 43934 19394 43986 19406
rect 5182 19346 5234 19358
rect 17166 19346 17218 19358
rect 1698 19294 1710 19346
rect 1762 19294 1774 19346
rect 5618 19294 5630 19346
rect 5682 19294 5694 19346
rect 11218 19294 11230 19346
rect 11282 19294 11294 19346
rect 12898 19294 12910 19346
rect 12962 19294 12974 19346
rect 5182 19282 5234 19294
rect 17166 19282 17218 19294
rect 18846 19346 18898 19358
rect 29710 19346 29762 19358
rect 35422 19346 35474 19358
rect 43710 19346 43762 19358
rect 19282 19294 19294 19346
rect 19346 19294 19358 19346
rect 20514 19294 20526 19346
rect 20578 19294 20590 19346
rect 21298 19294 21310 19346
rect 21362 19294 21374 19346
rect 24546 19294 24558 19346
rect 24610 19294 24622 19346
rect 26674 19294 26686 19346
rect 26738 19294 26750 19346
rect 28130 19294 28142 19346
rect 28194 19294 28206 19346
rect 30146 19294 30158 19346
rect 30210 19294 30222 19346
rect 30930 19294 30942 19346
rect 30994 19294 31006 19346
rect 37762 19294 37774 19346
rect 37826 19294 37838 19346
rect 39890 19294 39902 19346
rect 39954 19294 39966 19346
rect 40226 19294 40238 19346
rect 40290 19294 40302 19346
rect 48178 19294 48190 19346
rect 48242 19294 48254 19346
rect 18846 19282 18898 19294
rect 29710 19282 29762 19294
rect 35422 19282 35474 19294
rect 43710 19282 43762 19294
rect 13694 19234 13746 19246
rect 16382 19234 16434 19246
rect 4498 19182 4510 19234
rect 4562 19182 4574 19234
rect 7074 19182 7086 19234
rect 7138 19182 7150 19234
rect 8418 19182 8430 19234
rect 8482 19182 8494 19234
rect 15250 19182 15262 19234
rect 15314 19182 15326 19234
rect 13694 19170 13746 19182
rect 16382 19170 16434 19182
rect 16718 19234 16770 19246
rect 16718 19170 16770 19182
rect 16942 19234 16994 19246
rect 16942 19170 16994 19182
rect 18622 19234 18674 19246
rect 18622 19170 18674 19182
rect 19742 19234 19794 19246
rect 22094 19234 22146 19246
rect 29486 19234 29538 19246
rect 20178 19182 20190 19234
rect 20242 19182 20254 19234
rect 21410 19182 21422 19234
rect 21474 19182 21486 19234
rect 23314 19182 23326 19234
rect 23378 19182 23390 19234
rect 23874 19182 23886 19234
rect 23938 19182 23950 19234
rect 27570 19182 27582 19234
rect 27634 19182 27646 19234
rect 27906 19182 27918 19234
rect 27970 19182 27982 19234
rect 30482 19182 30494 19234
rect 30546 19182 30558 19234
rect 33842 19182 33854 19234
rect 33906 19182 33918 19234
rect 36978 19182 36990 19234
rect 37042 19182 37054 19234
rect 43026 19182 43038 19234
rect 43090 19182 43102 19234
rect 45378 19182 45390 19234
rect 45442 19182 45454 19234
rect 19742 19170 19794 19182
rect 22094 19170 22146 19182
rect 29486 19170 29538 19182
rect 6078 19122 6130 19134
rect 3826 19070 3838 19122
rect 3890 19070 3902 19122
rect 5954 19070 5966 19122
rect 6018 19070 6030 19122
rect 6078 19058 6130 19070
rect 6190 19122 6242 19134
rect 6190 19058 6242 19070
rect 7534 19122 7586 19134
rect 7534 19058 7586 19070
rect 7646 19122 7698 19134
rect 7646 19058 7698 19070
rect 7758 19122 7810 19134
rect 11678 19122 11730 19134
rect 9090 19070 9102 19122
rect 9154 19070 9166 19122
rect 7758 19058 7810 19070
rect 11678 19058 11730 19070
rect 12462 19122 12514 19134
rect 21758 19122 21810 19134
rect 34526 19122 34578 19134
rect 12562 19070 12574 19122
rect 12626 19070 12638 19122
rect 15474 19070 15486 19122
rect 15538 19070 15550 19122
rect 22754 19070 22766 19122
rect 22818 19070 22830 19122
rect 23090 19070 23102 19122
rect 23154 19070 23166 19122
rect 33058 19070 33070 19122
rect 33122 19070 33134 19122
rect 34178 19070 34190 19122
rect 34242 19070 34254 19122
rect 12462 19058 12514 19070
rect 21758 19058 21810 19070
rect 34526 19058 34578 19070
rect 34974 19122 35026 19134
rect 42354 19070 42366 19122
rect 42418 19070 42430 19122
rect 46050 19070 46062 19122
rect 46114 19070 46126 19122
rect 34974 19058 35026 19070
rect 6414 19010 6466 19022
rect 6414 18946 6466 18958
rect 7870 19010 7922 19022
rect 7870 18946 7922 18958
rect 11790 19010 11842 19022
rect 11790 18946 11842 18958
rect 12126 19010 12178 19022
rect 12126 18946 12178 18958
rect 12350 19010 12402 19022
rect 12350 18946 12402 18958
rect 16494 19010 16546 19022
rect 16494 18946 16546 18958
rect 17502 19010 17554 19022
rect 17502 18946 17554 18958
rect 18174 19010 18226 19022
rect 18174 18946 18226 18958
rect 18286 19010 18338 19022
rect 18286 18946 18338 18958
rect 18398 19010 18450 19022
rect 18398 18946 18450 18958
rect 21870 19010 21922 19022
rect 21870 18946 21922 18958
rect 22430 19010 22482 19022
rect 22430 18946 22482 18958
rect 34862 19010 34914 19022
rect 34862 18946 34914 18958
rect 35870 19010 35922 19022
rect 35870 18946 35922 18958
rect 36318 19010 36370 19022
rect 45054 19010 45106 19022
rect 44258 18958 44270 19010
rect 44322 18958 44334 19010
rect 36318 18946 36370 18958
rect 45054 18946 45106 18958
rect 1344 18842 48608 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 48608 18842
rect 1344 18756 48608 18790
rect 6526 18674 6578 18686
rect 5842 18622 5854 18674
rect 5906 18622 5918 18674
rect 6526 18610 6578 18622
rect 7086 18674 7138 18686
rect 24110 18674 24162 18686
rect 18498 18622 18510 18674
rect 18562 18622 18574 18674
rect 7086 18610 7138 18622
rect 24110 18610 24162 18622
rect 31502 18674 31554 18686
rect 31502 18610 31554 18622
rect 33070 18674 33122 18686
rect 33070 18610 33122 18622
rect 38110 18674 38162 18686
rect 38110 18610 38162 18622
rect 38894 18674 38946 18686
rect 38894 18610 38946 18622
rect 45166 18674 45218 18686
rect 45166 18610 45218 18622
rect 46174 18674 46226 18686
rect 46174 18610 46226 18622
rect 7310 18562 7362 18574
rect 7310 18498 7362 18510
rect 7422 18562 7474 18574
rect 20862 18562 20914 18574
rect 7634 18510 7646 18562
rect 7698 18510 7710 18562
rect 7422 18498 7474 18510
rect 20862 18498 20914 18510
rect 21198 18562 21250 18574
rect 31838 18562 31890 18574
rect 38334 18562 38386 18574
rect 22866 18510 22878 18562
rect 22930 18510 22942 18562
rect 23538 18510 23550 18562
rect 23602 18510 23614 18562
rect 24434 18510 24446 18562
rect 24498 18510 24510 18562
rect 32498 18510 32510 18562
rect 32562 18510 32574 18562
rect 33394 18510 33406 18562
rect 33458 18510 33470 18562
rect 21198 18498 21250 18510
rect 31838 18498 31890 18510
rect 38334 18498 38386 18510
rect 39006 18562 39058 18574
rect 39006 18498 39058 18510
rect 44494 18562 44546 18574
rect 47070 18562 47122 18574
rect 45490 18510 45502 18562
rect 45554 18510 45566 18562
rect 44494 18498 44546 18510
rect 47070 18498 47122 18510
rect 47854 18562 47906 18574
rect 47854 18498 47906 18510
rect 2046 18450 2098 18462
rect 12574 18450 12626 18462
rect 18846 18450 18898 18462
rect 2482 18398 2494 18450
rect 2546 18398 2558 18450
rect 6514 18398 6526 18450
rect 6578 18398 6590 18450
rect 8642 18398 8654 18450
rect 8706 18398 8718 18450
rect 9650 18398 9662 18450
rect 9714 18398 9726 18450
rect 12786 18398 12798 18450
rect 12850 18398 12862 18450
rect 13906 18398 13918 18450
rect 13970 18398 13982 18450
rect 14578 18398 14590 18450
rect 14642 18398 14654 18450
rect 17602 18398 17614 18450
rect 17666 18398 17678 18450
rect 18050 18398 18062 18450
rect 18114 18398 18126 18450
rect 2046 18386 2098 18398
rect 12574 18386 12626 18398
rect 18846 18386 18898 18398
rect 19630 18450 19682 18462
rect 19630 18386 19682 18398
rect 19854 18450 19906 18462
rect 19854 18386 19906 18398
rect 20302 18450 20354 18462
rect 23886 18450 23938 18462
rect 29038 18450 29090 18462
rect 30382 18450 30434 18462
rect 31166 18450 31218 18462
rect 21410 18398 21422 18450
rect 21474 18398 21486 18450
rect 22754 18398 22766 18450
rect 22818 18398 22830 18450
rect 23314 18398 23326 18450
rect 23378 18398 23390 18450
rect 24322 18398 24334 18450
rect 24386 18398 24398 18450
rect 25330 18398 25342 18450
rect 25394 18398 25406 18450
rect 29586 18398 29598 18450
rect 29650 18398 29662 18450
rect 30818 18398 30830 18450
rect 30882 18398 30894 18450
rect 20302 18386 20354 18398
rect 23886 18386 23938 18398
rect 29038 18386 29090 18398
rect 30382 18386 30434 18398
rect 31166 18386 31218 18398
rect 31502 18450 31554 18462
rect 31502 18386 31554 18398
rect 32174 18450 32226 18462
rect 37662 18450 37714 18462
rect 33842 18398 33854 18450
rect 33906 18398 33918 18450
rect 32174 18386 32226 18398
rect 37662 18386 37714 18398
rect 38222 18450 38274 18462
rect 45950 18450 46002 18462
rect 39666 18398 39678 18450
rect 39730 18398 39742 18450
rect 40898 18398 40910 18450
rect 40962 18398 40974 18450
rect 43810 18398 43822 18450
rect 43874 18398 43886 18450
rect 44706 18398 44718 18450
rect 44770 18398 44782 18450
rect 38222 18386 38274 18398
rect 45950 18386 46002 18398
rect 46174 18450 46226 18462
rect 46174 18386 46226 18398
rect 46398 18450 46450 18462
rect 46398 18386 46450 18398
rect 46734 18450 46786 18462
rect 46734 18386 46786 18398
rect 46846 18450 46898 18462
rect 46846 18386 46898 18398
rect 47182 18450 47234 18462
rect 48066 18398 48078 18450
rect 48130 18398 48142 18450
rect 47182 18386 47234 18398
rect 7198 18338 7250 18350
rect 19406 18338 19458 18350
rect 3154 18286 3166 18338
rect 3218 18286 3230 18338
rect 10882 18286 10894 18338
rect 10946 18286 10958 18338
rect 16706 18286 16718 18338
rect 16770 18286 16782 18338
rect 7198 18274 7250 18286
rect 19406 18274 19458 18286
rect 19742 18338 19794 18350
rect 37102 18338 37154 18350
rect 40350 18338 40402 18350
rect 22530 18286 22542 18338
rect 22594 18286 22606 18338
rect 24658 18286 24670 18338
rect 24722 18286 24734 18338
rect 26002 18286 26014 18338
rect 26066 18286 26078 18338
rect 28130 18286 28142 18338
rect 28194 18286 28206 18338
rect 28578 18286 28590 18338
rect 28642 18286 28654 18338
rect 29922 18286 29934 18338
rect 29986 18286 29998 18338
rect 34514 18286 34526 18338
rect 34578 18286 34590 18338
rect 36642 18286 36654 18338
rect 36706 18286 36718 18338
rect 39442 18286 39454 18338
rect 39506 18286 39518 18338
rect 42018 18286 42030 18338
rect 42082 18286 42094 18338
rect 19742 18274 19794 18286
rect 37102 18274 37154 18286
rect 40350 18274 40402 18286
rect 19182 18226 19234 18238
rect 8418 18174 8430 18226
rect 8482 18174 8494 18226
rect 13234 18174 13246 18226
rect 13298 18174 13310 18226
rect 18050 18174 18062 18226
rect 18114 18174 18126 18226
rect 19182 18162 19234 18174
rect 38894 18226 38946 18238
rect 38894 18162 38946 18174
rect 43822 18226 43874 18238
rect 43822 18162 43874 18174
rect 44158 18226 44210 18238
rect 44158 18162 44210 18174
rect 1344 18058 48608 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 48608 18058
rect 1344 17972 48608 18006
rect 20638 17890 20690 17902
rect 20638 17826 20690 17838
rect 23774 17890 23826 17902
rect 46398 17890 46450 17902
rect 43362 17838 43374 17890
rect 43426 17838 43438 17890
rect 23774 17826 23826 17838
rect 46398 17826 46450 17838
rect 25566 17778 25618 17790
rect 35086 17778 35138 17790
rect 42926 17778 42978 17790
rect 1922 17726 1934 17778
rect 1986 17726 1998 17778
rect 4610 17726 4622 17778
rect 4674 17726 4686 17778
rect 6290 17726 6302 17778
rect 6354 17726 6366 17778
rect 11106 17726 11118 17778
rect 11170 17726 11182 17778
rect 12898 17726 12910 17778
rect 12962 17726 12974 17778
rect 14130 17726 14142 17778
rect 14194 17726 14206 17778
rect 27122 17726 27134 17778
rect 27186 17726 27198 17778
rect 32946 17726 32958 17778
rect 33010 17726 33022 17778
rect 34626 17726 34638 17778
rect 34690 17726 34702 17778
rect 38434 17726 38446 17778
rect 38498 17726 38510 17778
rect 25566 17714 25618 17726
rect 35086 17714 35138 17726
rect 42926 17714 42978 17726
rect 44046 17778 44098 17790
rect 44046 17714 44098 17726
rect 47854 17778 47906 17790
rect 47854 17714 47906 17726
rect 3726 17666 3778 17678
rect 2258 17614 2270 17666
rect 2322 17614 2334 17666
rect 3726 17602 3778 17614
rect 5070 17666 5122 17678
rect 14926 17666 14978 17678
rect 17390 17666 17442 17678
rect 6626 17614 6638 17666
rect 6690 17614 6702 17666
rect 8194 17614 8206 17666
rect 8258 17614 8270 17666
rect 17042 17614 17054 17666
rect 17106 17614 17118 17666
rect 5070 17602 5122 17614
rect 14926 17602 14978 17614
rect 17390 17602 17442 17614
rect 19406 17666 19458 17678
rect 19406 17602 19458 17614
rect 19630 17666 19682 17678
rect 19630 17602 19682 17614
rect 19966 17666 20018 17678
rect 19966 17602 20018 17614
rect 20526 17666 20578 17678
rect 23886 17666 23938 17678
rect 21634 17614 21646 17666
rect 21698 17614 21710 17666
rect 22418 17614 22430 17666
rect 22482 17614 22494 17666
rect 23090 17614 23102 17666
rect 23154 17614 23166 17666
rect 20526 17602 20578 17614
rect 23886 17602 23938 17614
rect 24670 17666 24722 17678
rect 24670 17602 24722 17614
rect 25006 17666 25058 17678
rect 25006 17602 25058 17614
rect 25902 17666 25954 17678
rect 25902 17602 25954 17614
rect 28030 17666 28082 17678
rect 28030 17602 28082 17614
rect 28590 17666 28642 17678
rect 28590 17602 28642 17614
rect 29150 17666 29202 17678
rect 33294 17666 33346 17678
rect 30146 17614 30158 17666
rect 30210 17614 30222 17666
rect 29150 17602 29202 17614
rect 33294 17602 33346 17614
rect 33854 17666 33906 17678
rect 35646 17666 35698 17678
rect 34514 17614 34526 17666
rect 34578 17614 34590 17666
rect 33854 17602 33906 17614
rect 35646 17602 35698 17614
rect 35758 17666 35810 17678
rect 35758 17602 35810 17614
rect 35982 17666 36034 17678
rect 44718 17666 44770 17678
rect 38994 17614 39006 17666
rect 39058 17614 39070 17666
rect 41906 17614 41918 17666
rect 41970 17614 41982 17666
rect 43026 17614 43038 17666
rect 43090 17614 43102 17666
rect 43362 17614 43374 17666
rect 43426 17614 43438 17666
rect 35982 17602 36034 17614
rect 44718 17602 44770 17614
rect 45390 17666 45442 17678
rect 45390 17602 45442 17614
rect 46734 17666 46786 17678
rect 46734 17602 46786 17614
rect 3950 17554 4002 17566
rect 3950 17490 4002 17502
rect 6302 17554 6354 17566
rect 7534 17554 7586 17566
rect 7298 17502 7310 17554
rect 7362 17502 7374 17554
rect 6302 17490 6354 17502
rect 7534 17490 7586 17502
rect 7758 17554 7810 17566
rect 7758 17490 7810 17502
rect 7870 17554 7922 17566
rect 12462 17554 12514 17566
rect 14590 17554 14642 17566
rect 8978 17502 8990 17554
rect 9042 17502 9054 17554
rect 11778 17502 11790 17554
rect 11842 17502 11854 17554
rect 12562 17502 12574 17554
rect 12626 17502 12638 17554
rect 14354 17502 14366 17554
rect 14418 17502 14430 17554
rect 7870 17490 7922 17502
rect 12462 17490 12514 17502
rect 14590 17490 14642 17502
rect 14702 17554 14754 17566
rect 17950 17554 18002 17566
rect 15362 17502 15374 17554
rect 15426 17502 15438 17554
rect 14702 17490 14754 17502
rect 17950 17490 18002 17502
rect 19854 17554 19906 17566
rect 26014 17554 26066 17566
rect 21858 17502 21870 17554
rect 21922 17502 21934 17554
rect 22194 17502 22206 17554
rect 22258 17502 22270 17554
rect 23314 17502 23326 17554
rect 23378 17502 23390 17554
rect 19854 17490 19906 17502
rect 26014 17490 26066 17502
rect 27358 17554 27410 17566
rect 28478 17554 28530 17566
rect 27682 17502 27694 17554
rect 27746 17502 27758 17554
rect 27358 17490 27410 17502
rect 28478 17490 28530 17502
rect 29486 17554 29538 17566
rect 33406 17554 33458 17566
rect 30818 17502 30830 17554
rect 30882 17502 30894 17554
rect 29486 17490 29538 17502
rect 33406 17490 33458 17502
rect 33630 17554 33682 17566
rect 33630 17490 33682 17502
rect 34078 17554 34130 17566
rect 34078 17490 34130 17502
rect 34190 17554 34242 17566
rect 34190 17490 34242 17502
rect 36094 17554 36146 17566
rect 42814 17554 42866 17566
rect 40674 17502 40686 17554
rect 40738 17502 40750 17554
rect 36094 17490 36146 17502
rect 42814 17490 42866 17502
rect 45166 17554 45218 17566
rect 45166 17490 45218 17502
rect 45614 17554 45666 17566
rect 45614 17490 45666 17502
rect 45950 17554 46002 17566
rect 45950 17490 46002 17502
rect 46286 17554 46338 17566
rect 46286 17490 46338 17502
rect 46958 17554 47010 17566
rect 46958 17490 47010 17502
rect 47070 17554 47122 17566
rect 47506 17502 47518 17554
rect 47570 17502 47582 17554
rect 47070 17490 47122 17502
rect 3278 17442 3330 17454
rect 3278 17378 3330 17390
rect 3502 17442 3554 17454
rect 3502 17378 3554 17390
rect 3614 17442 3666 17454
rect 3614 17378 3666 17390
rect 5966 17442 6018 17454
rect 5966 17378 6018 17390
rect 6190 17442 6242 17454
rect 6190 17378 6242 17390
rect 7646 17442 7698 17454
rect 7646 17378 7698 17390
rect 11454 17442 11506 17454
rect 11454 17378 11506 17390
rect 12126 17442 12178 17454
rect 12126 17378 12178 17390
rect 12350 17442 12402 17454
rect 12350 17378 12402 17390
rect 13470 17442 13522 17454
rect 20078 17442 20130 17454
rect 13794 17390 13806 17442
rect 13858 17390 13870 17442
rect 16930 17390 16942 17442
rect 16994 17390 17006 17442
rect 13470 17378 13522 17390
rect 20078 17378 20130 17390
rect 20638 17442 20690 17454
rect 20638 17378 20690 17390
rect 23774 17442 23826 17454
rect 26686 17442 26738 17454
rect 24322 17390 24334 17442
rect 24386 17390 24398 17442
rect 26338 17390 26350 17442
rect 26402 17390 26414 17442
rect 23774 17378 23826 17390
rect 26686 17378 26738 17390
rect 28254 17442 28306 17454
rect 28254 17378 28306 17390
rect 44942 17442 44994 17454
rect 44942 17378 44994 17390
rect 45838 17442 45890 17454
rect 45838 17378 45890 17390
rect 46398 17442 46450 17454
rect 46398 17378 46450 17390
rect 1344 17274 48608 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 48608 17274
rect 1344 17188 48608 17222
rect 1710 17106 1762 17118
rect 1710 17042 1762 17054
rect 2718 17106 2770 17118
rect 2718 17042 2770 17054
rect 3726 17106 3778 17118
rect 4510 17106 4562 17118
rect 3726 17042 3778 17054
rect 4062 17050 4114 17062
rect 3166 16994 3218 17006
rect 4510 17042 4562 17054
rect 5518 17106 5570 17118
rect 5518 17042 5570 17054
rect 10558 17106 10610 17118
rect 10558 17042 10610 17054
rect 10782 17106 10834 17118
rect 10782 17042 10834 17054
rect 17390 17106 17442 17118
rect 17390 17042 17442 17054
rect 18622 17106 18674 17118
rect 18622 17042 18674 17054
rect 22430 17106 22482 17118
rect 22430 17042 22482 17054
rect 24334 17106 24386 17118
rect 24334 17042 24386 17054
rect 24558 17106 24610 17118
rect 29486 17106 29538 17118
rect 29138 17054 29150 17106
rect 29202 17054 29214 17106
rect 24558 17042 24610 17054
rect 29486 17042 29538 17054
rect 29822 17106 29874 17118
rect 29822 17042 29874 17054
rect 30830 17106 30882 17118
rect 30830 17042 30882 17054
rect 31950 17106 32002 17118
rect 31950 17042 32002 17054
rect 32174 17106 32226 17118
rect 40226 17054 40238 17106
rect 40290 17054 40302 17106
rect 32174 17042 32226 17054
rect 4062 16986 4114 16998
rect 24670 16994 24722 17006
rect 27022 16994 27074 17006
rect 30718 16994 30770 17006
rect 47966 16994 48018 17006
rect 3166 16930 3218 16942
rect 26226 16942 26238 16994
rect 26290 16942 26302 16994
rect 28354 16942 28366 16994
rect 28418 16942 28430 16994
rect 44930 16942 44942 16994
rect 44994 16942 45006 16994
rect 24670 16930 24722 16942
rect 27022 16930 27074 16942
rect 30718 16930 30770 16942
rect 47966 16930 48018 16942
rect 2270 16882 2322 16894
rect 2270 16818 2322 16830
rect 2606 16882 2658 16894
rect 2606 16818 2658 16830
rect 2830 16882 2882 16894
rect 2830 16818 2882 16830
rect 4174 16882 4226 16894
rect 9550 16882 9602 16894
rect 10446 16882 10498 16894
rect 17614 16882 17666 16894
rect 5842 16830 5854 16882
rect 5906 16830 5918 16882
rect 6626 16830 6638 16882
rect 6690 16830 6702 16882
rect 9986 16830 9998 16882
rect 10050 16830 10062 16882
rect 13794 16830 13806 16882
rect 13858 16830 13870 16882
rect 14802 16830 14814 16882
rect 14866 16830 14878 16882
rect 4174 16818 4226 16830
rect 9550 16818 9602 16830
rect 10446 16818 10498 16830
rect 17614 16818 17666 16830
rect 18062 16882 18114 16894
rect 18062 16818 18114 16830
rect 18398 16882 18450 16894
rect 18398 16818 18450 16830
rect 19070 16882 19122 16894
rect 22542 16882 22594 16894
rect 25790 16882 25842 16894
rect 20066 16830 20078 16882
rect 20130 16830 20142 16882
rect 23426 16830 23438 16882
rect 23490 16830 23502 16882
rect 23762 16830 23774 16882
rect 23826 16830 23838 16882
rect 19070 16818 19122 16830
rect 22542 16818 22594 16830
rect 25790 16818 25842 16830
rect 26574 16882 26626 16894
rect 26574 16818 26626 16830
rect 26910 16882 26962 16894
rect 26910 16818 26962 16830
rect 27246 16882 27298 16894
rect 27246 16818 27298 16830
rect 28702 16882 28754 16894
rect 28702 16818 28754 16830
rect 30942 16882 30994 16894
rect 30942 16818 30994 16830
rect 31278 16882 31330 16894
rect 31278 16818 31330 16830
rect 31502 16882 31554 16894
rect 31502 16818 31554 16830
rect 32062 16882 32114 16894
rect 36094 16882 36146 16894
rect 47294 16882 47346 16894
rect 33058 16830 33070 16882
rect 33122 16830 33134 16882
rect 36530 16830 36542 16882
rect 36594 16830 36606 16882
rect 40898 16830 40910 16882
rect 40962 16830 40974 16882
rect 44146 16830 44158 16882
rect 44210 16830 44222 16882
rect 32062 16818 32114 16830
rect 36094 16818 36146 16830
rect 47294 16818 47346 16830
rect 47518 16882 47570 16894
rect 47518 16818 47570 16830
rect 47742 16882 47794 16894
rect 47742 16818 47794 16830
rect 17502 16770 17554 16782
rect 4946 16718 4958 16770
rect 5010 16718 5022 16770
rect 8754 16718 8766 16770
rect 8818 16718 8830 16770
rect 10994 16718 11006 16770
rect 11058 16718 11070 16770
rect 13122 16718 13134 16770
rect 13186 16718 13198 16770
rect 15362 16718 15374 16770
rect 15426 16718 15438 16770
rect 17502 16706 17554 16718
rect 18510 16770 18562 16782
rect 18510 16706 18562 16718
rect 18846 16770 18898 16782
rect 25230 16770 25282 16782
rect 20962 16718 20974 16770
rect 21026 16718 21038 16770
rect 23202 16718 23214 16770
rect 23266 16718 23278 16770
rect 18846 16706 18898 16718
rect 25230 16706 25282 16718
rect 27582 16770 27634 16782
rect 27582 16706 27634 16718
rect 27694 16770 27746 16782
rect 27694 16706 27746 16718
rect 30382 16770 30434 16782
rect 39678 16770 39730 16782
rect 35410 16718 35422 16770
rect 35474 16718 35486 16770
rect 37202 16718 37214 16770
rect 37266 16718 37278 16770
rect 39330 16718 39342 16770
rect 39394 16718 39406 16770
rect 41682 16718 41694 16770
rect 41746 16718 41758 16770
rect 43810 16718 43822 16770
rect 43874 16718 43886 16770
rect 47058 16718 47070 16770
rect 47122 16718 47134 16770
rect 30382 16706 30434 16718
rect 39678 16706 39730 16718
rect 4062 16658 4114 16670
rect 27918 16658 27970 16670
rect 22978 16606 22990 16658
rect 23042 16606 23054 16658
rect 4062 16594 4114 16606
rect 27918 16594 27970 16606
rect 28030 16658 28082 16670
rect 28030 16594 28082 16606
rect 39902 16658 39954 16670
rect 39902 16594 39954 16606
rect 1344 16490 48608 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 48608 16490
rect 1344 16404 48608 16438
rect 4398 16322 4450 16334
rect 4398 16258 4450 16270
rect 12686 16322 12738 16334
rect 12686 16258 12738 16270
rect 16494 16322 16546 16334
rect 16494 16258 16546 16270
rect 21422 16322 21474 16334
rect 21422 16258 21474 16270
rect 27022 16322 27074 16334
rect 27022 16258 27074 16270
rect 2158 16210 2210 16222
rect 2158 16146 2210 16158
rect 3166 16210 3218 16222
rect 3166 16146 3218 16158
rect 4062 16210 4114 16222
rect 4062 16146 4114 16158
rect 6078 16210 6130 16222
rect 6078 16146 6130 16158
rect 7870 16210 7922 16222
rect 23886 16210 23938 16222
rect 31390 16210 31442 16222
rect 37102 16210 37154 16222
rect 41806 16210 41858 16222
rect 8306 16158 8318 16210
rect 8370 16158 8382 16210
rect 13906 16158 13918 16210
rect 13970 16158 13982 16210
rect 23426 16158 23438 16210
rect 23490 16158 23502 16210
rect 26674 16158 26686 16210
rect 26738 16158 26750 16210
rect 33058 16158 33070 16210
rect 33122 16158 33134 16210
rect 36418 16158 36430 16210
rect 36482 16158 36494 16210
rect 39218 16158 39230 16210
rect 39282 16158 39294 16210
rect 41346 16158 41358 16210
rect 41410 16158 41422 16210
rect 7870 16146 7922 16158
rect 23886 16146 23938 16158
rect 31390 16146 31442 16158
rect 37102 16146 37154 16158
rect 41806 16146 41858 16158
rect 42702 16210 42754 16222
rect 46050 16158 46062 16210
rect 46114 16158 46126 16210
rect 48178 16158 48190 16210
rect 48242 16158 48254 16210
rect 42702 16146 42754 16158
rect 5182 16098 5234 16110
rect 7310 16098 7362 16110
rect 11902 16098 11954 16110
rect 17054 16098 17106 16110
rect 24222 16098 24274 16110
rect 6738 16046 6750 16098
rect 6802 16046 6814 16098
rect 11218 16046 11230 16098
rect 11282 16046 11294 16098
rect 16034 16046 16046 16098
rect 16098 16046 16110 16098
rect 20738 16046 20750 16098
rect 20802 16046 20814 16098
rect 23090 16046 23102 16098
rect 23154 16046 23166 16098
rect 5182 16034 5234 16046
rect 7310 16034 7362 16046
rect 11902 16034 11954 16046
rect 17054 16034 17106 16046
rect 24222 16034 24274 16046
rect 24558 16098 24610 16110
rect 24558 16034 24610 16046
rect 25566 16098 25618 16110
rect 28254 16098 28306 16110
rect 30270 16098 30322 16110
rect 37886 16098 37938 16110
rect 42366 16098 42418 16110
rect 27682 16046 27694 16098
rect 27746 16046 27758 16098
rect 29586 16046 29598 16098
rect 29650 16046 29662 16098
rect 30818 16046 30830 16098
rect 30882 16046 30894 16098
rect 33618 16046 33630 16098
rect 33682 16046 33694 16098
rect 38434 16046 38446 16098
rect 38498 16046 38510 16098
rect 25566 16034 25618 16046
rect 28254 16034 28306 16046
rect 30270 16034 30322 16046
rect 37886 16034 37938 16046
rect 42366 16034 42418 16046
rect 42926 16098 42978 16110
rect 42926 16034 42978 16046
rect 43150 16098 43202 16110
rect 43150 16034 43202 16046
rect 43486 16098 43538 16110
rect 43486 16034 43538 16046
rect 43822 16098 43874 16110
rect 45378 16046 45390 16098
rect 45442 16046 45454 16098
rect 43822 16034 43874 16046
rect 4286 15986 4338 15998
rect 4286 15922 4338 15934
rect 4398 15986 4450 15998
rect 4398 15922 4450 15934
rect 4846 15986 4898 15998
rect 4846 15922 4898 15934
rect 6302 15986 6354 15998
rect 16382 15986 16434 15998
rect 10434 15934 10446 15986
rect 10498 15934 10510 15986
rect 6302 15922 6354 15934
rect 16382 15922 16434 15934
rect 16494 15986 16546 15998
rect 16494 15922 16546 15934
rect 17614 15986 17666 15998
rect 17614 15922 17666 15934
rect 19630 15986 19682 15998
rect 19630 15922 19682 15934
rect 21310 15986 21362 15998
rect 21310 15922 21362 15934
rect 21758 15986 21810 15998
rect 21758 15922 21810 15934
rect 22094 15986 22146 15998
rect 22094 15922 22146 15934
rect 22318 15986 22370 15998
rect 22318 15922 22370 15934
rect 23998 15986 24050 15998
rect 23998 15922 24050 15934
rect 24446 15986 24498 15998
rect 25902 15986 25954 15998
rect 25218 15934 25230 15986
rect 25282 15934 25294 15986
rect 24446 15922 24498 15934
rect 25902 15922 25954 15934
rect 26126 15986 26178 15998
rect 26126 15922 26178 15934
rect 26798 15986 26850 15998
rect 32622 15986 32674 15998
rect 37662 15986 37714 15998
rect 29362 15934 29374 15986
rect 29426 15934 29438 15986
rect 34290 15934 34302 15986
rect 34354 15934 34366 15986
rect 26798 15922 26850 15934
rect 32622 15922 32674 15934
rect 37662 15922 37714 15934
rect 38110 15986 38162 15998
rect 38110 15922 38162 15934
rect 41694 15986 41746 15998
rect 41694 15922 41746 15934
rect 42590 15986 42642 15998
rect 42590 15922 42642 15934
rect 43710 15986 43762 15998
rect 43710 15922 43762 15934
rect 2718 15874 2770 15886
rect 2718 15810 2770 15822
rect 3502 15874 3554 15886
rect 3502 15810 3554 15822
rect 4958 15874 5010 15886
rect 4958 15810 5010 15822
rect 5966 15874 6018 15886
rect 5966 15810 6018 15822
rect 6190 15874 6242 15886
rect 21982 15874 22034 15886
rect 19730 15822 19742 15874
rect 19794 15822 19806 15874
rect 6190 15810 6242 15822
rect 21982 15810 22034 15822
rect 24894 15874 24946 15886
rect 24894 15810 24946 15822
rect 25790 15874 25842 15886
rect 30382 15874 30434 15886
rect 27906 15822 27918 15874
rect 27970 15822 27982 15874
rect 28578 15822 28590 15874
rect 28642 15822 28654 15874
rect 25790 15810 25842 15822
rect 30382 15810 30434 15822
rect 30494 15874 30546 15886
rect 30494 15810 30546 15822
rect 31726 15874 31778 15886
rect 31726 15810 31778 15822
rect 31950 15874 32002 15886
rect 31950 15810 32002 15822
rect 32062 15874 32114 15886
rect 32062 15810 32114 15822
rect 32174 15874 32226 15886
rect 32174 15810 32226 15822
rect 37998 15874 38050 15886
rect 37998 15810 38050 15822
rect 41918 15874 41970 15886
rect 41918 15810 41970 15822
rect 1344 15706 48608 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 48608 15706
rect 1344 15620 48608 15654
rect 2158 15538 2210 15550
rect 2158 15474 2210 15486
rect 3502 15538 3554 15550
rect 8430 15538 8482 15550
rect 16270 15538 16322 15550
rect 33182 15538 33234 15550
rect 7634 15486 7646 15538
rect 7698 15486 7710 15538
rect 12226 15486 12238 15538
rect 12290 15486 12302 15538
rect 17490 15486 17502 15538
rect 17554 15486 17566 15538
rect 3502 15474 3554 15486
rect 8430 15474 8482 15486
rect 16270 15474 16322 15486
rect 33182 15474 33234 15486
rect 33294 15538 33346 15550
rect 33294 15474 33346 15486
rect 35310 15538 35362 15550
rect 35310 15474 35362 15486
rect 35422 15538 35474 15550
rect 35422 15474 35474 15486
rect 37326 15538 37378 15550
rect 37326 15474 37378 15486
rect 37774 15538 37826 15550
rect 37774 15474 37826 15486
rect 38222 15538 38274 15550
rect 38222 15474 38274 15486
rect 38670 15538 38722 15550
rect 38670 15474 38722 15486
rect 39790 15538 39842 15550
rect 39790 15474 39842 15486
rect 39902 15538 39954 15550
rect 39902 15474 39954 15486
rect 41134 15538 41186 15550
rect 41134 15474 41186 15486
rect 42478 15538 42530 15550
rect 42478 15474 42530 15486
rect 43486 15538 43538 15550
rect 43486 15474 43538 15486
rect 43934 15538 43986 15550
rect 43934 15474 43986 15486
rect 45054 15538 45106 15550
rect 45054 15474 45106 15486
rect 46174 15538 46226 15550
rect 46174 15474 46226 15486
rect 46958 15538 47010 15550
rect 46958 15474 47010 15486
rect 47182 15538 47234 15550
rect 47182 15474 47234 15486
rect 47742 15538 47794 15550
rect 47742 15474 47794 15486
rect 48078 15538 48130 15550
rect 48078 15474 48130 15486
rect 5854 15426 5906 15438
rect 4162 15374 4174 15426
rect 4226 15374 4238 15426
rect 4834 15374 4846 15426
rect 4898 15374 4910 15426
rect 5506 15374 5518 15426
rect 5570 15374 5582 15426
rect 5854 15362 5906 15374
rect 8318 15426 8370 15438
rect 8318 15362 8370 15374
rect 17950 15426 18002 15438
rect 17950 15362 18002 15374
rect 20526 15426 20578 15438
rect 33406 15426 33458 15438
rect 26002 15374 26014 15426
rect 26066 15374 26078 15426
rect 20526 15362 20578 15374
rect 33406 15362 33458 15374
rect 39678 15426 39730 15438
rect 39678 15362 39730 15374
rect 41246 15426 41298 15438
rect 41246 15362 41298 15374
rect 41582 15426 41634 15438
rect 47406 15426 47458 15438
rect 44258 15374 44270 15426
rect 44322 15374 44334 15426
rect 45378 15374 45390 15426
rect 45442 15374 45454 15426
rect 41582 15362 41634 15374
rect 47406 15362 47458 15374
rect 47518 15426 47570 15438
rect 47518 15362 47570 15374
rect 2606 15314 2658 15326
rect 6414 15314 6466 15326
rect 7982 15314 8034 15326
rect 3938 15262 3950 15314
rect 4002 15262 4014 15314
rect 4610 15262 4622 15314
rect 4674 15262 4686 15314
rect 5282 15262 5294 15314
rect 5346 15262 5358 15314
rect 6850 15262 6862 15314
rect 6914 15262 6926 15314
rect 2606 15250 2658 15262
rect 6414 15250 6466 15262
rect 7982 15250 8034 15262
rect 8654 15314 8706 15326
rect 8654 15250 8706 15262
rect 8766 15314 8818 15326
rect 8766 15250 8818 15262
rect 9886 15314 9938 15326
rect 12574 15314 12626 15326
rect 19070 15314 19122 15326
rect 31614 15314 31666 15326
rect 10322 15262 10334 15314
rect 10386 15262 10398 15314
rect 11442 15262 11454 15314
rect 11506 15262 11518 15314
rect 15810 15262 15822 15314
rect 15874 15262 15886 15314
rect 19394 15262 19406 15314
rect 19458 15262 19470 15314
rect 24434 15262 24446 15314
rect 24498 15262 24510 15314
rect 25218 15262 25230 15314
rect 25282 15262 25294 15314
rect 28578 15262 28590 15314
rect 28642 15262 28654 15314
rect 9886 15250 9938 15262
rect 12574 15250 12626 15262
rect 19070 15250 19122 15262
rect 31614 15250 31666 15262
rect 32062 15314 32114 15326
rect 32062 15250 32114 15262
rect 32174 15314 32226 15326
rect 34862 15314 34914 15326
rect 33954 15262 33966 15314
rect 34018 15262 34030 15314
rect 32174 15250 32226 15262
rect 34862 15250 34914 15262
rect 35198 15314 35250 15326
rect 35198 15250 35250 15262
rect 36430 15314 36482 15326
rect 36430 15250 36482 15262
rect 36878 15314 36930 15326
rect 36878 15250 36930 15262
rect 40910 15314 40962 15326
rect 40910 15250 40962 15262
rect 41806 15314 41858 15326
rect 41806 15250 41858 15262
rect 42814 15314 42866 15326
rect 42814 15250 42866 15262
rect 43150 15314 43202 15326
rect 43150 15250 43202 15262
rect 45838 15314 45890 15326
rect 45838 15250 45890 15262
rect 46846 15314 46898 15326
rect 46846 15250 46898 15262
rect 47966 15314 48018 15326
rect 47966 15250 48018 15262
rect 3166 15202 3218 15214
rect 11790 15202 11842 15214
rect 31838 15202 31890 15214
rect 35982 15202 36034 15214
rect 7186 15150 7198 15202
rect 7250 15150 7262 15202
rect 11218 15150 11230 15202
rect 11282 15150 11294 15202
rect 13010 15150 13022 15202
rect 13074 15150 13086 15202
rect 15138 15150 15150 15202
rect 15202 15150 15214 15202
rect 16706 15150 16718 15202
rect 16770 15150 16782 15202
rect 21634 15150 21646 15202
rect 21698 15150 21710 15202
rect 23762 15150 23774 15202
rect 23826 15150 23838 15202
rect 28130 15150 28142 15202
rect 28194 15150 28206 15202
rect 29250 15150 29262 15202
rect 29314 15150 29326 15202
rect 31378 15150 31390 15202
rect 31442 15150 31454 15202
rect 34066 15150 34078 15202
rect 34130 15150 34142 15202
rect 3166 15138 3218 15150
rect 11790 15138 11842 15150
rect 31838 15138 31890 15150
rect 35982 15138 36034 15150
rect 42142 15202 42194 15214
rect 42142 15138 42194 15150
rect 48078 15090 48130 15102
rect 48078 15026 48130 15038
rect 1344 14922 48608 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 48608 14922
rect 1344 14836 48608 14870
rect 13470 14754 13522 14766
rect 2370 14702 2382 14754
rect 2434 14751 2446 14754
rect 2706 14751 2718 14754
rect 2434 14705 2718 14751
rect 2434 14702 2446 14705
rect 2706 14702 2718 14705
rect 2770 14702 2782 14754
rect 13470 14690 13522 14702
rect 16494 14754 16546 14766
rect 16494 14690 16546 14702
rect 21422 14754 21474 14766
rect 21422 14690 21474 14702
rect 23662 14754 23714 14766
rect 23662 14690 23714 14702
rect 28478 14754 28530 14766
rect 28478 14690 28530 14702
rect 39790 14754 39842 14766
rect 39790 14690 39842 14702
rect 2382 14642 2434 14654
rect 2382 14578 2434 14590
rect 2830 14642 2882 14654
rect 2830 14578 2882 14590
rect 3278 14642 3330 14654
rect 3278 14578 3330 14590
rect 7870 14642 7922 14654
rect 7870 14578 7922 14590
rect 9438 14642 9490 14654
rect 9438 14578 9490 14590
rect 10446 14642 10498 14654
rect 13582 14642 13634 14654
rect 11554 14590 11566 14642
rect 11618 14590 11630 14642
rect 10446 14578 10498 14590
rect 13582 14578 13634 14590
rect 15262 14642 15314 14654
rect 26574 14642 26626 14654
rect 20738 14590 20750 14642
rect 20802 14590 20814 14642
rect 22194 14590 22206 14642
rect 22258 14590 22270 14642
rect 15262 14578 15314 14590
rect 26574 14578 26626 14590
rect 27134 14642 27186 14654
rect 27134 14578 27186 14590
rect 27582 14642 27634 14654
rect 27582 14578 27634 14590
rect 28030 14642 28082 14654
rect 28030 14578 28082 14590
rect 28590 14642 28642 14654
rect 28590 14578 28642 14590
rect 29262 14642 29314 14654
rect 34078 14642 34130 14654
rect 31490 14590 31502 14642
rect 31554 14590 31566 14642
rect 33618 14590 33630 14642
rect 33682 14590 33694 14642
rect 41346 14590 41358 14642
rect 41410 14590 41422 14642
rect 48178 14590 48190 14642
rect 48242 14590 48254 14642
rect 29262 14578 29314 14590
rect 34078 14578 34130 14590
rect 5182 14530 5234 14542
rect 5182 14466 5234 14478
rect 5518 14530 5570 14542
rect 7758 14530 7810 14542
rect 9102 14530 9154 14542
rect 7074 14478 7086 14530
rect 7138 14478 7150 14530
rect 8530 14478 8542 14530
rect 8594 14478 8606 14530
rect 5518 14466 5570 14478
rect 7758 14466 7810 14478
rect 9102 14466 9154 14478
rect 9214 14530 9266 14542
rect 9214 14466 9266 14478
rect 9662 14530 9714 14542
rect 9662 14466 9714 14478
rect 9886 14530 9938 14542
rect 9886 14466 9938 14478
rect 11118 14530 11170 14542
rect 12238 14530 12290 14542
rect 11890 14478 11902 14530
rect 11954 14478 11966 14530
rect 11118 14466 11170 14478
rect 12238 14466 12290 14478
rect 12686 14530 12738 14542
rect 15038 14530 15090 14542
rect 13794 14478 13806 14530
rect 13858 14478 13870 14530
rect 12686 14466 12738 14478
rect 15038 14466 15090 14478
rect 15710 14530 15762 14542
rect 15710 14466 15762 14478
rect 16606 14530 16658 14542
rect 16606 14466 16658 14478
rect 16942 14530 16994 14542
rect 21310 14530 21362 14542
rect 23886 14530 23938 14542
rect 17938 14478 17950 14530
rect 18002 14478 18014 14530
rect 22530 14478 22542 14530
rect 22594 14478 22606 14530
rect 16942 14466 16994 14478
rect 21310 14466 21362 14478
rect 23886 14466 23938 14478
rect 24222 14530 24274 14542
rect 25454 14530 25506 14542
rect 26462 14530 26514 14542
rect 24882 14478 24894 14530
rect 24946 14478 24958 14530
rect 26114 14478 26126 14530
rect 26178 14478 26190 14530
rect 24222 14466 24274 14478
rect 25454 14466 25506 14478
rect 26462 14466 26514 14478
rect 29038 14530 29090 14542
rect 29038 14466 29090 14478
rect 29374 14530 29426 14542
rect 29374 14466 29426 14478
rect 29710 14530 29762 14542
rect 33854 14530 33906 14542
rect 30818 14478 30830 14530
rect 30882 14478 30894 14530
rect 29710 14466 29762 14478
rect 33854 14466 33906 14478
rect 34190 14530 34242 14542
rect 34190 14466 34242 14478
rect 34526 14530 34578 14542
rect 34526 14466 34578 14478
rect 35198 14530 35250 14542
rect 35198 14466 35250 14478
rect 37326 14530 37378 14542
rect 38882 14478 38894 14530
rect 38946 14478 38958 14530
rect 44146 14478 44158 14530
rect 44210 14478 44222 14530
rect 45266 14478 45278 14530
rect 45330 14478 45342 14530
rect 37326 14466 37378 14478
rect 4846 14418 4898 14430
rect 4846 14354 4898 14366
rect 4958 14418 5010 14430
rect 4958 14354 5010 14366
rect 5966 14418 6018 14430
rect 5966 14354 6018 14366
rect 6190 14418 6242 14430
rect 6190 14354 6242 14366
rect 6638 14418 6690 14430
rect 12798 14418 12850 14430
rect 8306 14366 8318 14418
rect 8370 14366 8382 14418
rect 6638 14354 6690 14366
rect 12798 14354 12850 14366
rect 14254 14418 14306 14430
rect 14254 14354 14306 14366
rect 14478 14418 14530 14430
rect 14478 14354 14530 14366
rect 14814 14418 14866 14430
rect 14814 14354 14866 14366
rect 15486 14418 15538 14430
rect 22990 14418 23042 14430
rect 18610 14366 18622 14418
rect 18674 14366 18686 14418
rect 15486 14354 15538 14366
rect 22990 14354 23042 14366
rect 23326 14418 23378 14430
rect 23326 14354 23378 14366
rect 24110 14418 24162 14430
rect 34862 14418 34914 14430
rect 25778 14366 25790 14418
rect 25842 14366 25854 14418
rect 24110 14354 24162 14366
rect 34862 14354 34914 14366
rect 35422 14418 35474 14430
rect 35422 14354 35474 14366
rect 36318 14418 36370 14430
rect 36318 14354 36370 14366
rect 37774 14418 37826 14430
rect 37774 14354 37826 14366
rect 38222 14418 38274 14430
rect 38222 14354 38274 14366
rect 39454 14418 39506 14430
rect 39454 14354 39506 14366
rect 39678 14418 39730 14430
rect 43474 14366 43486 14418
rect 43538 14366 43550 14418
rect 46050 14366 46062 14418
rect 46114 14366 46126 14418
rect 39678 14354 39730 14366
rect 1822 14306 1874 14318
rect 1822 14242 1874 14254
rect 3614 14306 3666 14318
rect 3614 14242 3666 14254
rect 4062 14306 4114 14318
rect 4062 14242 4114 14254
rect 4622 14306 4674 14318
rect 4622 14242 4674 14254
rect 5742 14306 5794 14318
rect 5742 14242 5794 14254
rect 6526 14306 6578 14318
rect 6526 14242 6578 14254
rect 6750 14306 6802 14318
rect 6750 14242 6802 14254
rect 7534 14306 7586 14318
rect 7534 14242 7586 14254
rect 7982 14306 8034 14318
rect 12910 14306 12962 14318
rect 10770 14254 10782 14306
rect 10834 14254 10846 14306
rect 7982 14242 8034 14254
rect 12910 14242 12962 14254
rect 14590 14306 14642 14318
rect 14590 14242 14642 14254
rect 16494 14306 16546 14318
rect 21422 14306 21474 14318
rect 17266 14254 17278 14306
rect 17330 14254 17342 14306
rect 16494 14242 16546 14254
rect 21422 14242 21474 14254
rect 23550 14306 23602 14318
rect 26686 14306 26738 14318
rect 25106 14254 25118 14306
rect 25170 14254 25182 14306
rect 23550 14242 23602 14254
rect 26686 14242 26738 14254
rect 30382 14306 30434 14318
rect 30382 14242 30434 14254
rect 35310 14306 35362 14318
rect 35310 14242 35362 14254
rect 35870 14306 35922 14318
rect 39118 14306 39170 14318
rect 36978 14254 36990 14306
rect 37042 14254 37054 14306
rect 35870 14242 35922 14254
rect 39118 14242 39170 14254
rect 39342 14306 39394 14318
rect 39342 14242 39394 14254
rect 40910 14306 40962 14318
rect 40910 14242 40962 14254
rect 44942 14306 44994 14318
rect 44942 14242 44994 14254
rect 1344 14138 48608 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 48608 14138
rect 1344 14052 48608 14086
rect 2270 13970 2322 13982
rect 2270 13906 2322 13918
rect 2718 13970 2770 13982
rect 2718 13906 2770 13918
rect 6638 13970 6690 13982
rect 6638 13906 6690 13918
rect 7086 13970 7138 13982
rect 7086 13906 7138 13918
rect 7758 13970 7810 13982
rect 15262 13970 15314 13982
rect 9650 13918 9662 13970
rect 9714 13918 9726 13970
rect 7758 13906 7810 13918
rect 15262 13906 15314 13918
rect 17726 13970 17778 13982
rect 17726 13906 17778 13918
rect 23886 13970 23938 13982
rect 23886 13906 23938 13918
rect 26574 13970 26626 13982
rect 26574 13906 26626 13918
rect 28478 13970 28530 13982
rect 28478 13906 28530 13918
rect 28814 13970 28866 13982
rect 28814 13906 28866 13918
rect 29374 13970 29426 13982
rect 29374 13906 29426 13918
rect 30830 13970 30882 13982
rect 30830 13906 30882 13918
rect 31614 13970 31666 13982
rect 41022 13970 41074 13982
rect 33618 13918 33630 13970
rect 33682 13918 33694 13970
rect 31614 13906 31666 13918
rect 41022 13906 41074 13918
rect 41582 13970 41634 13982
rect 41582 13906 41634 13918
rect 43598 13970 43650 13982
rect 43598 13906 43650 13918
rect 46958 13970 47010 13982
rect 46958 13906 47010 13918
rect 47630 13970 47682 13982
rect 47630 13906 47682 13918
rect 8878 13858 8930 13870
rect 16270 13858 16322 13870
rect 4162 13806 4174 13858
rect 4226 13806 4238 13858
rect 14914 13806 14926 13858
rect 14978 13806 14990 13858
rect 15922 13806 15934 13858
rect 15986 13806 15998 13858
rect 8878 13794 8930 13806
rect 16270 13794 16322 13806
rect 16606 13858 16658 13870
rect 16606 13794 16658 13806
rect 23662 13858 23714 13870
rect 23662 13794 23714 13806
rect 24110 13858 24162 13870
rect 24110 13794 24162 13806
rect 25566 13858 25618 13870
rect 25566 13794 25618 13806
rect 45502 13858 45554 13870
rect 45502 13794 45554 13806
rect 45838 13858 45890 13870
rect 45838 13794 45890 13806
rect 46622 13858 46674 13870
rect 46622 13794 46674 13806
rect 6862 13746 6914 13758
rect 3490 13694 3502 13746
rect 3554 13694 3566 13746
rect 6862 13682 6914 13694
rect 7422 13746 7474 13758
rect 7422 13682 7474 13694
rect 7870 13746 7922 13758
rect 7870 13682 7922 13694
rect 7982 13746 8034 13758
rect 7982 13682 8034 13694
rect 8430 13746 8482 13758
rect 8430 13682 8482 13694
rect 8542 13746 8594 13758
rect 8542 13682 8594 13694
rect 8654 13746 8706 13758
rect 8654 13682 8706 13694
rect 10222 13746 10274 13758
rect 14366 13746 14418 13758
rect 16830 13746 16882 13758
rect 10658 13694 10670 13746
rect 10722 13694 10734 13746
rect 15698 13694 15710 13746
rect 15762 13694 15774 13746
rect 10222 13682 10274 13694
rect 14366 13682 14418 13694
rect 16830 13682 16882 13694
rect 17502 13746 17554 13758
rect 17502 13682 17554 13694
rect 17950 13746 18002 13758
rect 17950 13682 18002 13694
rect 18174 13746 18226 13758
rect 21422 13746 21474 13758
rect 20626 13694 20638 13746
rect 20690 13694 20702 13746
rect 18174 13682 18226 13694
rect 21422 13682 21474 13694
rect 21534 13746 21586 13758
rect 21534 13682 21586 13694
rect 21758 13746 21810 13758
rect 21758 13682 21810 13694
rect 21982 13746 22034 13758
rect 24222 13746 24274 13758
rect 23202 13694 23214 13746
rect 23266 13694 23278 13746
rect 23426 13694 23438 13746
rect 23490 13694 23502 13746
rect 21982 13682 22034 13694
rect 24222 13682 24274 13694
rect 25902 13746 25954 13758
rect 25902 13682 25954 13694
rect 26126 13746 26178 13758
rect 26126 13682 26178 13694
rect 27470 13746 27522 13758
rect 27470 13682 27522 13694
rect 30382 13746 30434 13758
rect 30382 13682 30434 13694
rect 31278 13746 31330 13758
rect 31278 13682 31330 13694
rect 33966 13746 34018 13758
rect 33966 13682 34018 13694
rect 34190 13746 34242 13758
rect 34190 13682 34242 13694
rect 34526 13746 34578 13758
rect 38446 13746 38498 13758
rect 34962 13694 34974 13746
rect 35026 13694 35038 13746
rect 34526 13682 34578 13694
rect 38446 13682 38498 13694
rect 38670 13746 38722 13758
rect 39230 13746 39282 13758
rect 38882 13694 38894 13746
rect 38946 13694 38958 13746
rect 38670 13682 38722 13694
rect 39230 13682 39282 13694
rect 39566 13746 39618 13758
rect 39566 13682 39618 13694
rect 39790 13746 39842 13758
rect 39790 13682 39842 13694
rect 40238 13746 40290 13758
rect 40238 13682 40290 13694
rect 43486 13746 43538 13758
rect 43486 13682 43538 13694
rect 43710 13746 43762 13758
rect 43710 13682 43762 13694
rect 43934 13746 43986 13758
rect 43934 13682 43986 13694
rect 46958 13746 47010 13758
rect 46958 13682 47010 13694
rect 47294 13746 47346 13758
rect 47294 13682 47346 13694
rect 47518 13746 47570 13758
rect 47518 13682 47570 13694
rect 47854 13746 47906 13758
rect 47854 13682 47906 13694
rect 3054 13634 3106 13646
rect 6750 13634 6802 13646
rect 13806 13634 13858 13646
rect 6290 13582 6302 13634
rect 6354 13582 6366 13634
rect 11330 13582 11342 13634
rect 11394 13582 11406 13634
rect 13458 13582 13470 13634
rect 13522 13582 13534 13634
rect 3054 13570 3106 13582
rect 6750 13570 6802 13582
rect 13806 13570 13858 13582
rect 16382 13634 16434 13646
rect 22318 13634 22370 13646
rect 19394 13582 19406 13634
rect 19458 13582 19470 13634
rect 16382 13570 16434 13582
rect 22318 13570 22370 13582
rect 23326 13634 23378 13646
rect 23326 13570 23378 13582
rect 24670 13634 24722 13646
rect 24670 13570 24722 13582
rect 25678 13634 25730 13646
rect 25678 13570 25730 13582
rect 27022 13634 27074 13646
rect 27022 13570 27074 13582
rect 27918 13634 27970 13646
rect 27918 13570 27970 13582
rect 29822 13634 29874 13646
rect 33070 13634 33122 13646
rect 32050 13582 32062 13634
rect 32114 13582 32126 13634
rect 29822 13570 29874 13582
rect 33070 13570 33122 13582
rect 34078 13634 34130 13646
rect 39342 13634 39394 13646
rect 35634 13582 35646 13634
rect 35698 13582 35710 13634
rect 37762 13582 37774 13634
rect 37826 13582 37838 13634
rect 34078 13570 34130 13582
rect 39342 13570 39394 13582
rect 41694 13634 41746 13646
rect 41694 13570 41746 13582
rect 9998 13522 10050 13534
rect 9998 13458 10050 13470
rect 22542 13522 22594 13534
rect 33294 13522 33346 13534
rect 22866 13470 22878 13522
rect 22930 13470 22942 13522
rect 26226 13470 26238 13522
rect 26290 13519 26302 13522
rect 27794 13519 27806 13522
rect 26290 13473 27806 13519
rect 26290 13470 26302 13473
rect 27794 13470 27806 13473
rect 27858 13470 27870 13522
rect 28018 13470 28030 13522
rect 28082 13519 28094 13522
rect 29026 13519 29038 13522
rect 28082 13473 29038 13519
rect 28082 13470 28094 13473
rect 29026 13470 29038 13473
rect 29090 13470 29102 13522
rect 22542 13458 22594 13470
rect 33294 13458 33346 13470
rect 38334 13522 38386 13534
rect 38334 13458 38386 13470
rect 41806 13522 41858 13534
rect 41806 13458 41858 13470
rect 1344 13354 48608 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 48608 13354
rect 1344 13268 48608 13302
rect 34078 13186 34130 13198
rect 2034 13134 2046 13186
rect 2098 13183 2110 13186
rect 2482 13183 2494 13186
rect 2098 13137 2494 13183
rect 2098 13134 2110 13137
rect 2482 13134 2494 13137
rect 2546 13183 2558 13186
rect 3042 13183 3054 13186
rect 2546 13137 3054 13183
rect 2546 13134 2558 13137
rect 3042 13134 3054 13137
rect 3106 13183 3118 13186
rect 4610 13183 4622 13186
rect 3106 13137 4622 13183
rect 3106 13134 3118 13137
rect 4610 13134 4622 13137
rect 4674 13134 4686 13186
rect 34078 13122 34130 13134
rect 34526 13186 34578 13198
rect 34526 13122 34578 13134
rect 2382 13074 2434 13086
rect 2382 13010 2434 13022
rect 4622 13074 4674 13086
rect 12126 13074 12178 13086
rect 28142 13074 28194 13086
rect 32622 13074 32674 13086
rect 7746 13022 7758 13074
rect 7810 13022 7822 13074
rect 9874 13022 9886 13074
rect 9938 13022 9950 13074
rect 11442 13022 11454 13074
rect 11506 13022 11518 13074
rect 16706 13022 16718 13074
rect 16770 13022 16782 13074
rect 20738 13022 20750 13074
rect 20802 13022 20814 13074
rect 27346 13022 27358 13074
rect 27410 13022 27422 13074
rect 29922 13022 29934 13074
rect 29986 13022 29998 13074
rect 32050 13022 32062 13074
rect 32114 13022 32126 13074
rect 4622 13010 4674 13022
rect 12126 13010 12178 13022
rect 28142 13010 28194 13022
rect 32622 13010 32674 13022
rect 33518 13074 33570 13086
rect 35858 13022 35870 13074
rect 35922 13022 35934 13074
rect 38546 13022 38558 13074
rect 38610 13022 38622 13074
rect 40674 13022 40686 13074
rect 40738 13022 40750 13074
rect 41010 13022 41022 13074
rect 41074 13022 41086 13074
rect 43138 13022 43150 13074
rect 43202 13022 43214 13074
rect 33518 13010 33570 13022
rect 5966 12962 6018 12974
rect 5966 12898 6018 12910
rect 6414 12962 6466 12974
rect 6414 12898 6466 12910
rect 6638 12962 6690 12974
rect 10334 12962 10386 12974
rect 7074 12910 7086 12962
rect 7138 12910 7150 12962
rect 6638 12898 6690 12910
rect 10334 12898 10386 12910
rect 10558 12962 10610 12974
rect 10558 12898 10610 12910
rect 10782 12962 10834 12974
rect 10782 12898 10834 12910
rect 11790 12962 11842 12974
rect 11790 12898 11842 12910
rect 12238 12962 12290 12974
rect 17054 12962 17106 12974
rect 13906 12910 13918 12962
rect 13970 12910 13982 12962
rect 12238 12898 12290 12910
rect 17054 12898 17106 12910
rect 17390 12962 17442 12974
rect 22430 12962 22482 12974
rect 17826 12910 17838 12962
rect 17890 12910 17902 12962
rect 18610 12910 18622 12962
rect 18674 12910 18686 12962
rect 17390 12898 17442 12910
rect 22430 12898 22482 12910
rect 22766 12962 22818 12974
rect 22766 12898 22818 12910
rect 23438 12962 23490 12974
rect 23438 12898 23490 12910
rect 23774 12962 23826 12974
rect 28030 12962 28082 12974
rect 24546 12910 24558 12962
rect 24610 12910 24622 12962
rect 25218 12910 25230 12962
rect 25282 12910 25294 12962
rect 23774 12898 23826 12910
rect 28030 12898 28082 12910
rect 28366 12962 28418 12974
rect 33742 12962 33794 12974
rect 29138 12910 29150 12962
rect 29202 12910 29214 12962
rect 33394 12910 33406 12962
rect 33458 12910 33470 12962
rect 28366 12898 28418 12910
rect 33742 12898 33794 12910
rect 34190 12962 34242 12974
rect 34190 12898 34242 12910
rect 34414 12962 34466 12974
rect 34414 12898 34466 12910
rect 35086 12962 35138 12974
rect 35086 12898 35138 12910
rect 35534 12962 35586 12974
rect 46510 12962 46562 12974
rect 36194 12910 36206 12962
rect 36258 12910 36270 12962
rect 37874 12910 37886 12962
rect 37938 12910 37950 12962
rect 43810 12910 43822 12962
rect 43874 12910 43886 12962
rect 35534 12898 35586 12910
rect 46510 12898 46562 12910
rect 46846 12962 46898 12974
rect 46846 12898 46898 12910
rect 47182 12962 47234 12974
rect 47182 12898 47234 12910
rect 12014 12850 12066 12862
rect 12014 12786 12066 12798
rect 12574 12850 12626 12862
rect 17166 12850 17218 12862
rect 14578 12798 14590 12850
rect 14642 12798 14654 12850
rect 12574 12786 12626 12798
rect 17166 12786 17218 12798
rect 21646 12850 21698 12862
rect 21646 12786 21698 12798
rect 21758 12850 21810 12862
rect 21758 12786 21810 12798
rect 21982 12850 22034 12862
rect 21982 12786 22034 12798
rect 22206 12850 22258 12862
rect 22206 12786 22258 12798
rect 23102 12850 23154 12862
rect 23102 12786 23154 12798
rect 23550 12850 23602 12862
rect 23550 12786 23602 12798
rect 28590 12850 28642 12862
rect 28590 12786 28642 12798
rect 33182 12850 33234 12862
rect 33182 12786 33234 12798
rect 34862 12850 34914 12862
rect 34862 12786 34914 12798
rect 46062 12850 46114 12862
rect 47842 12798 47854 12850
rect 47906 12798 47918 12850
rect 46062 12786 46114 12798
rect 1934 12738 1986 12750
rect 1934 12674 1986 12686
rect 2830 12738 2882 12750
rect 2830 12674 2882 12686
rect 3278 12738 3330 12750
rect 3278 12674 3330 12686
rect 3726 12738 3778 12750
rect 3726 12674 3778 12686
rect 4174 12738 4226 12750
rect 4174 12674 4226 12686
rect 5070 12738 5122 12750
rect 5070 12674 5122 12686
rect 5742 12738 5794 12750
rect 5742 12674 5794 12686
rect 6190 12738 6242 12750
rect 6190 12674 6242 12686
rect 10558 12738 10610 12750
rect 10558 12674 10610 12686
rect 11230 12738 11282 12750
rect 11230 12674 11282 12686
rect 11454 12738 11506 12750
rect 11454 12674 11506 12686
rect 22654 12738 22706 12750
rect 22654 12674 22706 12686
rect 24110 12738 24162 12750
rect 24110 12674 24162 12686
rect 35310 12738 35362 12750
rect 35310 12674 35362 12686
rect 37102 12738 37154 12750
rect 37102 12674 37154 12686
rect 44830 12738 44882 12750
rect 45726 12738 45778 12750
rect 45154 12686 45166 12738
rect 45218 12686 45230 12738
rect 44830 12674 44882 12686
rect 45726 12674 45778 12686
rect 45950 12738 46002 12750
rect 45950 12674 46002 12686
rect 46846 12738 46898 12750
rect 46846 12674 46898 12686
rect 47630 12738 47682 12750
rect 47630 12674 47682 12686
rect 48190 12738 48242 12750
rect 48190 12674 48242 12686
rect 1344 12570 48608 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 48608 12570
rect 1344 12484 48608 12518
rect 1934 12402 1986 12414
rect 1934 12338 1986 12350
rect 6750 12402 6802 12414
rect 7982 12402 8034 12414
rect 10334 12402 10386 12414
rect 7634 12350 7646 12402
rect 7698 12350 7710 12402
rect 9538 12350 9550 12402
rect 9602 12350 9614 12402
rect 6750 12338 6802 12350
rect 7982 12338 8034 12350
rect 10334 12338 10386 12350
rect 10670 12402 10722 12414
rect 10670 12338 10722 12350
rect 10894 12402 10946 12414
rect 10894 12338 10946 12350
rect 11678 12402 11730 12414
rect 11678 12338 11730 12350
rect 12126 12402 12178 12414
rect 12126 12338 12178 12350
rect 13022 12402 13074 12414
rect 13022 12338 13074 12350
rect 14030 12402 14082 12414
rect 14030 12338 14082 12350
rect 14254 12402 14306 12414
rect 14254 12338 14306 12350
rect 14590 12402 14642 12414
rect 14590 12338 14642 12350
rect 15150 12402 15202 12414
rect 15150 12338 15202 12350
rect 16270 12402 16322 12414
rect 16270 12338 16322 12350
rect 16494 12402 16546 12414
rect 16494 12338 16546 12350
rect 16718 12402 16770 12414
rect 16718 12338 16770 12350
rect 17838 12402 17890 12414
rect 17838 12338 17890 12350
rect 18510 12402 18562 12414
rect 18510 12338 18562 12350
rect 18622 12402 18674 12414
rect 18622 12338 18674 12350
rect 18734 12402 18786 12414
rect 18734 12338 18786 12350
rect 19854 12402 19906 12414
rect 19854 12338 19906 12350
rect 19966 12402 20018 12414
rect 19966 12338 20018 12350
rect 20302 12402 20354 12414
rect 20302 12338 20354 12350
rect 20414 12402 20466 12414
rect 20414 12338 20466 12350
rect 21310 12402 21362 12414
rect 21310 12338 21362 12350
rect 21534 12402 21586 12414
rect 21534 12338 21586 12350
rect 25342 12402 25394 12414
rect 25342 12338 25394 12350
rect 26350 12402 26402 12414
rect 26350 12338 26402 12350
rect 26462 12402 26514 12414
rect 26462 12338 26514 12350
rect 26574 12402 26626 12414
rect 26574 12338 26626 12350
rect 27806 12402 27858 12414
rect 27806 12338 27858 12350
rect 28478 12402 28530 12414
rect 28478 12338 28530 12350
rect 28590 12402 28642 12414
rect 28590 12338 28642 12350
rect 28702 12402 28754 12414
rect 28702 12338 28754 12350
rect 29374 12402 29426 12414
rect 29374 12338 29426 12350
rect 31614 12402 31666 12414
rect 34414 12402 34466 12414
rect 34066 12350 34078 12402
rect 34130 12350 34142 12402
rect 31614 12338 31666 12350
rect 34414 12338 34466 12350
rect 36654 12402 36706 12414
rect 36654 12338 36706 12350
rect 40350 12402 40402 12414
rect 40350 12338 40402 12350
rect 42814 12402 42866 12414
rect 42814 12338 42866 12350
rect 44158 12402 44210 12414
rect 44158 12338 44210 12350
rect 44942 12402 44994 12414
rect 44942 12338 44994 12350
rect 10110 12290 10162 12302
rect 3826 12238 3838 12290
rect 3890 12238 3902 12290
rect 8642 12238 8654 12290
rect 8706 12238 8718 12290
rect 10110 12226 10162 12238
rect 12574 12290 12626 12302
rect 12574 12226 12626 12238
rect 13918 12290 13970 12302
rect 13918 12226 13970 12238
rect 14478 12290 14530 12302
rect 14478 12226 14530 12238
rect 16382 12290 16434 12302
rect 16382 12226 16434 12238
rect 18174 12290 18226 12302
rect 18174 12226 18226 12238
rect 21198 12290 21250 12302
rect 27582 12290 27634 12302
rect 22530 12238 22542 12290
rect 22594 12238 22606 12290
rect 26002 12238 26014 12290
rect 26066 12238 26078 12290
rect 21198 12226 21250 12238
rect 27582 12226 27634 12238
rect 29822 12290 29874 12302
rect 29822 12226 29874 12238
rect 31278 12290 31330 12302
rect 31278 12226 31330 12238
rect 31390 12290 31442 12302
rect 31390 12226 31442 12238
rect 31838 12290 31890 12302
rect 31838 12226 31890 12238
rect 32062 12290 32114 12302
rect 32062 12226 32114 12238
rect 32174 12290 32226 12302
rect 41918 12290 41970 12302
rect 38994 12238 39006 12290
rect 39058 12238 39070 12290
rect 46050 12238 46062 12290
rect 46114 12238 46126 12290
rect 32174 12226 32226 12238
rect 41918 12226 41970 12238
rect 6974 12178 7026 12190
rect 8990 12178 9042 12190
rect 3042 12126 3054 12178
rect 3106 12126 3118 12178
rect 7298 12126 7310 12178
rect 7362 12126 7374 12178
rect 6974 12114 7026 12126
rect 8990 12114 9042 12126
rect 9886 12178 9938 12190
rect 9886 12114 9938 12126
rect 10446 12178 10498 12190
rect 10446 12114 10498 12126
rect 11006 12178 11058 12190
rect 11006 12114 11058 12126
rect 11566 12178 11618 12190
rect 11566 12114 11618 12126
rect 11902 12178 11954 12190
rect 11902 12114 11954 12126
rect 12350 12178 12402 12190
rect 12350 12114 12402 12126
rect 15038 12178 15090 12190
rect 15038 12114 15090 12126
rect 15374 12178 15426 12190
rect 15374 12114 15426 12126
rect 15598 12178 15650 12190
rect 15598 12114 15650 12126
rect 17614 12178 17666 12190
rect 17614 12114 17666 12126
rect 17838 12178 17890 12190
rect 17838 12114 17890 12126
rect 19182 12178 19234 12190
rect 19182 12114 19234 12126
rect 19294 12178 19346 12190
rect 19294 12114 19346 12126
rect 19742 12178 19794 12190
rect 19742 12114 19794 12126
rect 20526 12178 20578 12190
rect 20526 12114 20578 12126
rect 20974 12178 21026 12190
rect 25678 12178 25730 12190
rect 21858 12126 21870 12178
rect 21922 12126 21934 12178
rect 20974 12114 21026 12126
rect 25678 12114 25730 12126
rect 27022 12178 27074 12190
rect 27022 12114 27074 12126
rect 27918 12178 27970 12190
rect 27918 12114 27970 12126
rect 28142 12178 28194 12190
rect 29486 12178 29538 12190
rect 29026 12126 29038 12178
rect 29090 12126 29102 12178
rect 28142 12114 28194 12126
rect 29486 12114 29538 12126
rect 29598 12178 29650 12190
rect 33070 12178 33122 12190
rect 30818 12126 30830 12178
rect 30882 12126 30894 12178
rect 29598 12114 29650 12126
rect 33070 12114 33122 12126
rect 34750 12178 34802 12190
rect 34750 12114 34802 12126
rect 34862 12178 34914 12190
rect 34862 12114 34914 12126
rect 34974 12178 35026 12190
rect 34974 12114 35026 12126
rect 35422 12178 35474 12190
rect 35422 12114 35474 12126
rect 35534 12178 35586 12190
rect 36094 12178 36146 12190
rect 35858 12126 35870 12178
rect 35922 12126 35934 12178
rect 35534 12114 35586 12126
rect 36094 12114 36146 12126
rect 36318 12178 36370 12190
rect 36318 12114 36370 12126
rect 36542 12178 36594 12190
rect 39778 12126 39790 12178
rect 39842 12126 39854 12178
rect 41234 12126 41246 12178
rect 41298 12126 41310 12178
rect 45266 12126 45278 12178
rect 45330 12126 45342 12178
rect 36542 12114 36594 12126
rect 2270 12066 2322 12078
rect 2270 12002 2322 12014
rect 2830 12066 2882 12078
rect 6414 12066 6466 12078
rect 5954 12014 5966 12066
rect 6018 12014 6030 12066
rect 2830 12002 2882 12014
rect 6414 12002 6466 12014
rect 6862 12066 6914 12078
rect 30494 12066 30546 12078
rect 24658 12014 24670 12066
rect 24722 12014 24734 12066
rect 6862 12002 6914 12014
rect 30494 12002 30546 12014
rect 31502 12066 31554 12078
rect 42366 12066 42418 12078
rect 36866 12014 36878 12066
rect 36930 12014 36942 12066
rect 41122 12014 41134 12066
rect 41186 12014 41198 12066
rect 48178 12014 48190 12066
rect 48242 12014 48254 12066
rect 31502 12002 31554 12014
rect 42366 12002 42418 12014
rect 13022 11954 13074 11966
rect 13022 11890 13074 11902
rect 13134 11954 13186 11966
rect 13134 11890 13186 11902
rect 13358 11954 13410 11966
rect 13358 11890 13410 11902
rect 14590 11954 14642 11966
rect 14590 11890 14642 11902
rect 33294 11954 33346 11966
rect 33618 11902 33630 11954
rect 33682 11902 33694 11954
rect 33294 11890 33346 11902
rect 1344 11786 48608 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 48608 11786
rect 1344 11700 48608 11734
rect 7758 11618 7810 11630
rect 7758 11554 7810 11566
rect 22206 11618 22258 11630
rect 22206 11554 22258 11566
rect 23102 11618 23154 11630
rect 23102 11554 23154 11566
rect 34078 11618 34130 11630
rect 34078 11554 34130 11566
rect 34862 11618 34914 11630
rect 34862 11554 34914 11566
rect 37438 11618 37490 11630
rect 37438 11554 37490 11566
rect 46398 11618 46450 11630
rect 46398 11554 46450 11566
rect 1822 11506 1874 11518
rect 7534 11506 7586 11518
rect 5058 11454 5070 11506
rect 5122 11454 5134 11506
rect 1822 11442 1874 11454
rect 7534 11442 7586 11454
rect 12462 11506 12514 11518
rect 21310 11506 21362 11518
rect 14354 11454 14366 11506
rect 14418 11454 14430 11506
rect 16482 11454 16494 11506
rect 16546 11454 16558 11506
rect 20514 11454 20526 11506
rect 20578 11454 20590 11506
rect 12462 11442 12514 11454
rect 21310 11442 21362 11454
rect 21534 11506 21586 11518
rect 21534 11442 21586 11454
rect 22542 11506 22594 11518
rect 22542 11442 22594 11454
rect 23886 11506 23938 11518
rect 23886 11442 23938 11454
rect 24446 11506 24498 11518
rect 24446 11442 24498 11454
rect 24782 11506 24834 11518
rect 24782 11442 24834 11454
rect 25902 11506 25954 11518
rect 25902 11442 25954 11454
rect 26350 11506 26402 11518
rect 37102 11506 37154 11518
rect 31602 11454 31614 11506
rect 31666 11454 31678 11506
rect 33730 11454 33742 11506
rect 33794 11454 33806 11506
rect 35858 11454 35870 11506
rect 35922 11454 35934 11506
rect 26350 11442 26402 11454
rect 37102 11442 37154 11454
rect 37550 11506 37602 11518
rect 37550 11442 37602 11454
rect 39006 11506 39058 11518
rect 39006 11442 39058 11454
rect 40574 11506 40626 11518
rect 40574 11442 40626 11454
rect 41470 11506 41522 11518
rect 41470 11442 41522 11454
rect 43038 11506 43090 11518
rect 43038 11442 43090 11454
rect 43486 11506 43538 11518
rect 43486 11442 43538 11454
rect 5630 11394 5682 11406
rect 2258 11342 2270 11394
rect 2322 11342 2334 11394
rect 5630 11330 5682 11342
rect 6302 11394 6354 11406
rect 6302 11330 6354 11342
rect 6750 11394 6802 11406
rect 8990 11394 9042 11406
rect 10670 11394 10722 11406
rect 8082 11342 8094 11394
rect 8146 11342 8158 11394
rect 9426 11342 9438 11394
rect 9490 11342 9502 11394
rect 9650 11342 9662 11394
rect 9714 11342 9726 11394
rect 9874 11342 9886 11394
rect 9938 11342 9950 11394
rect 6750 11330 6802 11342
rect 8990 11330 9042 11342
rect 10670 11330 10722 11342
rect 11118 11394 11170 11406
rect 11118 11330 11170 11342
rect 12238 11394 12290 11406
rect 22318 11394 22370 11406
rect 26798 11394 26850 11406
rect 13570 11342 13582 11394
rect 13634 11342 13646 11394
rect 17602 11342 17614 11394
rect 17666 11342 17678 11394
rect 18386 11342 18398 11394
rect 18450 11342 18462 11394
rect 22754 11342 22766 11394
rect 22818 11342 22830 11394
rect 25330 11342 25342 11394
rect 25394 11342 25406 11394
rect 12238 11330 12290 11342
rect 22318 11330 22370 11342
rect 26798 11330 26850 11342
rect 27470 11394 27522 11406
rect 27470 11330 27522 11342
rect 29710 11394 29762 11406
rect 34526 11394 34578 11406
rect 30930 11342 30942 11394
rect 30994 11342 31006 11394
rect 29710 11330 29762 11342
rect 34526 11330 34578 11342
rect 35086 11394 35138 11406
rect 37998 11394 38050 11406
rect 35522 11342 35534 11394
rect 35586 11342 35598 11394
rect 35746 11342 35758 11394
rect 35810 11342 35822 11394
rect 35086 11330 35138 11342
rect 37998 11330 38050 11342
rect 40238 11394 40290 11406
rect 40238 11330 40290 11342
rect 41134 11394 41186 11406
rect 41134 11330 41186 11342
rect 42030 11394 42082 11406
rect 42030 11330 42082 11342
rect 42366 11394 42418 11406
rect 42366 11330 42418 11342
rect 45390 11394 45442 11406
rect 45390 11330 45442 11342
rect 45726 11394 45778 11406
rect 45726 11330 45778 11342
rect 45838 11394 45890 11406
rect 45838 11330 45890 11342
rect 46510 11394 46562 11406
rect 46510 11330 46562 11342
rect 47182 11394 47234 11406
rect 47182 11330 47234 11342
rect 47630 11394 47682 11406
rect 47630 11330 47682 11342
rect 6078 11282 6130 11294
rect 2930 11230 2942 11282
rect 2994 11230 3006 11282
rect 6078 11218 6130 11230
rect 7086 11282 7138 11294
rect 7086 11218 7138 11230
rect 8542 11282 8594 11294
rect 8542 11218 8594 11230
rect 11230 11282 11282 11294
rect 11230 11218 11282 11230
rect 11790 11282 11842 11294
rect 12686 11282 12738 11294
rect 12002 11230 12014 11282
rect 12066 11230 12078 11282
rect 11790 11218 11842 11230
rect 12686 11218 12738 11230
rect 16830 11282 16882 11294
rect 16830 11218 16882 11230
rect 17166 11282 17218 11294
rect 17166 11218 17218 11230
rect 23326 11282 23378 11294
rect 34190 11282 34242 11294
rect 25106 11230 25118 11282
rect 25170 11230 25182 11282
rect 23326 11218 23378 11230
rect 34190 11218 34242 11230
rect 44830 11282 44882 11294
rect 44830 11218 44882 11230
rect 44942 11282 44994 11294
rect 44942 11218 44994 11230
rect 46398 11282 46450 11294
rect 46398 11218 46450 11230
rect 46846 11282 46898 11294
rect 46846 11218 46898 11230
rect 47518 11282 47570 11294
rect 47518 11218 47570 11230
rect 5854 11170 5906 11182
rect 5854 11106 5906 11118
rect 6638 11170 6690 11182
rect 6638 11106 6690 11118
rect 6862 11170 6914 11182
rect 6862 11106 6914 11118
rect 8766 11170 8818 11182
rect 8766 11106 8818 11118
rect 8878 11170 8930 11182
rect 8878 11106 8930 11118
rect 11342 11170 11394 11182
rect 23214 11170 23266 11182
rect 12114 11118 12126 11170
rect 12178 11118 12190 11170
rect 21858 11118 21870 11170
rect 21922 11118 21934 11170
rect 11342 11106 11394 11118
rect 23214 11106 23266 11118
rect 26910 11170 26962 11182
rect 26910 11106 26962 11118
rect 27022 11170 27074 11182
rect 27022 11106 27074 11118
rect 27806 11170 27858 11182
rect 27806 11106 27858 11118
rect 28254 11170 28306 11182
rect 28254 11106 28306 11118
rect 29262 11170 29314 11182
rect 29262 11106 29314 11118
rect 30494 11170 30546 11182
rect 30494 11106 30546 11118
rect 34750 11170 34802 11182
rect 34750 11106 34802 11118
rect 38446 11170 38498 11182
rect 38446 11106 38498 11118
rect 42478 11170 42530 11182
rect 42478 11106 42530 11118
rect 42702 11170 42754 11182
rect 42702 11106 42754 11118
rect 45166 11170 45218 11182
rect 45166 11106 45218 11118
rect 45502 11170 45554 11182
rect 45502 11106 45554 11118
rect 46958 11170 47010 11182
rect 46958 11106 47010 11118
rect 47294 11170 47346 11182
rect 47294 11106 47346 11118
rect 1344 11002 48608 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 48608 11002
rect 1344 10916 48608 10950
rect 3054 10834 3106 10846
rect 3054 10770 3106 10782
rect 3502 10834 3554 10846
rect 3502 10770 3554 10782
rect 7198 10834 7250 10846
rect 7198 10770 7250 10782
rect 8094 10834 8146 10846
rect 8094 10770 8146 10782
rect 8654 10834 8706 10846
rect 8654 10770 8706 10782
rect 14030 10834 14082 10846
rect 14030 10770 14082 10782
rect 15038 10834 15090 10846
rect 15038 10770 15090 10782
rect 16046 10834 16098 10846
rect 16046 10770 16098 10782
rect 16270 10834 16322 10846
rect 16270 10770 16322 10782
rect 17726 10834 17778 10846
rect 17726 10770 17778 10782
rect 18174 10834 18226 10846
rect 18174 10770 18226 10782
rect 20414 10834 20466 10846
rect 20414 10770 20466 10782
rect 32398 10834 32450 10846
rect 32398 10770 32450 10782
rect 34862 10834 34914 10846
rect 34862 10770 34914 10782
rect 35534 10834 35586 10846
rect 35534 10770 35586 10782
rect 36990 10834 37042 10846
rect 36990 10770 37042 10782
rect 40014 10834 40066 10846
rect 40014 10770 40066 10782
rect 46958 10834 47010 10846
rect 46958 10770 47010 10782
rect 6974 10722 7026 10734
rect 13246 10722 13298 10734
rect 4498 10670 4510 10722
rect 4562 10670 4574 10722
rect 11890 10670 11902 10722
rect 11954 10670 11966 10722
rect 6974 10658 7026 10670
rect 13246 10658 13298 10670
rect 13358 10722 13410 10734
rect 13358 10658 13410 10670
rect 13806 10722 13858 10734
rect 14926 10722 14978 10734
rect 14242 10670 14254 10722
rect 14306 10670 14318 10722
rect 13806 10658 13858 10670
rect 14926 10658 14978 10670
rect 15486 10722 15538 10734
rect 15486 10658 15538 10670
rect 18958 10722 19010 10734
rect 20750 10722 20802 10734
rect 26126 10722 26178 10734
rect 19842 10670 19854 10722
rect 19906 10670 19918 10722
rect 23314 10670 23326 10722
rect 23378 10670 23390 10722
rect 18958 10658 19010 10670
rect 20750 10658 20802 10670
rect 26126 10658 26178 10670
rect 26462 10722 26514 10734
rect 26462 10658 26514 10670
rect 26686 10722 26738 10734
rect 30606 10722 30658 10734
rect 28018 10670 28030 10722
rect 28082 10670 28094 10722
rect 26686 10658 26738 10670
rect 30606 10658 30658 10670
rect 34190 10722 34242 10734
rect 34190 10658 34242 10670
rect 34302 10722 34354 10734
rect 34302 10658 34354 10670
rect 35310 10722 35362 10734
rect 35310 10658 35362 10670
rect 36206 10722 36258 10734
rect 36206 10658 36258 10670
rect 37550 10722 37602 10734
rect 37550 10658 37602 10670
rect 38894 10722 38946 10734
rect 46510 10722 46562 10734
rect 41010 10670 41022 10722
rect 41074 10670 41086 10722
rect 43138 10670 43150 10722
rect 43202 10670 43214 10722
rect 38894 10658 38946 10670
rect 46510 10658 46562 10670
rect 47182 10722 47234 10734
rect 47182 10658 47234 10670
rect 47294 10722 47346 10734
rect 47294 10658 47346 10670
rect 7310 10610 7362 10622
rect 3826 10558 3838 10610
rect 3890 10558 3902 10610
rect 7310 10546 7362 10558
rect 7422 10610 7474 10622
rect 13694 10610 13746 10622
rect 15262 10610 15314 10622
rect 12674 10558 12686 10610
rect 12738 10558 12750 10610
rect 14466 10558 14478 10610
rect 14530 10558 14542 10610
rect 7422 10546 7474 10558
rect 13694 10546 13746 10558
rect 15262 10546 15314 10558
rect 16382 10610 16434 10622
rect 16382 10546 16434 10558
rect 16494 10610 16546 10622
rect 16494 10546 16546 10558
rect 16942 10610 16994 10622
rect 16942 10546 16994 10558
rect 17838 10610 17890 10622
rect 17838 10546 17890 10558
rect 17950 10610 18002 10622
rect 17950 10546 18002 10558
rect 18510 10610 18562 10622
rect 18510 10546 18562 10558
rect 19182 10610 19234 10622
rect 19182 10546 19234 10558
rect 19518 10610 19570 10622
rect 19518 10546 19570 10558
rect 20974 10610 21026 10622
rect 20974 10546 21026 10558
rect 21086 10610 21138 10622
rect 21086 10546 21138 10558
rect 21198 10610 21250 10622
rect 22990 10610 23042 10622
rect 21858 10558 21870 10610
rect 21922 10558 21934 10610
rect 22082 10558 22094 10610
rect 22146 10558 22158 10610
rect 21198 10546 21250 10558
rect 22990 10546 23042 10558
rect 23774 10610 23826 10622
rect 23774 10546 23826 10558
rect 23998 10610 24050 10622
rect 30830 10610 30882 10622
rect 34526 10610 34578 10622
rect 25666 10558 25678 10610
rect 25730 10558 25742 10610
rect 27346 10558 27358 10610
rect 27410 10558 27422 10610
rect 31154 10558 31166 10610
rect 31218 10558 31230 10610
rect 23998 10546 24050 10558
rect 30830 10546 30882 10558
rect 34526 10546 34578 10558
rect 35646 10610 35698 10622
rect 35646 10546 35698 10558
rect 35870 10610 35922 10622
rect 35870 10546 35922 10558
rect 36542 10610 36594 10622
rect 36542 10546 36594 10558
rect 37998 10610 38050 10622
rect 37998 10546 38050 10558
rect 39230 10610 39282 10622
rect 39230 10546 39282 10558
rect 39678 10610 39730 10622
rect 39678 10546 39730 10558
rect 40014 10610 40066 10622
rect 40014 10546 40066 10558
rect 40350 10610 40402 10622
rect 46062 10610 46114 10622
rect 40898 10558 40910 10610
rect 40962 10558 40974 10610
rect 41794 10558 41806 10610
rect 41858 10558 41870 10610
rect 42466 10558 42478 10610
rect 42530 10558 42542 10610
rect 40350 10546 40402 10558
rect 46062 10546 46114 10558
rect 46734 10610 46786 10622
rect 46734 10546 46786 10558
rect 2158 10498 2210 10510
rect 2158 10434 2210 10446
rect 2494 10498 2546 10510
rect 9102 10498 9154 10510
rect 18734 10498 18786 10510
rect 23886 10498 23938 10510
rect 6626 10446 6638 10498
rect 6690 10446 6702 10498
rect 9762 10446 9774 10498
rect 9826 10446 9838 10498
rect 21970 10446 21982 10498
rect 22034 10446 22046 10498
rect 2494 10434 2546 10446
rect 9102 10434 9154 10446
rect 18734 10434 18786 10446
rect 23886 10434 23938 10446
rect 24446 10498 24498 10510
rect 24446 10434 24498 10446
rect 25230 10498 25282 10510
rect 25230 10434 25282 10446
rect 26238 10498 26290 10510
rect 30718 10498 30770 10510
rect 30146 10446 30158 10498
rect 30210 10446 30222 10498
rect 26238 10434 26290 10446
rect 30718 10434 30770 10446
rect 31950 10498 32002 10510
rect 31950 10434 32002 10446
rect 33182 10498 33234 10510
rect 33182 10434 33234 10446
rect 33630 10498 33682 10510
rect 46286 10498 46338 10510
rect 41010 10446 41022 10498
rect 41074 10446 41086 10498
rect 45266 10446 45278 10498
rect 45330 10446 45342 10498
rect 33630 10434 33682 10446
rect 46286 10434 46338 10446
rect 23550 10386 23602 10398
rect 21634 10334 21646 10386
rect 21698 10383 21710 10386
rect 21858 10383 21870 10386
rect 21698 10337 21870 10383
rect 21698 10334 21710 10337
rect 21858 10334 21870 10337
rect 21922 10334 21934 10386
rect 22530 10334 22542 10386
rect 22594 10334 22606 10386
rect 23550 10322 23602 10334
rect 37774 10386 37826 10398
rect 37774 10322 37826 10334
rect 38222 10386 38274 10398
rect 38222 10322 38274 10334
rect 38670 10386 38722 10398
rect 38670 10322 38722 10334
rect 1344 10218 48608 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 48608 10218
rect 1344 10132 48608 10166
rect 12798 10050 12850 10062
rect 2930 9998 2942 10050
rect 2994 10047 3006 10050
rect 3602 10047 3614 10050
rect 2994 10001 3614 10047
rect 2994 9998 3006 10001
rect 3602 9998 3614 10001
rect 3666 9998 3678 10050
rect 10210 9998 10222 10050
rect 10274 10047 10286 10050
rect 11554 10047 11566 10050
rect 10274 10001 11566 10047
rect 10274 9998 10286 10001
rect 11554 9998 11566 10001
rect 11618 9998 11630 10050
rect 12798 9986 12850 9998
rect 42814 10050 42866 10062
rect 42814 9986 42866 9998
rect 2942 9938 2994 9950
rect 2942 9874 2994 9886
rect 4622 9938 4674 9950
rect 4622 9874 4674 9886
rect 6190 9938 6242 9950
rect 6190 9874 6242 9886
rect 10110 9938 10162 9950
rect 10110 9874 10162 9886
rect 11006 9938 11058 9950
rect 11006 9874 11058 9886
rect 12014 9938 12066 9950
rect 12014 9874 12066 9886
rect 12574 9938 12626 9950
rect 12574 9874 12626 9886
rect 12910 9938 12962 9950
rect 12910 9874 12962 9886
rect 15374 9938 15426 9950
rect 19070 9938 19122 9950
rect 16370 9886 16382 9938
rect 16434 9886 16446 9938
rect 18498 9886 18510 9938
rect 18562 9886 18574 9938
rect 21634 9886 21646 9938
rect 21698 9886 21710 9938
rect 23762 9886 23774 9938
rect 23826 9886 23838 9938
rect 25666 9886 25678 9938
rect 25730 9886 25742 9938
rect 27794 9886 27806 9938
rect 27858 9886 27870 9938
rect 32050 9886 32062 9938
rect 32114 9886 32126 9938
rect 35298 9886 35310 9938
rect 35362 9886 35374 9938
rect 46050 9886 46062 9938
rect 46114 9886 46126 9938
rect 48178 9886 48190 9938
rect 48242 9886 48254 9938
rect 15374 9874 15426 9886
rect 19070 9874 19122 9886
rect 3838 9826 3890 9838
rect 3838 9762 3890 9774
rect 7870 9826 7922 9838
rect 7870 9762 7922 9774
rect 8206 9826 8258 9838
rect 8206 9762 8258 9774
rect 8542 9826 8594 9838
rect 8542 9762 8594 9774
rect 9326 9826 9378 9838
rect 9326 9762 9378 9774
rect 11678 9826 11730 9838
rect 36094 9826 36146 9838
rect 15698 9774 15710 9826
rect 15762 9774 15774 9826
rect 24546 9774 24558 9826
rect 24610 9774 24622 9826
rect 24882 9774 24894 9826
rect 24946 9774 24958 9826
rect 28242 9774 28254 9826
rect 28306 9774 28318 9826
rect 29250 9774 29262 9826
rect 29314 9774 29326 9826
rect 32498 9774 32510 9826
rect 32562 9774 32574 9826
rect 11678 9762 11730 9774
rect 36094 9762 36146 9774
rect 36990 9826 37042 9838
rect 36990 9762 37042 9774
rect 37214 9826 37266 9838
rect 37214 9762 37266 9774
rect 37998 9826 38050 9838
rect 37998 9762 38050 9774
rect 40014 9826 40066 9838
rect 42366 9826 42418 9838
rect 42130 9774 42142 9826
rect 42194 9774 42206 9826
rect 40014 9762 40066 9774
rect 42366 9762 42418 9774
rect 43038 9826 43090 9838
rect 43038 9762 43090 9774
rect 43262 9826 43314 9838
rect 44034 9774 44046 9826
rect 44098 9774 44110 9826
rect 45266 9774 45278 9826
rect 45330 9774 45342 9826
rect 43262 9762 43314 9774
rect 2046 9714 2098 9726
rect 2046 9650 2098 9662
rect 7310 9714 7362 9726
rect 7310 9650 7362 9662
rect 7534 9714 7586 9726
rect 7534 9650 7586 9662
rect 13806 9714 13858 9726
rect 13806 9650 13858 9662
rect 14814 9714 14866 9726
rect 14814 9650 14866 9662
rect 20750 9714 20802 9726
rect 37550 9714 37602 9726
rect 29922 9662 29934 9714
rect 29986 9662 29998 9714
rect 33170 9662 33182 9714
rect 33234 9662 33246 9714
rect 20750 9650 20802 9662
rect 37550 9650 37602 9662
rect 39566 9714 39618 9726
rect 39566 9650 39618 9662
rect 41022 9714 41074 9726
rect 41022 9650 41074 9662
rect 43486 9714 43538 9726
rect 44258 9662 44270 9714
rect 44322 9662 44334 9714
rect 43486 9650 43538 9662
rect 2382 9602 2434 9614
rect 2382 9538 2434 9550
rect 3390 9602 3442 9614
rect 3390 9538 3442 9550
rect 4286 9602 4338 9614
rect 4286 9538 4338 9550
rect 5070 9602 5122 9614
rect 5070 9538 5122 9550
rect 6638 9602 6690 9614
rect 6638 9538 6690 9550
rect 6974 9602 7026 9614
rect 6974 9538 7026 9550
rect 7646 9602 7698 9614
rect 7646 9538 7698 9550
rect 8318 9602 8370 9614
rect 8318 9538 8370 9550
rect 8990 9602 9042 9614
rect 8990 9538 9042 9550
rect 9214 9602 9266 9614
rect 9214 9538 9266 9550
rect 10446 9602 10498 9614
rect 10446 9538 10498 9550
rect 13918 9602 13970 9614
rect 13918 9538 13970 9550
rect 14142 9602 14194 9614
rect 14142 9538 14194 9550
rect 19406 9602 19458 9614
rect 20190 9602 20242 9614
rect 35758 9602 35810 9614
rect 37102 9602 37154 9614
rect 19842 9550 19854 9602
rect 19906 9550 19918 9602
rect 28466 9550 28478 9602
rect 28530 9550 28542 9602
rect 36418 9550 36430 9602
rect 36482 9550 36494 9602
rect 19406 9538 19458 9550
rect 20190 9538 20242 9550
rect 35758 9538 35810 9550
rect 37102 9538 37154 9550
rect 39678 9602 39730 9614
rect 39678 9538 39730 9550
rect 44942 9602 44994 9614
rect 44942 9538 44994 9550
rect 1344 9434 48608 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 48608 9434
rect 1344 9348 48608 9382
rect 2942 9266 2994 9278
rect 2942 9202 2994 9214
rect 3390 9266 3442 9278
rect 3390 9202 3442 9214
rect 7310 9266 7362 9278
rect 7310 9202 7362 9214
rect 9662 9266 9714 9278
rect 9662 9202 9714 9214
rect 10446 9266 10498 9278
rect 10446 9202 10498 9214
rect 16046 9266 16098 9278
rect 16046 9202 16098 9214
rect 17726 9266 17778 9278
rect 17726 9202 17778 9214
rect 18286 9266 18338 9278
rect 18286 9202 18338 9214
rect 23326 9266 23378 9278
rect 23326 9202 23378 9214
rect 24558 9266 24610 9278
rect 24558 9202 24610 9214
rect 25454 9266 25506 9278
rect 25454 9202 25506 9214
rect 26014 9266 26066 9278
rect 26014 9202 26066 9214
rect 26462 9266 26514 9278
rect 26462 9202 26514 9214
rect 27806 9266 27858 9278
rect 27806 9202 27858 9214
rect 28142 9266 28194 9278
rect 28142 9202 28194 9214
rect 28590 9266 28642 9278
rect 28590 9202 28642 9214
rect 29710 9266 29762 9278
rect 29710 9202 29762 9214
rect 30830 9266 30882 9278
rect 30830 9202 30882 9214
rect 32062 9266 32114 9278
rect 32062 9202 32114 9214
rect 36654 9266 36706 9278
rect 36654 9202 36706 9214
rect 37102 9266 37154 9278
rect 37102 9202 37154 9214
rect 37886 9266 37938 9278
rect 37886 9202 37938 9214
rect 38782 9266 38834 9278
rect 38782 9202 38834 9214
rect 40014 9266 40066 9278
rect 40014 9202 40066 9214
rect 44942 9266 44994 9278
rect 44942 9202 44994 9214
rect 46734 9266 46786 9278
rect 46734 9202 46786 9214
rect 47406 9266 47458 9278
rect 47406 9202 47458 9214
rect 7534 9154 7586 9166
rect 7534 9090 7586 9102
rect 8430 9154 8482 9166
rect 8430 9090 8482 9102
rect 14254 9154 14306 9166
rect 14254 9090 14306 9102
rect 15038 9154 15090 9166
rect 15038 9090 15090 9102
rect 16942 9154 16994 9166
rect 22094 9154 22146 9166
rect 17378 9102 17390 9154
rect 17442 9102 17454 9154
rect 16942 9090 16994 9102
rect 22094 9090 22146 9102
rect 23214 9154 23266 9166
rect 29150 9154 29202 9166
rect 27234 9102 27246 9154
rect 27298 9102 27310 9154
rect 23214 9090 23266 9102
rect 29150 9090 29202 9102
rect 29486 9154 29538 9166
rect 29486 9090 29538 9102
rect 29822 9154 29874 9166
rect 29822 9090 29874 9102
rect 30046 9154 30098 9166
rect 30046 9090 30098 9102
rect 30606 9154 30658 9166
rect 30606 9090 30658 9102
rect 31166 9154 31218 9166
rect 31166 9090 31218 9102
rect 31950 9154 32002 9166
rect 31950 9090 32002 9102
rect 37662 9154 37714 9166
rect 37662 9090 37714 9102
rect 38558 9154 38610 9166
rect 38558 9090 38610 9102
rect 38894 9154 38946 9166
rect 38894 9090 38946 9102
rect 39118 9154 39170 9166
rect 39118 9090 39170 9102
rect 40126 9154 40178 9166
rect 40126 9090 40178 9102
rect 40910 9154 40962 9166
rect 40910 9090 40962 9102
rect 41022 9154 41074 9166
rect 46398 9154 46450 9166
rect 45266 9102 45278 9154
rect 45330 9102 45342 9154
rect 41022 9090 41074 9102
rect 46398 9090 46450 9102
rect 47294 9154 47346 9166
rect 47294 9090 47346 9102
rect 2046 9042 2098 9054
rect 7982 9042 8034 9054
rect 8878 9042 8930 9054
rect 3714 8990 3726 9042
rect 3778 8990 3790 9042
rect 8194 8990 8206 9042
rect 8258 8990 8270 9042
rect 2046 8978 2098 8990
rect 7982 8978 8034 8990
rect 8878 8978 8930 8990
rect 9998 9042 10050 9054
rect 14030 9042 14082 9054
rect 13570 8990 13582 9042
rect 13634 8990 13646 9042
rect 9998 8978 10050 8990
rect 14030 8978 14082 8990
rect 14702 9042 14754 9054
rect 14702 8978 14754 8990
rect 14926 9042 14978 9054
rect 14926 8978 14978 8990
rect 15262 9042 15314 9054
rect 21758 9042 21810 9054
rect 18610 8990 18622 9042
rect 18674 8990 18686 9042
rect 15262 8978 15314 8990
rect 21758 8978 21810 8990
rect 22206 9042 22258 9054
rect 30830 9042 30882 9054
rect 27010 8990 27022 9042
rect 27074 8990 27086 9042
rect 22206 8978 22258 8990
rect 30830 8978 30882 8990
rect 31390 9042 31442 9054
rect 31390 8978 31442 8990
rect 31838 9042 31890 9054
rect 37886 9042 37938 9054
rect 36082 8990 36094 9042
rect 36146 8990 36158 9042
rect 31838 8978 31890 8990
rect 37886 8978 37938 8990
rect 38222 9042 38274 9054
rect 38222 8978 38274 8990
rect 39678 9042 39730 9054
rect 39678 8978 39730 8990
rect 40350 9042 40402 9054
rect 40350 8978 40402 8990
rect 41246 9042 41298 9054
rect 46622 9042 46674 9054
rect 44482 8990 44494 9042
rect 44546 8990 44558 9042
rect 41246 8978 41298 8990
rect 46622 8978 46674 8990
rect 47070 9042 47122 9054
rect 47070 8978 47122 8990
rect 47854 9042 47906 9054
rect 47854 8978 47906 8990
rect 2494 8930 2546 8942
rect 7422 8930 7474 8942
rect 14478 8930 14530 8942
rect 4386 8878 4398 8930
rect 4450 8878 4462 8930
rect 6514 8878 6526 8930
rect 6578 8878 6590 8930
rect 7858 8878 7870 8930
rect 7922 8878 7934 8930
rect 10770 8878 10782 8930
rect 10834 8878 10846 8930
rect 12898 8878 12910 8930
rect 12962 8878 12974 8930
rect 2494 8866 2546 8878
rect 7422 8866 7474 8878
rect 14478 8866 14530 8878
rect 16494 8930 16546 8942
rect 21870 8930 21922 8942
rect 19282 8878 19294 8930
rect 19346 8878 19358 8930
rect 21410 8878 21422 8930
rect 21474 8878 21486 8930
rect 16494 8866 16546 8878
rect 21870 8866 21922 8878
rect 22766 8930 22818 8942
rect 22766 8866 22818 8878
rect 23886 8930 23938 8942
rect 23886 8866 23938 8878
rect 32510 8930 32562 8942
rect 45726 8930 45778 8942
rect 33282 8878 33294 8930
rect 33346 8878 33358 8930
rect 35410 8878 35422 8930
rect 35474 8878 35486 8930
rect 41682 8878 41694 8930
rect 41746 8878 41758 8930
rect 43810 8878 43822 8930
rect 43874 8878 43886 8930
rect 32510 8866 32562 8878
rect 45726 8866 45778 8878
rect 47966 8930 48018 8942
rect 47966 8866 48018 8878
rect 8766 8818 8818 8830
rect 47406 8818 47458 8830
rect 2482 8766 2494 8818
rect 2546 8815 2558 8818
rect 2706 8815 2718 8818
rect 2546 8769 2718 8815
rect 2546 8766 2558 8769
rect 2706 8766 2718 8769
rect 2770 8815 2782 8818
rect 3266 8815 3278 8818
rect 2770 8769 3278 8815
rect 2770 8766 2782 8769
rect 3266 8766 3278 8769
rect 3330 8766 3342 8818
rect 15810 8766 15822 8818
rect 15874 8815 15886 8818
rect 16482 8815 16494 8818
rect 15874 8769 16494 8815
rect 15874 8766 15886 8769
rect 16482 8766 16494 8769
rect 16546 8766 16558 8818
rect 23874 8766 23886 8818
rect 23938 8815 23950 8818
rect 24658 8815 24670 8818
rect 23938 8769 24670 8815
rect 23938 8766 23950 8769
rect 24658 8766 24670 8769
rect 24722 8766 24734 8818
rect 27906 8766 27918 8818
rect 27970 8815 27982 8818
rect 28466 8815 28478 8818
rect 27970 8769 28478 8815
rect 27970 8766 27982 8769
rect 28466 8766 28478 8769
rect 28530 8766 28542 8818
rect 8766 8754 8818 8766
rect 47406 8754 47458 8766
rect 1344 8650 48608 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 48608 8650
rect 1344 8564 48608 8598
rect 4846 8482 4898 8494
rect 4846 8418 4898 8430
rect 7422 8482 7474 8494
rect 7422 8418 7474 8430
rect 8878 8482 8930 8494
rect 8878 8418 8930 8430
rect 36318 8482 36370 8494
rect 36318 8418 36370 8430
rect 1934 8370 1986 8382
rect 1934 8306 1986 8318
rect 3278 8370 3330 8382
rect 3278 8306 3330 8318
rect 4174 8370 4226 8382
rect 4174 8306 4226 8318
rect 4958 8370 5010 8382
rect 8654 8370 8706 8382
rect 19182 8370 19234 8382
rect 6402 8367 6414 8370
rect 4958 8306 5010 8318
rect 6193 8321 6414 8367
rect 3726 8258 3778 8270
rect 3726 8194 3778 8206
rect 2382 8146 2434 8158
rect 2382 8082 2434 8094
rect 5742 8146 5794 8158
rect 5842 8094 5854 8146
rect 5906 8143 5918 8146
rect 6193 8143 6239 8321
rect 6402 8318 6414 8321
rect 6466 8318 6478 8370
rect 12786 8318 12798 8370
rect 12850 8318 12862 8370
rect 13458 8318 13470 8370
rect 13522 8318 13534 8370
rect 8654 8306 8706 8318
rect 19182 8306 19234 8318
rect 22654 8370 22706 8382
rect 22654 8306 22706 8318
rect 28590 8370 28642 8382
rect 28590 8306 28642 8318
rect 32062 8370 32114 8382
rect 37102 8370 37154 8382
rect 32498 8318 32510 8370
rect 32562 8318 32574 8370
rect 46050 8318 46062 8370
rect 46114 8318 46126 8370
rect 48178 8318 48190 8370
rect 48242 8318 48254 8370
rect 32062 8306 32114 8318
rect 37102 8306 37154 8318
rect 6862 8258 6914 8270
rect 6402 8206 6414 8258
rect 6466 8206 6478 8258
rect 6862 8194 6914 8206
rect 7310 8258 7362 8270
rect 8206 8258 8258 8270
rect 7970 8206 7982 8258
rect 8034 8206 8046 8258
rect 7310 8194 7362 8206
rect 8206 8194 8258 8206
rect 9102 8258 9154 8270
rect 9102 8194 9154 8206
rect 9326 8258 9378 8270
rect 18174 8258 18226 8270
rect 10658 8206 10670 8258
rect 10722 8206 10734 8258
rect 12002 8206 12014 8258
rect 12066 8206 12078 8258
rect 12338 8206 12350 8258
rect 12402 8206 12414 8258
rect 16258 8206 16270 8258
rect 16322 8206 16334 8258
rect 17490 8206 17502 8258
rect 17554 8206 17566 8258
rect 9326 8194 9378 8206
rect 18174 8194 18226 8206
rect 19518 8258 19570 8270
rect 19518 8194 19570 8206
rect 19854 8258 19906 8270
rect 21534 8258 21586 8270
rect 27806 8258 27858 8270
rect 20178 8206 20190 8258
rect 20242 8206 20254 8258
rect 23650 8206 23662 8258
rect 23714 8206 23726 8258
rect 25890 8206 25902 8258
rect 25954 8206 25966 8258
rect 19854 8194 19906 8206
rect 21534 8194 21586 8206
rect 27806 8194 27858 8206
rect 33854 8258 33906 8270
rect 33854 8194 33906 8206
rect 34526 8258 34578 8270
rect 34526 8194 34578 8206
rect 34750 8258 34802 8270
rect 34750 8194 34802 8206
rect 35870 8258 35922 8270
rect 35870 8194 35922 8206
rect 36206 8258 36258 8270
rect 36206 8194 36258 8206
rect 37774 8258 37826 8270
rect 37774 8194 37826 8206
rect 37998 8258 38050 8270
rect 37998 8194 38050 8206
rect 38894 8258 38946 8270
rect 38894 8194 38946 8206
rect 39566 8258 39618 8270
rect 39566 8194 39618 8206
rect 39790 8258 39842 8270
rect 39790 8194 39842 8206
rect 40910 8258 40962 8270
rect 40910 8194 40962 8206
rect 41022 8258 41074 8270
rect 42142 8258 42194 8270
rect 41906 8206 41918 8258
rect 41970 8206 41982 8258
rect 41022 8194 41074 8206
rect 42142 8194 42194 8206
rect 42590 8258 42642 8270
rect 42590 8194 42642 8206
rect 42814 8258 42866 8270
rect 42814 8194 42866 8206
rect 43822 8258 43874 8270
rect 43822 8194 43874 8206
rect 44158 8258 44210 8270
rect 45378 8206 45390 8258
rect 45442 8206 45454 8258
rect 44158 8194 44210 8206
rect 5906 8097 6239 8143
rect 8094 8146 8146 8158
rect 16830 8146 16882 8158
rect 5906 8094 5918 8097
rect 10434 8094 10446 8146
rect 10498 8094 10510 8146
rect 12786 8094 12798 8146
rect 12850 8094 12862 8146
rect 15586 8094 15598 8146
rect 15650 8094 15662 8146
rect 5742 8082 5794 8094
rect 8094 8082 8146 8094
rect 16830 8082 16882 8094
rect 17054 8146 17106 8158
rect 17054 8082 17106 8094
rect 18510 8146 18562 8158
rect 18510 8082 18562 8094
rect 18846 8146 18898 8158
rect 18846 8082 18898 8094
rect 19070 8146 19122 8158
rect 19070 8082 19122 8094
rect 20414 8146 20466 8158
rect 20414 8082 20466 8094
rect 21422 8146 21474 8158
rect 26350 8146 26402 8158
rect 23762 8094 23774 8146
rect 23826 8094 23838 8146
rect 21422 8082 21474 8094
rect 26350 8082 26402 8094
rect 29486 8146 29538 8158
rect 30382 8146 30434 8158
rect 29586 8094 29598 8146
rect 29650 8094 29662 8146
rect 29486 8082 29538 8094
rect 30382 8082 30434 8094
rect 31278 8146 31330 8158
rect 31278 8082 31330 8094
rect 34190 8146 34242 8158
rect 34190 8082 34242 8094
rect 35086 8146 35138 8158
rect 35086 8082 35138 8094
rect 35422 8146 35474 8158
rect 35422 8082 35474 8094
rect 35758 8146 35810 8158
rect 35758 8082 35810 8094
rect 41358 8146 41410 8158
rect 43150 8146 43202 8158
rect 41570 8094 41582 8146
rect 41634 8094 41646 8146
rect 41358 8082 41410 8094
rect 43150 8082 43202 8094
rect 2830 8034 2882 8046
rect 2830 7970 2882 7982
rect 4622 8034 4674 8046
rect 4622 7970 4674 7982
rect 5630 8034 5682 8046
rect 5630 7970 5682 7982
rect 6750 8034 6802 8046
rect 6750 7970 6802 7982
rect 6974 8034 7026 8046
rect 6974 7970 7026 7982
rect 7758 8034 7810 8046
rect 7758 7970 7810 7982
rect 9774 8034 9826 8046
rect 9774 7970 9826 7982
rect 10222 8034 10274 8046
rect 11454 8034 11506 8046
rect 11106 7982 11118 8034
rect 11170 7982 11182 8034
rect 10222 7970 10274 7982
rect 11454 7970 11506 7982
rect 16718 8034 16770 8046
rect 16718 7970 16770 7982
rect 16942 8034 16994 8046
rect 18622 8034 18674 8046
rect 17826 7982 17838 8034
rect 17890 7982 17902 8034
rect 16942 7970 16994 7982
rect 18622 7970 18674 7982
rect 19630 8034 19682 8046
rect 19630 7970 19682 7982
rect 21198 8034 21250 8046
rect 21198 7970 21250 7982
rect 21982 8034 22034 8046
rect 23326 8034 23378 8046
rect 29150 8034 29202 8046
rect 22978 7982 22990 8034
rect 23042 7982 23054 8034
rect 26450 7982 26462 8034
rect 26514 7982 26526 8034
rect 28130 7982 28142 8034
rect 28194 7982 28206 8034
rect 21982 7970 22034 7982
rect 23326 7970 23378 7982
rect 29150 7970 29202 7982
rect 29262 8034 29314 8046
rect 29262 7970 29314 7982
rect 29374 8034 29426 8046
rect 29374 7970 29426 7982
rect 30270 8034 30322 8046
rect 30270 7970 30322 7982
rect 30830 8034 30882 8046
rect 30830 7970 30882 7982
rect 32958 8034 33010 8046
rect 32958 7970 33010 7982
rect 33294 8034 33346 8046
rect 33294 7970 33346 7982
rect 34414 8034 34466 8046
rect 34414 7970 34466 7982
rect 35198 8034 35250 8046
rect 35198 7970 35250 7982
rect 35534 8034 35586 8046
rect 35534 7970 35586 7982
rect 36318 8034 36370 8046
rect 38446 8034 38498 8046
rect 37426 7982 37438 8034
rect 37490 7982 37502 8034
rect 36318 7970 36370 7982
rect 38446 7970 38498 7982
rect 38670 8034 38722 8046
rect 38670 7970 38722 7982
rect 38782 8034 38834 8046
rect 40238 8034 40290 8046
rect 39218 7982 39230 8034
rect 39282 7982 39294 8034
rect 38782 7970 38834 7982
rect 40238 7970 40290 7982
rect 41694 8034 41746 8046
rect 41694 7970 41746 7982
rect 42478 8034 42530 8046
rect 42478 7970 42530 7982
rect 43262 8034 43314 8046
rect 43262 7970 43314 7982
rect 43374 8034 43426 8046
rect 43374 7970 43426 7982
rect 44942 8034 44994 8046
rect 44942 7970 44994 7982
rect 1344 7866 48608 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 48608 7866
rect 1344 7780 48608 7814
rect 1822 7698 1874 7710
rect 1822 7634 1874 7646
rect 6974 7698 7026 7710
rect 8654 7698 8706 7710
rect 8082 7646 8094 7698
rect 8146 7646 8158 7698
rect 6974 7634 7026 7646
rect 8654 7634 8706 7646
rect 9102 7698 9154 7710
rect 10334 7698 10386 7710
rect 15150 7698 15202 7710
rect 9986 7646 9998 7698
rect 10050 7646 10062 7698
rect 10882 7646 10894 7698
rect 10946 7646 10958 7698
rect 9102 7634 9154 7646
rect 10334 7634 10386 7646
rect 15150 7634 15202 7646
rect 15934 7698 15986 7710
rect 15934 7634 15986 7646
rect 16382 7698 16434 7710
rect 16382 7634 16434 7646
rect 16942 7698 16994 7710
rect 16942 7634 16994 7646
rect 18846 7698 18898 7710
rect 18846 7634 18898 7646
rect 19294 7698 19346 7710
rect 19294 7634 19346 7646
rect 19854 7698 19906 7710
rect 19854 7634 19906 7646
rect 23102 7698 23154 7710
rect 23102 7634 23154 7646
rect 23438 7698 23490 7710
rect 23438 7634 23490 7646
rect 23886 7698 23938 7710
rect 23886 7634 23938 7646
rect 27582 7698 27634 7710
rect 27582 7634 27634 7646
rect 27806 7698 27858 7710
rect 33742 7698 33794 7710
rect 38894 7698 38946 7710
rect 32274 7646 32286 7698
rect 32338 7646 32350 7698
rect 35858 7646 35870 7698
rect 35922 7646 35934 7698
rect 27806 7634 27858 7646
rect 33742 7634 33794 7646
rect 38894 7634 38946 7646
rect 40126 7698 40178 7710
rect 40126 7634 40178 7646
rect 40238 7698 40290 7710
rect 40238 7634 40290 7646
rect 40350 7698 40402 7710
rect 40350 7634 40402 7646
rect 41470 7698 41522 7710
rect 43822 7698 43874 7710
rect 42802 7646 42814 7698
rect 42866 7646 42878 7698
rect 41470 7634 41522 7646
rect 43822 7634 43874 7646
rect 44270 7698 44322 7710
rect 44270 7634 44322 7646
rect 45054 7698 45106 7710
rect 45054 7634 45106 7646
rect 45614 7698 45666 7710
rect 45614 7634 45666 7646
rect 46622 7698 46674 7710
rect 46622 7634 46674 7646
rect 46846 7698 46898 7710
rect 46846 7634 46898 7646
rect 47406 7698 47458 7710
rect 47406 7634 47458 7646
rect 47854 7698 47906 7710
rect 47854 7634 47906 7646
rect 6638 7586 6690 7598
rect 13806 7586 13858 7598
rect 15822 7586 15874 7598
rect 4162 7534 4174 7586
rect 4226 7534 4238 7586
rect 10770 7534 10782 7586
rect 10834 7534 10846 7586
rect 14802 7534 14814 7586
rect 14866 7534 14878 7586
rect 6638 7522 6690 7534
rect 13806 7522 13858 7534
rect 15822 7522 15874 7534
rect 20638 7586 20690 7598
rect 20638 7522 20690 7534
rect 21086 7586 21138 7598
rect 21086 7522 21138 7534
rect 21982 7586 22034 7598
rect 25790 7586 25842 7598
rect 24210 7534 24222 7586
rect 24274 7534 24286 7586
rect 21982 7522 22034 7534
rect 25790 7522 25842 7534
rect 26574 7586 26626 7598
rect 26574 7522 26626 7534
rect 27470 7586 27522 7598
rect 33070 7586 33122 7598
rect 34750 7586 34802 7598
rect 28802 7534 28814 7586
rect 28866 7534 28878 7586
rect 31378 7534 31390 7586
rect 31442 7534 31454 7586
rect 33394 7534 33406 7586
rect 33458 7534 33470 7586
rect 27470 7522 27522 7534
rect 33070 7522 33122 7534
rect 34750 7522 34802 7534
rect 35198 7586 35250 7598
rect 35198 7522 35250 7534
rect 36766 7586 36818 7598
rect 36766 7522 36818 7534
rect 37214 7586 37266 7598
rect 37214 7522 37266 7534
rect 39118 7586 39170 7598
rect 48190 7586 48242 7598
rect 41234 7534 41246 7586
rect 41298 7534 41310 7586
rect 44594 7534 44606 7586
rect 44658 7534 44670 7586
rect 39118 7522 39170 7534
rect 48190 7522 48242 7534
rect 6974 7474 7026 7486
rect 3490 7422 3502 7474
rect 3554 7422 3566 7474
rect 6974 7410 7026 7422
rect 7310 7474 7362 7486
rect 7310 7410 7362 7422
rect 7534 7474 7586 7486
rect 7534 7410 7586 7422
rect 7758 7474 7810 7486
rect 14366 7474 14418 7486
rect 12226 7422 12238 7474
rect 12290 7422 12302 7474
rect 7758 7410 7810 7422
rect 14366 7410 14418 7422
rect 17278 7474 17330 7486
rect 17278 7410 17330 7422
rect 17726 7474 17778 7486
rect 17726 7410 17778 7422
rect 17838 7474 17890 7486
rect 17838 7410 17890 7422
rect 19630 7474 19682 7486
rect 19630 7410 19682 7422
rect 20302 7474 20354 7486
rect 21198 7474 21250 7486
rect 20962 7422 20974 7474
rect 21026 7422 21038 7474
rect 20302 7410 20354 7422
rect 21198 7410 21250 7422
rect 22206 7474 22258 7486
rect 22206 7410 22258 7422
rect 24558 7474 24610 7486
rect 26910 7474 26962 7486
rect 25554 7422 25566 7474
rect 25618 7422 25630 7474
rect 24558 7410 24610 7422
rect 26910 7410 26962 7422
rect 27134 7474 27186 7486
rect 36206 7474 36258 7486
rect 28018 7422 28030 7474
rect 28082 7422 28094 7474
rect 31266 7422 31278 7474
rect 31330 7422 31342 7474
rect 32162 7422 32174 7474
rect 32226 7422 32238 7474
rect 35522 7422 35534 7474
rect 35586 7422 35598 7474
rect 27134 7410 27186 7422
rect 36206 7410 36258 7422
rect 36990 7474 37042 7486
rect 36990 7410 37042 7422
rect 38110 7474 38162 7486
rect 38110 7410 38162 7422
rect 38670 7474 38722 7486
rect 38670 7410 38722 7422
rect 39678 7474 39730 7486
rect 41134 7474 41186 7486
rect 40898 7422 40910 7474
rect 40962 7422 40974 7474
rect 39678 7410 39730 7422
rect 41134 7410 41186 7422
rect 41806 7474 41858 7486
rect 41806 7410 41858 7422
rect 41918 7474 41970 7486
rect 41918 7410 41970 7422
rect 42254 7474 42306 7486
rect 42254 7410 42306 7422
rect 42478 7474 42530 7486
rect 42478 7410 42530 7422
rect 43710 7474 43762 7486
rect 43710 7410 43762 7422
rect 44046 7474 44098 7486
rect 44046 7410 44098 7422
rect 45166 7474 45218 7486
rect 45166 7410 45218 7422
rect 46958 7474 47010 7486
rect 46958 7410 47010 7422
rect 47294 7474 47346 7486
rect 47294 7410 47346 7422
rect 2718 7362 2770 7374
rect 2718 7298 2770 7310
rect 3166 7362 3218 7374
rect 9774 7362 9826 7374
rect 6290 7310 6302 7362
rect 6354 7310 6366 7362
rect 3166 7298 3218 7310
rect 9774 7298 9826 7310
rect 17502 7362 17554 7374
rect 17502 7298 17554 7310
rect 18510 7362 18562 7374
rect 18510 7298 18562 7310
rect 26350 7362 26402 7374
rect 26350 7298 26402 7310
rect 26686 7362 26738 7374
rect 34302 7362 34354 7374
rect 30930 7310 30942 7362
rect 30994 7310 31006 7362
rect 26686 7298 26738 7310
rect 34302 7298 34354 7310
rect 36430 7362 36482 7374
rect 36430 7298 36482 7310
rect 36878 7362 36930 7374
rect 36878 7298 36930 7310
rect 38334 7362 38386 7374
rect 38334 7298 38386 7310
rect 38782 7362 38834 7374
rect 38782 7298 38834 7310
rect 43262 7362 43314 7374
rect 43262 7298 43314 7310
rect 19966 7250 20018 7262
rect 16146 7198 16158 7250
rect 16210 7247 16222 7250
rect 16706 7247 16718 7250
rect 16210 7201 16718 7247
rect 16210 7198 16222 7201
rect 16706 7198 16718 7201
rect 16770 7198 16782 7250
rect 19966 7186 20018 7198
rect 20414 7250 20466 7262
rect 20414 7186 20466 7198
rect 22430 7250 22482 7262
rect 22430 7186 22482 7198
rect 22654 7250 22706 7262
rect 22654 7186 22706 7198
rect 35534 7250 35586 7262
rect 45054 7250 45106 7262
rect 37762 7198 37774 7250
rect 37826 7198 37838 7250
rect 35534 7186 35586 7198
rect 45054 7186 45106 7198
rect 47406 7250 47458 7262
rect 47406 7186 47458 7198
rect 1344 7082 48608 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 48608 7082
rect 1344 6996 48608 7030
rect 11454 6914 11506 6926
rect 2818 6862 2830 6914
rect 2882 6911 2894 6914
rect 3490 6911 3502 6914
rect 2882 6865 3502 6911
rect 2882 6862 2894 6865
rect 3490 6862 3502 6865
rect 3554 6911 3566 6914
rect 4610 6911 4622 6914
rect 3554 6865 4622 6911
rect 3554 6862 3566 6865
rect 4610 6862 4622 6865
rect 4674 6862 4686 6914
rect 11454 6850 11506 6862
rect 11678 6914 11730 6926
rect 11678 6850 11730 6862
rect 35310 6914 35362 6926
rect 35310 6850 35362 6862
rect 38110 6914 38162 6926
rect 38110 6850 38162 6862
rect 38222 6914 38274 6926
rect 38222 6850 38274 6862
rect 39454 6914 39506 6926
rect 39454 6850 39506 6862
rect 39566 6914 39618 6926
rect 39566 6850 39618 6862
rect 2830 6802 2882 6814
rect 2830 6738 2882 6750
rect 4622 6802 4674 6814
rect 4622 6738 4674 6750
rect 8430 6802 8482 6814
rect 8430 6738 8482 6750
rect 13022 6802 13074 6814
rect 17838 6802 17890 6814
rect 27470 6802 27522 6814
rect 14130 6750 14142 6802
rect 14194 6750 14206 6802
rect 27010 6750 27022 6802
rect 27074 6750 27086 6802
rect 13022 6738 13074 6750
rect 17838 6738 17890 6750
rect 27470 6738 27522 6750
rect 28366 6802 28418 6814
rect 28366 6738 28418 6750
rect 32398 6802 32450 6814
rect 32398 6738 32450 6750
rect 34862 6802 34914 6814
rect 48302 6802 48354 6814
rect 39106 6750 39118 6802
rect 39170 6750 39182 6802
rect 44258 6750 44270 6802
rect 44322 6750 44334 6802
rect 34862 6738 34914 6750
rect 48302 6738 48354 6750
rect 3838 6690 3890 6702
rect 6750 6690 6802 6702
rect 5842 6638 5854 6690
rect 5906 6638 5918 6690
rect 3838 6626 3890 6638
rect 6750 6626 6802 6638
rect 6974 6690 7026 6702
rect 6974 6626 7026 6638
rect 7422 6690 7474 6702
rect 7422 6626 7474 6638
rect 8990 6690 9042 6702
rect 8990 6626 9042 6638
rect 9214 6690 9266 6702
rect 9214 6626 9266 6638
rect 9550 6690 9602 6702
rect 9550 6626 9602 6638
rect 9662 6690 9714 6702
rect 9662 6626 9714 6638
rect 10446 6690 10498 6702
rect 10446 6626 10498 6638
rect 10670 6690 10722 6702
rect 10670 6626 10722 6638
rect 11230 6690 11282 6702
rect 11230 6626 11282 6638
rect 12126 6690 12178 6702
rect 17950 6690 18002 6702
rect 13682 6638 13694 6690
rect 13746 6638 13758 6690
rect 16258 6638 16270 6690
rect 16322 6638 16334 6690
rect 17042 6638 17054 6690
rect 17106 6638 17118 6690
rect 12126 6626 12178 6638
rect 17950 6626 18002 6638
rect 18174 6690 18226 6702
rect 18174 6626 18226 6638
rect 19518 6690 19570 6702
rect 19518 6626 19570 6638
rect 19854 6690 19906 6702
rect 19854 6626 19906 6638
rect 20078 6690 20130 6702
rect 20078 6626 20130 6638
rect 21534 6690 21586 6702
rect 21534 6626 21586 6638
rect 21870 6690 21922 6702
rect 21870 6626 21922 6638
rect 22094 6690 22146 6702
rect 27358 6690 27410 6702
rect 23538 6638 23550 6690
rect 23602 6638 23614 6690
rect 24210 6638 24222 6690
rect 24274 6638 24286 6690
rect 24882 6638 24894 6690
rect 24946 6638 24958 6690
rect 22094 6626 22146 6638
rect 27358 6626 27410 6638
rect 29934 6690 29986 6702
rect 29934 6626 29986 6638
rect 30270 6690 30322 6702
rect 30270 6626 30322 6638
rect 31278 6690 31330 6702
rect 31278 6626 31330 6638
rect 31502 6690 31554 6702
rect 31502 6626 31554 6638
rect 32174 6690 32226 6702
rect 33070 6690 33122 6702
rect 32722 6638 32734 6690
rect 32786 6638 32798 6690
rect 32174 6626 32226 6638
rect 33070 6626 33122 6638
rect 33294 6690 33346 6702
rect 35422 6690 35474 6702
rect 37102 6690 37154 6702
rect 40350 6690 40402 6702
rect 44718 6690 44770 6702
rect 33618 6638 33630 6690
rect 33682 6638 33694 6690
rect 34290 6638 34302 6690
rect 34354 6638 34366 6690
rect 36306 6638 36318 6690
rect 36370 6638 36382 6690
rect 38770 6638 38782 6690
rect 38834 6638 38846 6690
rect 40114 6638 40126 6690
rect 40178 6638 40190 6690
rect 41346 6638 41358 6690
rect 41410 6638 41422 6690
rect 33294 6626 33346 6638
rect 35422 6626 35474 6638
rect 37102 6626 37154 6638
rect 40350 6626 40402 6638
rect 44718 6626 44770 6638
rect 45054 6690 45106 6702
rect 45054 6626 45106 6638
rect 46958 6690 47010 6702
rect 46958 6626 47010 6638
rect 47294 6690 47346 6702
rect 47294 6626 47346 6638
rect 47854 6690 47906 6702
rect 47854 6626 47906 6638
rect 3390 6578 3442 6590
rect 3390 6514 3442 6526
rect 4286 6578 4338 6590
rect 4286 6514 4338 6526
rect 11006 6578 11058 6590
rect 11006 6514 11058 6526
rect 12574 6578 12626 6590
rect 12574 6514 12626 6526
rect 17502 6578 17554 6590
rect 17502 6514 17554 6526
rect 18622 6578 18674 6590
rect 18622 6514 18674 6526
rect 18846 6578 18898 6590
rect 18846 6514 18898 6526
rect 22430 6578 22482 6590
rect 22430 6514 22482 6526
rect 27582 6578 27634 6590
rect 27582 6514 27634 6526
rect 27806 6578 27858 6590
rect 27806 6514 27858 6526
rect 30606 6578 30658 6590
rect 30606 6514 30658 6526
rect 30830 6578 30882 6590
rect 30830 6514 30882 6526
rect 35758 6578 35810 6590
rect 38558 6578 38610 6590
rect 35970 6526 35982 6578
rect 36034 6526 36046 6578
rect 37762 6526 37774 6578
rect 37826 6526 37838 6578
rect 35758 6514 35810 6526
rect 38558 6514 38610 6526
rect 39006 6578 39058 6590
rect 39006 6514 39058 6526
rect 39790 6578 39842 6590
rect 44942 6578 44994 6590
rect 42130 6526 42142 6578
rect 42194 6526 42206 6578
rect 39790 6514 39842 6526
rect 44942 6514 44994 6526
rect 45390 6578 45442 6590
rect 45390 6514 45442 6526
rect 46062 6578 46114 6590
rect 46062 6514 46114 6526
rect 46622 6578 46674 6590
rect 46622 6514 46674 6526
rect 47518 6578 47570 6590
rect 47518 6514 47570 6526
rect 5182 6466 5234 6478
rect 5182 6402 5234 6414
rect 6190 6466 6242 6478
rect 6190 6402 6242 6414
rect 6302 6466 6354 6478
rect 6302 6402 6354 6414
rect 6414 6466 6466 6478
rect 6414 6402 6466 6414
rect 7086 6466 7138 6478
rect 7086 6402 7138 6414
rect 8094 6466 8146 6478
rect 8094 6402 8146 6414
rect 8318 6466 8370 6478
rect 8318 6402 8370 6414
rect 8542 6466 8594 6478
rect 8542 6402 8594 6414
rect 9326 6466 9378 6478
rect 17726 6466 17778 6478
rect 10098 6414 10110 6466
rect 10162 6414 10174 6466
rect 13458 6414 13470 6466
rect 13522 6414 13534 6466
rect 9326 6402 9378 6414
rect 17726 6402 17778 6414
rect 18398 6466 18450 6478
rect 18398 6402 18450 6414
rect 19966 6466 20018 6478
rect 20750 6466 20802 6478
rect 20402 6414 20414 6466
rect 20466 6414 20478 6466
rect 19966 6402 20018 6414
rect 20750 6402 20802 6414
rect 22094 6466 22146 6478
rect 22094 6402 22146 6414
rect 22990 6466 23042 6478
rect 29486 6466 29538 6478
rect 23762 6414 23774 6466
rect 23826 6414 23838 6466
rect 22990 6402 23042 6414
rect 29486 6402 29538 6414
rect 30494 6466 30546 6478
rect 33182 6466 33234 6478
rect 36094 6466 36146 6478
rect 31826 6414 31838 6466
rect 31890 6414 31902 6466
rect 34066 6414 34078 6466
rect 34130 6414 34142 6466
rect 30494 6402 30546 6414
rect 33182 6402 33234 6414
rect 36094 6402 36146 6414
rect 37438 6466 37490 6478
rect 37438 6402 37490 6414
rect 40238 6466 40290 6478
rect 40238 6402 40290 6414
rect 40910 6466 40962 6478
rect 40910 6402 40962 6414
rect 46174 6466 46226 6478
rect 46174 6402 46226 6414
rect 46398 6466 46450 6478
rect 46398 6402 46450 6414
rect 46958 6466 47010 6478
rect 46958 6402 47010 6414
rect 47630 6466 47682 6478
rect 47630 6402 47682 6414
rect 1344 6298 48608 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 48608 6298
rect 1344 6212 48608 6246
rect 3502 6130 3554 6142
rect 9774 6130 9826 6142
rect 7074 6078 7086 6130
rect 7138 6078 7150 6130
rect 3502 6066 3554 6078
rect 9774 6066 9826 6078
rect 13470 6130 13522 6142
rect 13470 6066 13522 6078
rect 14478 6130 14530 6142
rect 14478 6066 14530 6078
rect 16382 6130 16434 6142
rect 16382 6066 16434 6078
rect 16718 6130 16770 6142
rect 16718 6066 16770 6078
rect 16830 6130 16882 6142
rect 16830 6066 16882 6078
rect 17502 6130 17554 6142
rect 17502 6066 17554 6078
rect 19294 6130 19346 6142
rect 19294 6066 19346 6078
rect 20974 6130 21026 6142
rect 20974 6066 21026 6078
rect 22094 6130 22146 6142
rect 22094 6066 22146 6078
rect 22990 6130 23042 6142
rect 22990 6066 23042 6078
rect 23886 6130 23938 6142
rect 23886 6066 23938 6078
rect 24334 6130 24386 6142
rect 28366 6130 28418 6142
rect 26114 6078 26126 6130
rect 26178 6078 26190 6130
rect 24334 6066 24386 6078
rect 28366 6066 28418 6078
rect 29934 6130 29986 6142
rect 29934 6066 29986 6078
rect 31726 6130 31778 6142
rect 31726 6066 31778 6078
rect 34750 6130 34802 6142
rect 34750 6066 34802 6078
rect 35198 6130 35250 6142
rect 35198 6066 35250 6078
rect 36206 6130 36258 6142
rect 36206 6066 36258 6078
rect 37214 6130 37266 6142
rect 37214 6066 37266 6078
rect 37662 6130 37714 6142
rect 37662 6066 37714 6078
rect 39342 6130 39394 6142
rect 39342 6066 39394 6078
rect 40238 6130 40290 6142
rect 40238 6066 40290 6078
rect 44718 6130 44770 6142
rect 44718 6066 44770 6078
rect 8430 6018 8482 6030
rect 8430 5954 8482 5966
rect 11006 6018 11058 6030
rect 11006 5954 11058 5966
rect 11454 6018 11506 6030
rect 11454 5954 11506 5966
rect 13694 6018 13746 6030
rect 13694 5954 13746 5966
rect 22542 6018 22594 6030
rect 24558 6018 24610 6030
rect 23314 5966 23326 6018
rect 23378 5966 23390 6018
rect 22542 5954 22594 5966
rect 24558 5954 24610 5966
rect 25566 6018 25618 6030
rect 25566 5954 25618 5966
rect 27134 6018 27186 6030
rect 27134 5954 27186 5966
rect 27694 6018 27746 6030
rect 27694 5954 27746 5966
rect 28590 6018 28642 6030
rect 28590 5954 28642 5966
rect 29262 6018 29314 6030
rect 29262 5954 29314 5966
rect 31950 6018 32002 6030
rect 31950 5954 32002 5966
rect 33518 6018 33570 6030
rect 33966 6018 34018 6030
rect 39566 6018 39618 6030
rect 33730 5966 33742 6018
rect 33794 5966 33806 6018
rect 36418 5966 36430 6018
rect 36482 5966 36494 6018
rect 33518 5954 33570 5966
rect 33966 5954 34018 5966
rect 39566 5954 39618 5966
rect 44382 6018 44434 6030
rect 44382 5954 44434 5966
rect 44494 6018 44546 6030
rect 46050 5966 46062 6018
rect 46114 5966 46126 6018
rect 44494 5954 44546 5966
rect 7422 5906 7474 5918
rect 3826 5854 3838 5906
rect 3890 5854 3902 5906
rect 7422 5842 7474 5854
rect 7646 5906 7698 5918
rect 7646 5842 7698 5854
rect 7982 5906 8034 5918
rect 7982 5842 8034 5854
rect 8094 5906 8146 5918
rect 8766 5906 8818 5918
rect 9998 5906 10050 5918
rect 8642 5854 8654 5906
rect 8706 5854 8718 5906
rect 8978 5854 8990 5906
rect 9042 5854 9054 5906
rect 8094 5842 8146 5854
rect 8766 5842 8818 5854
rect 9998 5842 10050 5854
rect 10222 5906 10274 5918
rect 10222 5842 10274 5854
rect 10670 5906 10722 5918
rect 11342 5906 11394 5918
rect 11218 5854 11230 5906
rect 11282 5854 11294 5906
rect 10670 5842 10722 5854
rect 11342 5842 11394 5854
rect 12910 5906 12962 5918
rect 12910 5842 12962 5854
rect 13134 5906 13186 5918
rect 13134 5842 13186 5854
rect 14142 5906 14194 5918
rect 14142 5842 14194 5854
rect 14254 5906 14306 5918
rect 14254 5842 14306 5854
rect 14702 5906 14754 5918
rect 14702 5842 14754 5854
rect 14926 5906 14978 5918
rect 14926 5842 14978 5854
rect 15486 5906 15538 5918
rect 15486 5842 15538 5854
rect 15598 5906 15650 5918
rect 15598 5842 15650 5854
rect 16046 5906 16098 5918
rect 16046 5842 16098 5854
rect 16606 5906 16658 5918
rect 16606 5842 16658 5854
rect 17614 5906 17666 5918
rect 17614 5842 17666 5854
rect 17726 5906 17778 5918
rect 18622 5906 18674 5918
rect 18050 5854 18062 5906
rect 18114 5854 18126 5906
rect 17726 5842 17778 5854
rect 18622 5842 18674 5854
rect 19070 5906 19122 5918
rect 19070 5842 19122 5854
rect 19966 5906 20018 5918
rect 19966 5842 20018 5854
rect 20190 5906 20242 5918
rect 20190 5842 20242 5854
rect 21534 5906 21586 5918
rect 21534 5842 21586 5854
rect 22318 5906 22370 5918
rect 22318 5842 22370 5854
rect 24110 5906 24162 5918
rect 24110 5842 24162 5854
rect 25118 5906 25170 5918
rect 25118 5842 25170 5854
rect 25342 5906 25394 5918
rect 25342 5842 25394 5854
rect 25790 5906 25842 5918
rect 27358 5906 27410 5918
rect 26338 5854 26350 5906
rect 26402 5854 26414 5906
rect 25790 5842 25842 5854
rect 27358 5842 27410 5854
rect 27918 5906 27970 5918
rect 27918 5842 27970 5854
rect 28478 5906 28530 5918
rect 28478 5842 28530 5854
rect 28814 5906 28866 5918
rect 28814 5842 28866 5854
rect 29374 5906 29426 5918
rect 29374 5842 29426 5854
rect 30382 5906 30434 5918
rect 30382 5842 30434 5854
rect 30606 5906 30658 5918
rect 30606 5842 30658 5854
rect 31054 5906 31106 5918
rect 31054 5842 31106 5854
rect 31502 5906 31554 5918
rect 31502 5842 31554 5854
rect 31614 5906 31666 5918
rect 31614 5842 31666 5854
rect 33070 5906 33122 5918
rect 33070 5842 33122 5854
rect 34414 5906 34466 5918
rect 34414 5842 34466 5854
rect 35758 5906 35810 5918
rect 35758 5842 35810 5854
rect 36654 5906 36706 5918
rect 41010 5854 41022 5906
rect 41074 5854 41086 5906
rect 45266 5854 45278 5906
rect 45330 5854 45342 5906
rect 36654 5842 36706 5854
rect 10110 5794 10162 5806
rect 4610 5742 4622 5794
rect 4674 5742 4686 5794
rect 6738 5742 6750 5794
rect 6802 5742 6814 5794
rect 10110 5730 10162 5742
rect 12350 5794 12402 5806
rect 12350 5730 12402 5742
rect 13582 5794 13634 5806
rect 13582 5730 13634 5742
rect 15822 5794 15874 5806
rect 15822 5730 15874 5742
rect 19182 5794 19234 5806
rect 21758 5794 21810 5806
rect 19618 5742 19630 5794
rect 19682 5742 19694 5794
rect 21186 5742 21198 5794
rect 21250 5742 21262 5794
rect 19182 5730 19234 5742
rect 21758 5730 21810 5742
rect 22206 5794 22258 5806
rect 22206 5730 22258 5742
rect 24222 5794 24274 5806
rect 24222 5730 24274 5742
rect 27246 5794 27298 5806
rect 27246 5730 27298 5742
rect 29038 5794 29090 5806
rect 29038 5730 29090 5742
rect 30830 5794 30882 5806
rect 30830 5730 30882 5742
rect 32510 5794 32562 5806
rect 34066 5742 34078 5794
rect 34130 5742 34142 5794
rect 36754 5742 36766 5794
rect 36818 5742 36830 5794
rect 41794 5742 41806 5794
rect 41858 5742 41870 5794
rect 43922 5742 43934 5794
rect 43986 5742 43998 5794
rect 48178 5742 48190 5794
rect 48242 5742 48254 5794
rect 32510 5730 32562 5742
rect 10558 5682 10610 5694
rect 33182 5682 33234 5694
rect 12562 5630 12574 5682
rect 12626 5630 12638 5682
rect 10558 5618 10610 5630
rect 33182 5618 33234 5630
rect 35870 5682 35922 5694
rect 35870 5618 35922 5630
rect 39678 5682 39730 5694
rect 39678 5618 39730 5630
rect 1344 5514 48608 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 48608 5514
rect 1344 5428 48608 5462
rect 5630 5346 5682 5358
rect 5630 5282 5682 5294
rect 6638 5346 6690 5358
rect 6638 5282 6690 5294
rect 7310 5346 7362 5358
rect 7310 5282 7362 5294
rect 7422 5346 7474 5358
rect 7422 5282 7474 5294
rect 13470 5346 13522 5358
rect 19630 5346 19682 5358
rect 18722 5294 18734 5346
rect 18786 5343 18798 5346
rect 19282 5343 19294 5346
rect 18786 5297 19294 5343
rect 18786 5294 18798 5297
rect 19282 5294 19294 5297
rect 19346 5294 19358 5346
rect 13470 5282 13522 5294
rect 19630 5282 19682 5294
rect 19742 5346 19794 5358
rect 19742 5282 19794 5294
rect 22094 5346 22146 5358
rect 23774 5346 23826 5358
rect 23426 5294 23438 5346
rect 23490 5294 23502 5346
rect 22094 5282 22146 5294
rect 23774 5282 23826 5294
rect 24334 5346 24386 5358
rect 24334 5282 24386 5294
rect 24446 5346 24498 5358
rect 24446 5282 24498 5294
rect 33854 5346 33906 5358
rect 33854 5282 33906 5294
rect 4622 5234 4674 5246
rect 4622 5170 4674 5182
rect 5070 5234 5122 5246
rect 5070 5170 5122 5182
rect 5742 5234 5794 5246
rect 5742 5170 5794 5182
rect 6414 5234 6466 5246
rect 12462 5234 12514 5246
rect 18846 5234 18898 5246
rect 11666 5182 11678 5234
rect 11730 5182 11742 5234
rect 16146 5182 16158 5234
rect 16210 5182 16222 5234
rect 18274 5182 18286 5234
rect 18338 5182 18350 5234
rect 6414 5170 6466 5182
rect 12462 5170 12514 5182
rect 18846 5170 18898 5182
rect 19294 5234 19346 5246
rect 29262 5234 29314 5246
rect 26450 5182 26462 5234
rect 26514 5182 26526 5234
rect 28578 5182 28590 5234
rect 28642 5182 28654 5234
rect 19294 5170 19346 5182
rect 29262 5170 29314 5182
rect 30158 5234 30210 5246
rect 35086 5234 35138 5246
rect 33394 5182 33406 5234
rect 33458 5182 33470 5234
rect 34626 5182 34638 5234
rect 34690 5182 34702 5234
rect 30158 5170 30210 5182
rect 35086 5170 35138 5182
rect 35646 5234 35698 5246
rect 35646 5170 35698 5182
rect 35982 5234 36034 5246
rect 35982 5170 36034 5182
rect 37102 5234 37154 5246
rect 42478 5234 42530 5246
rect 40002 5182 40014 5234
rect 40066 5182 40078 5234
rect 42130 5182 42142 5234
rect 42194 5182 42206 5234
rect 37102 5170 37154 5182
rect 42478 5170 42530 5182
rect 45390 5234 45442 5246
rect 45390 5170 45442 5182
rect 8094 5122 8146 5134
rect 6962 5070 6974 5122
rect 7026 5070 7038 5122
rect 7970 5070 7982 5122
rect 8034 5070 8046 5122
rect 8094 5058 8146 5070
rect 8206 5122 8258 5134
rect 12014 5122 12066 5134
rect 8754 5070 8766 5122
rect 8818 5070 8830 5122
rect 9538 5070 9550 5122
rect 9602 5070 9614 5122
rect 8206 5058 8258 5070
rect 12014 5058 12066 5070
rect 12350 5122 12402 5134
rect 12350 5058 12402 5070
rect 12574 5122 12626 5134
rect 12574 5058 12626 5070
rect 13582 5122 13634 5134
rect 13582 5058 13634 5070
rect 14366 5122 14418 5134
rect 20414 5122 20466 5134
rect 22206 5122 22258 5134
rect 23998 5122 24050 5134
rect 29150 5122 29202 5134
rect 33742 5122 33794 5134
rect 36990 5122 37042 5134
rect 46510 5122 46562 5134
rect 15474 5070 15486 5122
rect 15538 5070 15550 5122
rect 20626 5070 20638 5122
rect 20690 5070 20702 5122
rect 23090 5070 23102 5122
rect 23154 5070 23166 5122
rect 25330 5070 25342 5122
rect 25394 5070 25406 5122
rect 25778 5070 25790 5122
rect 25842 5070 25854 5122
rect 29698 5070 29710 5122
rect 29762 5070 29774 5122
rect 30482 5070 30494 5122
rect 30546 5070 30558 5122
rect 34402 5070 34414 5122
rect 34466 5070 34478 5122
rect 34738 5070 34750 5122
rect 34802 5070 34814 5122
rect 39218 5070 39230 5122
rect 39282 5070 39294 5122
rect 14366 5058 14418 5070
rect 20414 5058 20466 5070
rect 22206 5058 22258 5070
rect 23998 5058 24050 5070
rect 29150 5058 29202 5070
rect 33742 5058 33794 5070
rect 36990 5058 37042 5070
rect 46510 5058 46562 5070
rect 46958 5122 47010 5134
rect 46958 5058 47010 5070
rect 47070 5122 47122 5134
rect 47070 5058 47122 5070
rect 47518 5122 47570 5134
rect 47518 5058 47570 5070
rect 47854 5122 47906 5134
rect 47854 5058 47906 5070
rect 7758 5010 7810 5022
rect 7758 4946 7810 4958
rect 13806 5010 13858 5022
rect 19966 5010 20018 5022
rect 22542 5010 22594 5022
rect 24782 5010 24834 5022
rect 29374 5010 29426 5022
rect 34078 5010 34130 5022
rect 14130 4958 14142 5010
rect 14194 4958 14206 5010
rect 20290 4958 20302 5010
rect 20354 4958 20366 5010
rect 22754 4958 22766 5010
rect 22818 4958 22830 5010
rect 24994 4958 25006 5010
rect 25058 4958 25070 5010
rect 31266 4958 31278 5010
rect 31330 4958 31342 5010
rect 13806 4946 13858 4958
rect 19966 4946 20018 4958
rect 22542 4946 22594 4958
rect 24782 4946 24834 4958
rect 29374 4946 29426 4958
rect 34078 4946 34130 4958
rect 38894 5010 38946 5022
rect 38894 4946 38946 4958
rect 47630 5010 47682 5022
rect 47630 4946 47682 4958
rect 14254 4898 14306 4910
rect 14254 4834 14306 4846
rect 15038 4898 15090 4910
rect 15038 4834 15090 4846
rect 21422 4898 21474 4910
rect 21422 4834 21474 4846
rect 22878 4898 22930 4910
rect 22878 4834 22930 4846
rect 25118 4898 25170 4910
rect 25118 4834 25170 4846
rect 35198 4898 35250 4910
rect 35198 4834 35250 4846
rect 36094 4898 36146 4910
rect 36094 4834 36146 4846
rect 42590 4898 42642 4910
rect 42590 4834 42642 4846
rect 43038 4898 43090 4910
rect 43038 4834 43090 4846
rect 44158 4898 44210 4910
rect 44158 4834 44210 4846
rect 44942 4898 44994 4910
rect 44942 4834 44994 4846
rect 46734 4898 46786 4910
rect 46734 4834 46786 4846
rect 1344 4730 48608 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 48608 4730
rect 1344 4644 48608 4678
rect 5294 4562 5346 4574
rect 5294 4498 5346 4510
rect 5854 4562 5906 4574
rect 5854 4498 5906 4510
rect 9886 4562 9938 4574
rect 9886 4498 9938 4510
rect 10222 4562 10274 4574
rect 10222 4498 10274 4510
rect 24110 4562 24162 4574
rect 24110 4498 24162 4510
rect 24558 4562 24610 4574
rect 24558 4498 24610 4510
rect 25790 4562 25842 4574
rect 25790 4498 25842 4510
rect 26238 4562 26290 4574
rect 26238 4498 26290 4510
rect 26798 4562 26850 4574
rect 26798 4498 26850 4510
rect 30718 4562 30770 4574
rect 30718 4498 30770 4510
rect 31278 4562 31330 4574
rect 31278 4498 31330 4510
rect 31726 4562 31778 4574
rect 31726 4498 31778 4510
rect 31838 4562 31890 4574
rect 31838 4498 31890 4510
rect 40126 4562 40178 4574
rect 40126 4498 40178 4510
rect 41246 4562 41298 4574
rect 41246 4498 41298 4510
rect 44942 4562 44994 4574
rect 44942 4498 44994 4510
rect 25230 4450 25282 4462
rect 31390 4450 31442 4462
rect 39566 4450 39618 4462
rect 16034 4398 16046 4450
rect 16098 4398 16110 4450
rect 28130 4398 28142 4450
rect 28194 4398 28206 4450
rect 35186 4398 35198 4450
rect 35250 4398 35262 4450
rect 38434 4398 38446 4450
rect 38498 4398 38510 4450
rect 25230 4386 25282 4398
rect 31390 4386 31442 4398
rect 39566 4386 39618 4398
rect 41134 4450 41186 4462
rect 43698 4398 43710 4450
rect 43762 4398 43774 4450
rect 46050 4398 46062 4450
rect 46114 4398 46126 4450
rect 41134 4386 41186 4398
rect 31950 4338 32002 4350
rect 6178 4286 6190 4338
rect 6242 4286 6254 4338
rect 13570 4286 13582 4338
rect 13634 4286 13646 4338
rect 16818 4286 16830 4338
rect 16882 4286 16894 4338
rect 17602 4286 17614 4338
rect 17666 4286 17678 4338
rect 20738 4286 20750 4338
rect 20802 4286 20814 4338
rect 27458 4286 27470 4338
rect 27522 4286 27534 4338
rect 32274 4286 32286 4338
rect 32338 4286 32350 4338
rect 35970 4286 35982 4338
rect 36034 4286 36046 4338
rect 39106 4286 39118 4338
rect 39170 4286 39182 4338
rect 44370 4286 44382 4338
rect 44434 4286 44446 4338
rect 45266 4286 45278 4338
rect 45330 4286 45342 4338
rect 31950 4274 32002 4286
rect 10334 4226 10386 4238
rect 6850 4174 6862 4226
rect 6914 4174 6926 4226
rect 8978 4174 8990 4226
rect 9042 4174 9054 4226
rect 10658 4174 10670 4226
rect 10722 4174 10734 4226
rect 12786 4174 12798 4226
rect 12850 4174 12862 4226
rect 13906 4174 13918 4226
rect 13970 4174 13982 4226
rect 18274 4174 18286 4226
rect 18338 4174 18350 4226
rect 20402 4174 20414 4226
rect 20466 4174 20478 4226
rect 21522 4174 21534 4226
rect 21586 4174 21598 4226
rect 23650 4174 23662 4226
rect 23714 4174 23726 4226
rect 30258 4174 30270 4226
rect 30322 4174 30334 4226
rect 33058 4174 33070 4226
rect 33122 4174 33134 4226
rect 36306 4174 36318 4226
rect 36370 4174 36382 4226
rect 41570 4174 41582 4226
rect 41634 4174 41646 4226
rect 48178 4174 48190 4226
rect 48242 4174 48254 4226
rect 10334 4162 10386 4174
rect 25342 4114 25394 4126
rect 25342 4050 25394 4062
rect 39678 4114 39730 4126
rect 39678 4050 39730 4062
rect 1344 3946 48608 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 48608 3946
rect 1344 3860 48608 3894
rect 7534 3778 7586 3790
rect 13134 3778 13186 3790
rect 19518 3778 19570 3790
rect 10322 3726 10334 3778
rect 10386 3775 10398 3778
rect 11218 3775 11230 3778
rect 10386 3729 11230 3775
rect 10386 3726 10398 3729
rect 11218 3726 11230 3729
rect 11282 3726 11294 3778
rect 17602 3726 17614 3778
rect 17666 3775 17678 3778
rect 18834 3775 18846 3778
rect 17666 3729 18846 3775
rect 17666 3726 17678 3729
rect 18834 3726 18846 3729
rect 18898 3726 18910 3778
rect 7534 3714 7586 3726
rect 13134 3714 13186 3726
rect 19518 3714 19570 3726
rect 22094 3778 22146 3790
rect 22418 3726 22430 3778
rect 22482 3775 22494 3778
rect 22866 3775 22878 3778
rect 22482 3729 22878 3775
rect 22482 3726 22494 3729
rect 22866 3726 22878 3729
rect 22930 3726 22942 3778
rect 22094 3714 22146 3726
rect 6414 3666 6466 3678
rect 6414 3602 6466 3614
rect 6862 3666 6914 3678
rect 6862 3602 6914 3614
rect 7310 3666 7362 3678
rect 7310 3602 7362 3614
rect 7646 3666 7698 3678
rect 7646 3602 7698 3614
rect 8430 3666 8482 3678
rect 8430 3602 8482 3614
rect 8878 3666 8930 3678
rect 8878 3602 8930 3614
rect 9998 3666 10050 3678
rect 9998 3602 10050 3614
rect 10446 3666 10498 3678
rect 10446 3602 10498 3614
rect 11342 3666 11394 3678
rect 11342 3602 11394 3614
rect 12238 3666 12290 3678
rect 12238 3602 12290 3614
rect 13246 3666 13298 3678
rect 13246 3602 13298 3614
rect 14142 3666 14194 3678
rect 14142 3602 14194 3614
rect 14590 3666 14642 3678
rect 14590 3602 14642 3614
rect 15038 3666 15090 3678
rect 15038 3602 15090 3614
rect 15822 3666 15874 3678
rect 15822 3602 15874 3614
rect 16494 3666 16546 3678
rect 16494 3602 16546 3614
rect 17726 3666 17778 3678
rect 17726 3602 17778 3614
rect 18398 3666 18450 3678
rect 18398 3602 18450 3614
rect 18846 3666 18898 3678
rect 18846 3602 18898 3614
rect 19294 3666 19346 3678
rect 19294 3602 19346 3614
rect 19630 3666 19682 3678
rect 19630 3602 19682 3614
rect 20078 3666 20130 3678
rect 20078 3602 20130 3614
rect 20974 3666 21026 3678
rect 20974 3602 21026 3614
rect 21422 3666 21474 3678
rect 21422 3602 21474 3614
rect 21870 3666 21922 3678
rect 21870 3602 21922 3614
rect 22206 3666 22258 3678
rect 22206 3602 22258 3614
rect 22766 3666 22818 3678
rect 22766 3602 22818 3614
rect 23214 3666 23266 3678
rect 23214 3602 23266 3614
rect 24110 3666 24162 3678
rect 28590 3666 28642 3678
rect 25330 3614 25342 3666
rect 25394 3614 25406 3666
rect 27458 3614 27470 3666
rect 27522 3614 27534 3666
rect 24110 3602 24162 3614
rect 28590 3602 28642 3614
rect 35534 3666 35586 3678
rect 43822 3666 43874 3678
rect 36754 3614 36766 3666
rect 36818 3614 36830 3666
rect 38882 3614 38894 3666
rect 38946 3614 38958 3666
rect 39778 3614 39790 3666
rect 39842 3614 39854 3666
rect 41906 3614 41918 3666
rect 41970 3614 41982 3666
rect 35534 3602 35586 3614
rect 43822 3602 43874 3614
rect 45054 3666 45106 3678
rect 45054 3602 45106 3614
rect 23662 3554 23714 3566
rect 47630 3554 47682 3566
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 35970 3502 35982 3554
rect 36034 3502 36046 3554
rect 42578 3502 42590 3554
rect 42642 3502 42654 3554
rect 23662 3490 23714 3502
rect 47630 3490 47682 3502
rect 9550 3442 9602 3454
rect 9550 3378 9602 3390
rect 10894 3442 10946 3454
rect 10894 3378 10946 3390
rect 11790 3442 11842 3454
rect 11790 3378 11842 3390
rect 12686 3442 12738 3454
rect 12686 3378 12738 3390
rect 17390 3442 17442 3454
rect 17390 3378 17442 3390
rect 46958 3442 47010 3454
rect 46958 3378 47010 3390
rect 48190 3442 48242 3454
rect 48190 3378 48242 3390
rect 1344 3162 48608 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 48608 3162
rect 1344 3076 48608 3110
<< via1 >>
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 19182 46062 19234 46114
rect 22094 46062 22146 46114
rect 25230 46062 25282 46114
rect 36990 46062 37042 46114
rect 44606 46062 44658 46114
rect 16046 45950 16098 46002
rect 30270 45950 30322 46002
rect 35086 45950 35138 46002
rect 40350 45950 40402 46002
rect 46846 45950 46898 46002
rect 9662 45838 9714 45890
rect 13134 45838 13186 45890
rect 19742 45838 19794 45890
rect 21086 45838 21138 45890
rect 27134 45838 27186 45890
rect 31166 45838 31218 45890
rect 32174 45838 32226 45890
rect 35982 45838 36034 45890
rect 38894 45838 38946 45890
rect 42366 45838 42418 45890
rect 43934 45838 43986 45890
rect 47966 45838 48018 45890
rect 3838 45726 3890 45778
rect 5518 45726 5570 45778
rect 6974 45726 7026 45778
rect 8542 45726 8594 45778
rect 9326 45726 9378 45778
rect 10110 45726 10162 45778
rect 11678 45726 11730 45778
rect 12574 45726 12626 45778
rect 13918 45726 13970 45778
rect 16942 45726 16994 45778
rect 27470 45726 27522 45778
rect 28702 45726 28754 45778
rect 32958 45726 33010 45778
rect 39230 45726 39282 45778
rect 42702 45726 42754 45778
rect 46510 45726 46562 45778
rect 7982 45614 8034 45666
rect 9438 45614 9490 45666
rect 10894 45614 10946 45666
rect 11342 45614 11394 45666
rect 39118 45614 39170 45666
rect 42814 45614 42866 45666
rect 42926 45614 42978 45666
rect 46734 45614 46786 45666
rect 47406 45614 47458 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 13022 45278 13074 45330
rect 24446 45278 24498 45330
rect 26686 45278 26738 45330
rect 30942 45278 30994 45330
rect 39678 45278 39730 45330
rect 2942 45166 2994 45218
rect 5630 45166 5682 45218
rect 8206 45166 8258 45218
rect 25454 45166 25506 45218
rect 44830 45166 44882 45218
rect 47406 45166 47458 45218
rect 3278 45054 3330 45106
rect 3390 45054 3442 45106
rect 4958 45054 5010 45106
rect 9550 45054 9602 45106
rect 12686 45054 12738 45106
rect 13022 45054 13074 45106
rect 13246 45054 13298 45106
rect 14030 45054 14082 45106
rect 17502 45054 17554 45106
rect 17950 45054 18002 45106
rect 21086 45054 21138 45106
rect 24334 45054 24386 45106
rect 24670 45054 24722 45106
rect 25566 45054 25618 45106
rect 26350 45054 26402 45106
rect 29934 45054 29986 45106
rect 32510 45054 32562 45106
rect 33182 45054 33234 45106
rect 36430 45054 36482 45106
rect 39902 45054 39954 45106
rect 40238 45054 40290 45106
rect 41022 45054 41074 45106
rect 44158 45054 44210 45106
rect 44606 45054 44658 45106
rect 44942 45054 44994 45106
rect 48190 45054 48242 45106
rect 3054 44942 3106 44994
rect 7758 44942 7810 44994
rect 8990 44942 9042 44994
rect 10334 44942 10386 44994
rect 12462 44942 12514 44994
rect 14702 44942 14754 44994
rect 16830 44942 16882 44994
rect 18622 44942 18674 44994
rect 20750 44942 20802 44994
rect 21870 44942 21922 44994
rect 23998 44942 24050 44994
rect 26126 44942 26178 44994
rect 27134 44942 27186 44994
rect 29262 44942 29314 44994
rect 30494 44942 30546 44994
rect 31390 44942 31442 44994
rect 31950 44942 32002 44994
rect 33966 44942 34018 44994
rect 36094 44942 36146 44994
rect 37214 44942 37266 44994
rect 39342 44942 39394 44994
rect 39790 44942 39842 44994
rect 41694 44942 41746 44994
rect 43822 44942 43874 44994
rect 45278 44942 45330 44994
rect 8094 44830 8146 44882
rect 8430 44830 8482 44882
rect 25454 44830 25506 44882
rect 26014 44830 26066 44882
rect 44382 44830 44434 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 15374 44494 15426 44546
rect 21310 44494 21362 44546
rect 33742 44494 33794 44546
rect 37214 44494 37266 44546
rect 45838 44494 45890 44546
rect 2606 44382 2658 44434
rect 4734 44382 4786 44434
rect 6190 44382 6242 44434
rect 9102 44382 9154 44434
rect 10222 44382 10274 44434
rect 19630 44382 19682 44434
rect 26014 44382 26066 44434
rect 32398 44382 32450 44434
rect 36318 44382 36370 44434
rect 44270 44382 44322 44434
rect 1934 44270 1986 44322
rect 7758 44270 7810 44322
rect 8654 44270 8706 44322
rect 9662 44270 9714 44322
rect 12238 44270 12290 44322
rect 16046 44270 16098 44322
rect 16830 44270 16882 44322
rect 24222 44270 24274 44322
rect 24558 44270 24610 44322
rect 25454 44270 25506 44322
rect 26910 44270 26962 44322
rect 27134 44270 27186 44322
rect 28366 44270 28418 44322
rect 29598 44270 29650 44322
rect 32734 44270 32786 44322
rect 35982 44270 36034 44322
rect 39118 44270 39170 44322
rect 40014 44270 40066 44322
rect 40350 44270 40402 44322
rect 41358 44270 41410 44322
rect 45054 44270 45106 44322
rect 5742 44158 5794 44210
rect 5854 44158 5906 44210
rect 6302 44158 6354 44210
rect 7422 44158 7474 44210
rect 9550 44158 9602 44210
rect 10334 44158 10386 44210
rect 10670 44158 10722 44210
rect 10894 44158 10946 44210
rect 12574 44158 12626 44210
rect 17502 44158 17554 44210
rect 21422 44158 21474 44210
rect 23326 44158 23378 44210
rect 27806 44158 27858 44210
rect 28254 44158 28306 44210
rect 30270 44158 30322 44210
rect 39902 44158 39954 44210
rect 42142 44158 42194 44210
rect 47742 44158 47794 44210
rect 48078 44158 48130 44210
rect 5518 44046 5570 44098
rect 9326 44046 9378 44098
rect 10110 44046 10162 44098
rect 20078 44046 20130 44098
rect 20526 44046 20578 44098
rect 21870 44046 21922 44098
rect 22318 44046 22370 44098
rect 22990 44046 23042 44098
rect 26462 44046 26514 44098
rect 28030 44046 28082 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 3278 43710 3330 43762
rect 3390 43710 3442 43762
rect 6526 43710 6578 43762
rect 7310 43710 7362 43762
rect 7758 43710 7810 43762
rect 9998 43710 10050 43762
rect 12574 43710 12626 43762
rect 12798 43710 12850 43762
rect 13022 43710 13074 43762
rect 13134 43710 13186 43762
rect 14814 43710 14866 43762
rect 24334 43710 24386 43762
rect 24558 43710 24610 43762
rect 25230 43710 25282 43762
rect 27806 43710 27858 43762
rect 34078 43710 34130 43762
rect 44606 43710 44658 43762
rect 4846 43598 4898 43650
rect 7198 43598 7250 43650
rect 8654 43598 8706 43650
rect 12462 43598 12514 43650
rect 13918 43598 13970 43650
rect 14030 43598 14082 43650
rect 14702 43598 14754 43650
rect 15374 43598 15426 43650
rect 20974 43598 21026 43650
rect 22766 43598 22818 43650
rect 24222 43598 24274 43650
rect 25118 43598 25170 43650
rect 25678 43598 25730 43650
rect 26574 43598 26626 43650
rect 26686 43598 26738 43650
rect 27470 43598 27522 43650
rect 27918 43598 27970 43650
rect 30942 43598 30994 43650
rect 33406 43598 33458 43650
rect 34750 43598 34802 43650
rect 34862 43598 34914 43650
rect 38334 43598 38386 43650
rect 38782 43598 38834 43650
rect 44830 43598 44882 43650
rect 3502 43486 3554 43538
rect 3838 43486 3890 43538
rect 5406 43486 5458 43538
rect 6078 43486 6130 43538
rect 6750 43486 6802 43538
rect 7870 43486 7922 43538
rect 8766 43486 8818 43538
rect 10334 43486 10386 43538
rect 13246 43486 13298 43538
rect 13582 43486 13634 43538
rect 15262 43486 15314 43538
rect 15486 43486 15538 43538
rect 15710 43486 15762 43538
rect 16158 43486 16210 43538
rect 16382 43486 16434 43538
rect 16830 43486 16882 43538
rect 17502 43486 17554 43538
rect 22654 43486 22706 43538
rect 22990 43486 23042 43538
rect 23774 43486 23826 43538
rect 25454 43486 25506 43538
rect 26462 43486 26514 43538
rect 27022 43486 27074 43538
rect 28030 43486 28082 43538
rect 28478 43486 28530 43538
rect 29038 43486 29090 43538
rect 29710 43486 29762 43538
rect 30158 43486 30210 43538
rect 31166 43486 31218 43538
rect 31614 43486 31666 43538
rect 32062 43486 32114 43538
rect 33294 43486 33346 43538
rect 33966 43486 34018 43538
rect 37550 43486 37602 43538
rect 38110 43486 38162 43538
rect 38558 43486 38610 43538
rect 39118 43486 39170 43538
rect 43038 43486 43090 43538
rect 43934 43486 43986 43538
rect 44942 43486 44994 43538
rect 48190 43486 48242 43538
rect 1822 43374 1874 43426
rect 4510 43374 4562 43426
rect 5742 43374 5794 43426
rect 6638 43374 6690 43426
rect 9662 43374 9714 43426
rect 10782 43374 10834 43426
rect 11342 43374 11394 43426
rect 11790 43374 11842 43426
rect 12238 43374 12290 43426
rect 14926 43374 14978 43426
rect 16270 43374 16322 43426
rect 18174 43374 18226 43426
rect 20302 43374 20354 43426
rect 20862 43374 20914 43426
rect 21982 43374 22034 43426
rect 22430 43374 22482 43426
rect 23438 43374 23490 43426
rect 24334 43374 24386 43426
rect 26126 43374 26178 43426
rect 29374 43374 29426 43426
rect 31054 43374 31106 43426
rect 32510 43374 32562 43426
rect 35422 43374 35474 43426
rect 38446 43374 38498 43426
rect 40014 43374 40066 43426
rect 40238 43374 40290 43426
rect 41134 43374 41186 43426
rect 44382 43374 44434 43426
rect 45278 43374 45330 43426
rect 47406 43374 47458 43426
rect 11342 43262 11394 43314
rect 12238 43262 12290 43314
rect 14030 43262 14082 43314
rect 21198 43262 21250 43314
rect 34750 43262 34802 43314
rect 39118 43262 39170 43314
rect 39454 43262 39506 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 6302 42926 6354 42978
rect 18958 42926 19010 42978
rect 22318 42926 22370 42978
rect 37102 42926 37154 42978
rect 39342 42926 39394 42978
rect 45838 42926 45890 42978
rect 3166 42814 3218 42866
rect 3726 42814 3778 42866
rect 4734 42814 4786 42866
rect 7870 42814 7922 42866
rect 9550 42814 9602 42866
rect 14142 42814 14194 42866
rect 22878 42814 22930 42866
rect 23662 42814 23714 42866
rect 29262 42814 29314 42866
rect 29486 42814 29538 42866
rect 30046 42814 30098 42866
rect 30942 42814 30994 42866
rect 34078 42814 34130 42866
rect 35310 42814 35362 42866
rect 36206 42814 36258 42866
rect 39678 42814 39730 42866
rect 43262 42814 43314 42866
rect 43710 42814 43762 42866
rect 1822 42702 1874 42754
rect 2270 42702 2322 42754
rect 4062 42702 4114 42754
rect 4846 42702 4898 42754
rect 5630 42702 5682 42754
rect 5966 42702 6018 42754
rect 6974 42702 7026 42754
rect 13694 42702 13746 42754
rect 14590 42702 14642 42754
rect 15710 42702 15762 42754
rect 17950 42702 18002 42754
rect 21422 42702 21474 42754
rect 21982 42702 22034 42754
rect 22990 42702 23042 42754
rect 26462 42702 26514 42754
rect 27694 42702 27746 42754
rect 27918 42702 27970 42754
rect 28142 42702 28194 42754
rect 30270 42702 30322 42754
rect 31278 42702 31330 42754
rect 31838 42702 31890 42754
rect 33742 42702 33794 42754
rect 34190 42702 34242 42754
rect 35534 42702 35586 42754
rect 38110 42702 38162 42754
rect 38334 42702 38386 42754
rect 42478 42702 42530 42754
rect 43934 42702 43986 42754
rect 45054 42702 45106 42754
rect 2830 42590 2882 42642
rect 3054 42590 3106 42642
rect 5742 42590 5794 42642
rect 6414 42590 6466 42642
rect 7534 42590 7586 42642
rect 7758 42590 7810 42642
rect 8654 42590 8706 42642
rect 8878 42590 8930 42642
rect 9998 42590 10050 42642
rect 11454 42590 11506 42642
rect 11678 42590 11730 42642
rect 12014 42590 12066 42642
rect 12910 42590 12962 42642
rect 16158 42590 16210 42642
rect 17390 42590 17442 42642
rect 21758 42590 21810 42642
rect 24334 42590 24386 42642
rect 25342 42590 25394 42642
rect 25790 42590 25842 42642
rect 26126 42590 26178 42642
rect 26798 42590 26850 42642
rect 37102 42590 37154 42642
rect 37214 42590 37266 42642
rect 38558 42590 38610 42642
rect 39006 42590 39058 42642
rect 41806 42590 41858 42642
rect 43150 42590 43202 42642
rect 43374 42590 43426 42642
rect 48190 42590 48242 42642
rect 6302 42478 6354 42530
rect 7086 42478 7138 42530
rect 7310 42478 7362 42530
rect 8766 42478 8818 42530
rect 12126 42478 12178 42530
rect 12350 42478 12402 42530
rect 12574 42478 12626 42530
rect 13358 42478 13410 42530
rect 13582 42478 13634 42530
rect 16942 42478 16994 42530
rect 17502 42478 17554 42530
rect 17726 42478 17778 42530
rect 21310 42478 21362 42530
rect 24446 42478 24498 42530
rect 24670 42478 24722 42530
rect 25230 42478 25282 42530
rect 26238 42478 26290 42530
rect 26686 42478 26738 42530
rect 26910 42478 26962 42530
rect 27134 42478 27186 42530
rect 27918 42478 27970 42530
rect 29486 42478 29538 42530
rect 39230 42478 39282 42530
rect 44270 42478 44322 42530
rect 47854 42478 47906 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 12126 42142 12178 42194
rect 22318 42142 22370 42194
rect 22542 42142 22594 42194
rect 23102 42142 23154 42194
rect 23326 42142 23378 42194
rect 26462 42142 26514 42194
rect 39790 42142 39842 42194
rect 19630 42030 19682 42082
rect 21198 42030 21250 42082
rect 21534 42030 21586 42082
rect 21870 42030 21922 42082
rect 22206 42030 22258 42082
rect 25230 42030 25282 42082
rect 25342 42030 25394 42082
rect 26126 42030 26178 42082
rect 26238 42030 26290 42082
rect 34638 42030 34690 42082
rect 36430 42030 36482 42082
rect 36990 42030 37042 42082
rect 37662 42030 37714 42082
rect 37998 42030 38050 42082
rect 38222 42030 38274 42082
rect 38894 42030 38946 42082
rect 41470 42030 41522 42082
rect 43374 42030 43426 42082
rect 4622 41918 4674 41970
rect 4958 41918 5010 41970
rect 5742 41918 5794 41970
rect 8318 41918 8370 41970
rect 9438 41918 9490 41970
rect 10222 41918 10274 41970
rect 13134 41918 13186 41970
rect 16830 41918 16882 41970
rect 17950 41918 18002 41970
rect 18398 41918 18450 41970
rect 18622 41918 18674 41970
rect 20526 41918 20578 41970
rect 22766 41918 22818 41970
rect 24222 41918 24274 41970
rect 24670 41918 24722 41970
rect 25566 41918 25618 41970
rect 29486 41918 29538 41970
rect 30046 41918 30098 41970
rect 30718 41918 30770 41970
rect 31950 41918 32002 41970
rect 32398 41918 32450 41970
rect 32510 41918 32562 41970
rect 33070 41918 33122 41970
rect 35870 41918 35922 41970
rect 36766 41918 36818 41970
rect 37326 41918 37378 41970
rect 37774 41918 37826 41970
rect 38782 41918 38834 41970
rect 39678 41918 39730 41970
rect 41134 41918 41186 41970
rect 42142 41918 42194 41970
rect 42702 41918 42754 41970
rect 42926 41918 42978 41970
rect 43822 41918 43874 41970
rect 44830 41918 44882 41970
rect 44942 41918 44994 41970
rect 47406 41918 47458 41970
rect 48078 41918 48130 41970
rect 1710 41806 1762 41858
rect 3838 41806 3890 41858
rect 7870 41806 7922 41858
rect 9774 41806 9826 41858
rect 10110 41806 10162 41858
rect 11566 41806 11618 41858
rect 12686 41806 12738 41858
rect 13918 41806 13970 41858
rect 16046 41806 16098 41858
rect 17502 41806 17554 41858
rect 18174 41806 18226 41858
rect 19070 41806 19122 41858
rect 23214 41806 23266 41858
rect 23774 41806 23826 41858
rect 26686 41806 26738 41858
rect 28814 41806 28866 41858
rect 30606 41806 30658 41858
rect 31166 41806 31218 41858
rect 33518 41806 33570 41858
rect 34414 41806 34466 41858
rect 36878 41806 36930 41858
rect 40238 41806 40290 41858
rect 41806 41806 41858 41858
rect 45278 41806 45330 41858
rect 11790 41694 11842 41746
rect 13470 41694 13522 41746
rect 40350 41694 40402 41746
rect 44046 41694 44098 41746
rect 44382 41694 44434 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 16046 41358 16098 41410
rect 19070 41358 19122 41410
rect 19406 41358 19458 41410
rect 22094 41358 22146 41410
rect 22878 41358 22930 41410
rect 23326 41358 23378 41410
rect 30158 41358 30210 41410
rect 30494 41358 30546 41410
rect 31502 41358 31554 41410
rect 32846 41358 32898 41410
rect 33182 41358 33234 41410
rect 44158 41358 44210 41410
rect 47070 41358 47122 41410
rect 4622 41246 4674 41298
rect 8878 41246 8930 41298
rect 10670 41246 10722 41298
rect 14590 41246 14642 41298
rect 15934 41246 15986 41298
rect 21422 41246 21474 41298
rect 22878 41246 22930 41298
rect 23326 41246 23378 41298
rect 26238 41246 26290 41298
rect 27134 41246 27186 41298
rect 27918 41246 27970 41298
rect 28590 41246 28642 41298
rect 29934 41246 29986 41298
rect 36430 41246 36482 41298
rect 37662 41246 37714 41298
rect 38334 41246 38386 41298
rect 38446 41246 38498 41298
rect 2718 41134 2770 41186
rect 4734 41134 4786 41186
rect 7534 41134 7586 41186
rect 8318 41134 8370 41186
rect 11118 41134 11170 41186
rect 11342 41134 11394 41186
rect 12462 41134 12514 41186
rect 13470 41134 13522 41186
rect 21870 41134 21922 41186
rect 25118 41134 25170 41186
rect 26686 41134 26738 41186
rect 31838 41134 31890 41186
rect 32174 41134 32226 41186
rect 33630 41134 33682 41186
rect 37438 41134 37490 41186
rect 37550 41134 37602 41186
rect 38670 41134 38722 41186
rect 39678 41134 39730 41186
rect 39902 41134 39954 41186
rect 40686 41134 40738 41186
rect 42478 41134 42530 41186
rect 42814 41134 42866 41186
rect 43486 41134 43538 41186
rect 45614 41134 45666 41186
rect 2270 41022 2322 41074
rect 3838 41022 3890 41074
rect 4062 41022 4114 41074
rect 4398 41022 4450 41074
rect 7198 41022 7250 41074
rect 11678 41022 11730 41074
rect 12798 41022 12850 41074
rect 13694 41022 13746 41074
rect 19182 41022 19234 41074
rect 23886 41022 23938 41074
rect 24110 41022 24162 41074
rect 24782 41022 24834 41074
rect 27470 41022 27522 41074
rect 27694 41022 27746 41074
rect 28030 41022 28082 41074
rect 31166 41022 31218 41074
rect 31950 41022 32002 41074
rect 33070 41022 33122 41074
rect 34302 41022 34354 41074
rect 37998 41022 38050 41074
rect 39118 41022 39170 41074
rect 41134 41022 41186 41074
rect 44942 41022 44994 41074
rect 5854 40910 5906 40962
rect 9326 40910 9378 40962
rect 9774 40910 9826 40962
rect 10110 40910 10162 40962
rect 10558 40910 10610 40962
rect 10782 40910 10834 40962
rect 11566 40910 11618 40962
rect 12238 40910 12290 40962
rect 14030 40910 14082 40962
rect 15486 40910 15538 40962
rect 15822 40910 15874 40962
rect 18286 40910 18338 40962
rect 20526 40910 20578 40962
rect 21310 40910 21362 40962
rect 21534 40910 21586 40962
rect 22318 40910 22370 40962
rect 24446 40910 24498 40962
rect 24894 40910 24946 40962
rect 25790 40910 25842 40962
rect 29598 40910 29650 40962
rect 31390 40910 31442 40962
rect 32510 40910 32562 40962
rect 37774 40910 37826 40962
rect 40798 40910 40850 40962
rect 41470 40910 41522 40962
rect 45278 40910 45330 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 2494 40574 2546 40626
rect 3278 40574 3330 40626
rect 4062 40574 4114 40626
rect 5070 40574 5122 40626
rect 7982 40574 8034 40626
rect 10110 40574 10162 40626
rect 11118 40574 11170 40626
rect 11678 40574 11730 40626
rect 16942 40574 16994 40626
rect 17726 40574 17778 40626
rect 21758 40574 21810 40626
rect 25342 40574 25394 40626
rect 25566 40574 25618 40626
rect 26238 40574 26290 40626
rect 27022 40574 27074 40626
rect 27134 40574 27186 40626
rect 27470 40574 27522 40626
rect 35982 40574 36034 40626
rect 37102 40574 37154 40626
rect 38334 40574 38386 40626
rect 38558 40574 38610 40626
rect 38782 40574 38834 40626
rect 39230 40574 39282 40626
rect 40238 40574 40290 40626
rect 46510 40574 46562 40626
rect 46958 40574 47010 40626
rect 47630 40574 47682 40626
rect 2270 40462 2322 40514
rect 2606 40462 2658 40514
rect 2830 40462 2882 40514
rect 3390 40462 3442 40514
rect 6974 40462 7026 40514
rect 9550 40462 9602 40514
rect 10782 40462 10834 40514
rect 10894 40462 10946 40514
rect 11006 40462 11058 40514
rect 12014 40462 12066 40514
rect 12574 40462 12626 40514
rect 13470 40462 13522 40514
rect 16718 40462 16770 40514
rect 17614 40462 17666 40514
rect 23102 40462 23154 40514
rect 24110 40462 24162 40514
rect 25790 40462 25842 40514
rect 25902 40462 25954 40514
rect 29150 40462 29202 40514
rect 30158 40462 30210 40514
rect 32510 40462 32562 40514
rect 33070 40462 33122 40514
rect 35534 40462 35586 40514
rect 35870 40462 35922 40514
rect 36206 40462 36258 40514
rect 36430 40462 36482 40514
rect 36878 40462 36930 40514
rect 39790 40462 39842 40514
rect 40350 40462 40402 40514
rect 41694 40462 41746 40514
rect 44158 40462 44210 40514
rect 46286 40462 46338 40514
rect 47406 40462 47458 40514
rect 47854 40462 47906 40514
rect 3166 40350 3218 40402
rect 3726 40350 3778 40402
rect 6862 40350 6914 40402
rect 7198 40350 7250 40402
rect 7422 40350 7474 40402
rect 8654 40350 8706 40402
rect 9102 40350 9154 40402
rect 11230 40350 11282 40402
rect 11566 40350 11618 40402
rect 11790 40350 11842 40402
rect 13134 40350 13186 40402
rect 15262 40350 15314 40402
rect 15710 40350 15762 40402
rect 16606 40350 16658 40402
rect 17502 40350 17554 40402
rect 18062 40350 18114 40402
rect 18398 40350 18450 40402
rect 21982 40350 22034 40402
rect 22990 40350 23042 40402
rect 24446 40350 24498 40402
rect 26462 40350 26514 40402
rect 27246 40350 27298 40402
rect 27918 40350 27970 40402
rect 28590 40350 28642 40402
rect 30270 40350 30322 40402
rect 31166 40350 31218 40402
rect 33294 40350 33346 40402
rect 33742 40350 33794 40402
rect 35086 40350 35138 40402
rect 36766 40350 36818 40402
rect 37326 40350 37378 40402
rect 38446 40350 38498 40402
rect 40014 40350 40066 40402
rect 41022 40350 41074 40402
rect 44494 40350 44546 40402
rect 44942 40350 44994 40402
rect 45502 40350 45554 40402
rect 45838 40350 45890 40402
rect 47070 40350 47122 40402
rect 47518 40350 47570 40402
rect 4622 40238 4674 40290
rect 13582 40238 13634 40290
rect 14478 40238 14530 40290
rect 16270 40238 16322 40290
rect 19070 40238 19122 40290
rect 21198 40238 21250 40290
rect 29038 40238 29090 40290
rect 35198 40238 35250 40290
rect 37774 40238 37826 40290
rect 43822 40238 43874 40290
rect 4398 40126 4450 40178
rect 7646 40126 7698 40178
rect 9774 40126 9826 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 11790 39790 11842 39842
rect 21422 39790 21474 39842
rect 21758 39790 21810 39842
rect 25006 39790 25058 39842
rect 28254 39790 28306 39842
rect 36318 39790 36370 39842
rect 2494 39678 2546 39730
rect 4622 39678 4674 39730
rect 8542 39678 8594 39730
rect 9662 39678 9714 39730
rect 16942 39678 16994 39730
rect 19406 39678 19458 39730
rect 19966 39678 20018 39730
rect 20638 39678 20690 39730
rect 24558 39678 24610 39730
rect 26014 39678 26066 39730
rect 27358 39678 27410 39730
rect 27806 39678 27858 39730
rect 29262 39678 29314 39730
rect 33406 39678 33458 39730
rect 35086 39678 35138 39730
rect 35982 39678 36034 39730
rect 37550 39678 37602 39730
rect 38222 39678 38274 39730
rect 42478 39678 42530 39730
rect 42702 39678 42754 39730
rect 44382 39678 44434 39730
rect 45278 39678 45330 39730
rect 1822 39566 1874 39618
rect 5630 39566 5682 39618
rect 11118 39566 11170 39618
rect 11678 39566 11730 39618
rect 12350 39566 12402 39618
rect 13022 39566 13074 39618
rect 13806 39566 13858 39618
rect 14142 39566 14194 39618
rect 17950 39566 18002 39618
rect 20750 39566 20802 39618
rect 21982 39566 22034 39618
rect 22318 39566 22370 39618
rect 22878 39566 22930 39618
rect 24110 39566 24162 39618
rect 24446 39566 24498 39618
rect 26126 39566 26178 39618
rect 29486 39566 29538 39618
rect 30158 39566 30210 39618
rect 31166 39566 31218 39618
rect 31838 39566 31890 39618
rect 32510 39566 32562 39618
rect 33182 39566 33234 39618
rect 33742 39566 33794 39618
rect 34414 39566 34466 39618
rect 35534 39566 35586 39618
rect 36430 39566 36482 39618
rect 36990 39566 37042 39618
rect 37214 39566 37266 39618
rect 37438 39566 37490 39618
rect 41134 39566 41186 39618
rect 41582 39566 41634 39618
rect 41694 39566 41746 39618
rect 42030 39566 42082 39618
rect 42254 39566 42306 39618
rect 43038 39566 43090 39618
rect 43374 39566 43426 39618
rect 43822 39566 43874 39618
rect 44046 39566 44098 39618
rect 48078 39566 48130 39618
rect 6414 39454 6466 39506
rect 9998 39454 10050 39506
rect 10334 39454 10386 39506
rect 11230 39454 11282 39506
rect 11790 39454 11842 39506
rect 12574 39454 12626 39506
rect 13470 39454 13522 39506
rect 14814 39454 14866 39506
rect 18846 39454 18898 39506
rect 20526 39454 20578 39506
rect 21534 39454 21586 39506
rect 22206 39454 22258 39506
rect 23214 39454 23266 39506
rect 24894 39454 24946 39506
rect 26798 39454 26850 39506
rect 28142 39454 28194 39506
rect 32174 39454 32226 39506
rect 32734 39454 32786 39506
rect 33630 39454 33682 39506
rect 40350 39454 40402 39506
rect 44830 39454 44882 39506
rect 47406 39454 47458 39506
rect 5070 39342 5122 39394
rect 8878 39342 8930 39394
rect 9214 39342 9266 39394
rect 10894 39342 10946 39394
rect 11454 39342 11506 39394
rect 12798 39342 12850 39394
rect 13582 39342 13634 39394
rect 17390 39342 17442 39394
rect 25006 39342 25058 39394
rect 30606 39342 30658 39394
rect 37662 39342 37714 39394
rect 42478 39342 42530 39394
rect 43262 39342 43314 39394
rect 43822 39342 43874 39394
rect 44942 39342 44994 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 4286 39006 4338 39058
rect 4622 39006 4674 39058
rect 5966 39006 6018 39058
rect 8094 39006 8146 39058
rect 9886 39006 9938 39058
rect 11118 39006 11170 39058
rect 11342 39006 11394 39058
rect 14926 39006 14978 39058
rect 15934 39006 15986 39058
rect 17838 39006 17890 39058
rect 17950 39006 18002 39058
rect 20974 39006 21026 39058
rect 22654 39006 22706 39058
rect 23214 39006 23266 39058
rect 28590 39006 28642 39058
rect 29038 39006 29090 39058
rect 32062 39006 32114 39058
rect 35198 39006 35250 39058
rect 36766 39006 36818 39058
rect 40014 39006 40066 39058
rect 41022 39006 41074 39058
rect 42030 39006 42082 39058
rect 42366 39006 42418 39058
rect 44270 39006 44322 39058
rect 44830 39006 44882 39058
rect 2494 38894 2546 38946
rect 4846 38894 4898 38946
rect 8318 38894 8370 38946
rect 9662 38894 9714 38946
rect 10558 38894 10610 38946
rect 11006 38894 11058 38946
rect 13918 38894 13970 38946
rect 14366 38894 14418 38946
rect 15374 38894 15426 38946
rect 15598 38894 15650 38946
rect 19854 38894 19906 38946
rect 20302 38894 20354 38946
rect 21310 38894 21362 38946
rect 21758 38894 21810 38946
rect 21870 38894 21922 38946
rect 22318 38894 22370 38946
rect 22430 38894 22482 38946
rect 22990 38894 23042 38946
rect 24558 38894 24610 38946
rect 25454 38894 25506 38946
rect 27694 38894 27746 38946
rect 29150 38894 29202 38946
rect 31278 38894 31330 38946
rect 34078 38894 34130 38946
rect 37550 38894 37602 38946
rect 40910 38894 40962 38946
rect 42478 38894 42530 38946
rect 44494 38894 44546 38946
rect 3166 38782 3218 38834
rect 3838 38782 3890 38834
rect 4174 38782 4226 38834
rect 4398 38782 4450 38834
rect 4958 38782 5010 38834
rect 5630 38782 5682 38834
rect 5854 38782 5906 38834
rect 6190 38782 6242 38834
rect 6974 38782 7026 38834
rect 7646 38782 7698 38834
rect 8206 38782 8258 38834
rect 9550 38782 9602 38834
rect 10334 38782 10386 38834
rect 10670 38782 10722 38834
rect 13022 38782 13074 38834
rect 14254 38782 14306 38834
rect 14590 38782 14642 38834
rect 16046 38782 16098 38834
rect 16382 38782 16434 38834
rect 17278 38782 17330 38834
rect 17726 38782 17778 38834
rect 20750 38782 20802 38834
rect 20974 38782 21026 38834
rect 22878 38782 22930 38834
rect 23662 38782 23714 38834
rect 26014 38782 26066 38834
rect 26238 38782 26290 38834
rect 27246 38782 27298 38834
rect 27470 38782 27522 38834
rect 27806 38782 27858 38834
rect 29710 38782 29762 38834
rect 30046 38782 30098 38834
rect 33406 38782 33458 38834
rect 34750 38782 34802 38834
rect 34974 38782 35026 38834
rect 36542 38782 36594 38834
rect 38110 38782 38162 38834
rect 38782 38782 38834 38834
rect 43038 38782 43090 38834
rect 43150 38782 43202 38834
rect 43262 38782 43314 38834
rect 43710 38782 43762 38834
rect 44158 38782 44210 38834
rect 48078 38782 48130 38834
rect 3390 38670 3442 38722
rect 6414 38670 6466 38722
rect 6862 38670 6914 38722
rect 8878 38670 8930 38722
rect 12014 38670 12066 38722
rect 12574 38670 12626 38722
rect 13134 38670 13186 38722
rect 15262 38670 15314 38722
rect 18398 38670 18450 38722
rect 18958 38670 19010 38722
rect 19406 38670 19458 38722
rect 20414 38670 20466 38722
rect 21646 38670 21698 38722
rect 24110 38670 24162 38722
rect 25566 38670 25618 38722
rect 27022 38670 27074 38722
rect 28926 38670 28978 38722
rect 32510 38670 32562 38722
rect 33182 38670 33234 38722
rect 34862 38670 34914 38722
rect 35758 38670 35810 38722
rect 36094 38670 36146 38722
rect 36878 38670 36930 38722
rect 39454 38670 39506 38722
rect 39790 38670 39842 38722
rect 40126 38670 40178 38722
rect 41582 38670 41634 38722
rect 43822 38670 43874 38722
rect 47406 38670 47458 38722
rect 16382 38558 16434 38610
rect 16718 38558 16770 38610
rect 18510 38558 18562 38610
rect 19406 38558 19458 38610
rect 20078 38558 20130 38610
rect 45278 38614 45330 38666
rect 25230 38558 25282 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 3614 38222 3666 38274
rect 5630 38222 5682 38274
rect 6190 38222 6242 38274
rect 31390 38222 31442 38274
rect 3166 38110 3218 38162
rect 5070 38110 5122 38162
rect 8318 38110 8370 38162
rect 15038 38110 15090 38162
rect 15598 38110 15650 38162
rect 16270 38110 16322 38162
rect 20302 38110 20354 38162
rect 23998 38110 24050 38162
rect 25678 38110 25730 38162
rect 29598 38110 29650 38162
rect 34862 38110 34914 38162
rect 35870 38110 35922 38162
rect 37102 38110 37154 38162
rect 44046 38110 44098 38162
rect 44942 38110 44994 38162
rect 3726 37998 3778 38050
rect 4174 37998 4226 38050
rect 4734 37998 4786 38050
rect 6414 37998 6466 38050
rect 6638 37998 6690 38050
rect 7086 37998 7138 38050
rect 10334 37998 10386 38050
rect 11230 37998 11282 38050
rect 12462 37998 12514 38050
rect 13582 37998 13634 38050
rect 13918 37998 13970 38050
rect 15374 37998 15426 38050
rect 16158 37998 16210 38050
rect 17502 37998 17554 38050
rect 21310 37998 21362 38050
rect 23550 37998 23602 38050
rect 23886 37998 23938 38050
rect 24334 37998 24386 38050
rect 28478 37998 28530 38050
rect 30046 37998 30098 38050
rect 30270 37998 30322 38050
rect 31950 37998 32002 38050
rect 41134 37998 41186 38050
rect 47630 37998 47682 38050
rect 8654 37886 8706 37938
rect 9662 37886 9714 37938
rect 10446 37886 10498 37938
rect 10894 37886 10946 37938
rect 18174 37886 18226 37938
rect 21534 37886 21586 37938
rect 21646 37886 21698 37938
rect 22318 37886 22370 37938
rect 24670 37886 24722 37938
rect 26014 37886 26066 37938
rect 27582 37886 27634 37938
rect 27806 37886 27858 37938
rect 28142 37886 28194 37938
rect 29262 37886 29314 37938
rect 30942 37886 30994 37938
rect 31502 37886 31554 37938
rect 32734 37886 32786 37938
rect 36206 37886 36258 37938
rect 36990 37886 37042 37938
rect 37774 37886 37826 37938
rect 40686 37886 40738 37938
rect 40798 37886 40850 37938
rect 41918 37886 41970 37938
rect 45166 37886 45218 37938
rect 46846 37886 46898 37938
rect 2270 37774 2322 37826
rect 3614 37774 3666 37826
rect 4062 37774 4114 37826
rect 4286 37774 4338 37826
rect 5742 37774 5794 37826
rect 6526 37774 6578 37826
rect 7646 37774 7698 37826
rect 8990 37774 9042 37826
rect 9326 37774 9378 37826
rect 10670 37774 10722 37826
rect 11006 37774 11058 37826
rect 11566 37774 11618 37826
rect 11902 37774 11954 37826
rect 12014 37774 12066 37826
rect 12126 37774 12178 37826
rect 13022 37774 13074 37826
rect 20750 37774 20802 37826
rect 22654 37774 22706 37826
rect 25230 37774 25282 37826
rect 28254 37774 28306 37826
rect 29486 37774 29538 37826
rect 31390 37774 31442 37826
rect 35310 37774 35362 37826
rect 36318 37774 36370 37826
rect 36542 37774 36594 37826
rect 37214 37774 37266 37826
rect 37662 37774 37714 37826
rect 38222 37774 38274 37826
rect 38782 37774 38834 37826
rect 39118 37774 39170 37826
rect 39902 37774 39954 37826
rect 40350 37774 40402 37826
rect 46734 37774 46786 37826
rect 48190 37774 48242 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 5406 37438 5458 37490
rect 6638 37438 6690 37490
rect 7646 37438 7698 37490
rect 21646 37438 21698 37490
rect 34414 37438 34466 37490
rect 41022 37438 41074 37490
rect 43486 37438 43538 37490
rect 6862 37326 6914 37378
rect 10670 37326 10722 37378
rect 14702 37326 14754 37378
rect 16494 37326 16546 37378
rect 19182 37326 19234 37378
rect 20302 37326 20354 37378
rect 21534 37326 21586 37378
rect 23774 37326 23826 37378
rect 29262 37326 29314 37378
rect 34302 37326 34354 37378
rect 34862 37326 34914 37378
rect 35198 37326 35250 37378
rect 36990 37326 37042 37378
rect 41134 37326 41186 37378
rect 43038 37326 43090 37378
rect 47070 37326 47122 37378
rect 1822 37214 1874 37266
rect 4846 37214 4898 37266
rect 5294 37214 5346 37266
rect 5518 37214 5570 37266
rect 5742 37214 5794 37266
rect 6190 37214 6242 37266
rect 6302 37214 6354 37266
rect 6974 37214 7026 37266
rect 8430 37214 8482 37266
rect 8766 37214 8818 37266
rect 9774 37214 9826 37266
rect 10222 37214 10274 37266
rect 11006 37214 11058 37266
rect 15934 37214 15986 37266
rect 17502 37214 17554 37266
rect 18734 37214 18786 37266
rect 19070 37214 19122 37266
rect 19406 37214 19458 37266
rect 23214 37214 23266 37266
rect 30046 37214 30098 37266
rect 30830 37214 30882 37266
rect 31054 37214 31106 37266
rect 31726 37214 31778 37266
rect 32510 37214 32562 37266
rect 33518 37214 33570 37266
rect 34638 37214 34690 37266
rect 35422 37214 35474 37266
rect 35870 37214 35922 37266
rect 36766 37214 36818 37266
rect 37102 37214 37154 37266
rect 37438 37214 37490 37266
rect 41694 37214 41746 37266
rect 41918 37214 41970 37266
rect 42702 37214 42754 37266
rect 44494 37214 44546 37266
rect 47742 37214 47794 37266
rect 2494 37102 2546 37154
rect 4622 37102 4674 37154
rect 5966 37102 6018 37154
rect 8990 37102 9042 37154
rect 11790 37102 11842 37154
rect 13918 37102 13970 37154
rect 14366 37102 14418 37154
rect 18398 37102 18450 37154
rect 19742 37102 19794 37154
rect 22318 37102 22370 37154
rect 22990 37102 23042 37154
rect 26350 37102 26402 37154
rect 26798 37102 26850 37154
rect 27134 37102 27186 37154
rect 31838 37102 31890 37154
rect 33966 37102 34018 37154
rect 38222 37102 38274 37154
rect 40350 37102 40402 37154
rect 43934 37102 43986 37154
rect 44942 37102 44994 37154
rect 17390 36990 17442 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 5854 36654 5906 36706
rect 8430 36654 8482 36706
rect 9998 36654 10050 36706
rect 10446 36654 10498 36706
rect 14702 36654 14754 36706
rect 15038 36654 15090 36706
rect 21870 36654 21922 36706
rect 27582 36654 27634 36706
rect 37998 36654 38050 36706
rect 46846 36654 46898 36706
rect 4510 36542 4562 36594
rect 7310 36542 7362 36594
rect 8766 36542 8818 36594
rect 10894 36542 10946 36594
rect 15374 36542 15426 36594
rect 17502 36542 17554 36594
rect 21310 36542 21362 36594
rect 23774 36542 23826 36594
rect 31054 36542 31106 36594
rect 35086 36542 35138 36594
rect 36318 36542 36370 36594
rect 38670 36542 38722 36594
rect 40798 36542 40850 36594
rect 43150 36542 43202 36594
rect 45838 36542 45890 36594
rect 47630 36542 47682 36594
rect 4062 36430 4114 36482
rect 4398 36430 4450 36482
rect 6526 36430 6578 36482
rect 7198 36430 7250 36482
rect 8206 36430 8258 36482
rect 9214 36430 9266 36482
rect 9438 36430 9490 36482
rect 10558 36430 10610 36482
rect 11342 36430 11394 36482
rect 11902 36430 11954 36482
rect 12350 36430 12402 36482
rect 12462 36430 12514 36482
rect 13918 36430 13970 36482
rect 14142 36430 14194 36482
rect 15038 36430 15090 36482
rect 18286 36430 18338 36482
rect 18734 36430 18786 36482
rect 18846 36430 18898 36482
rect 19966 36430 20018 36482
rect 20414 36430 20466 36482
rect 20526 36430 20578 36482
rect 21534 36430 21586 36482
rect 22206 36430 22258 36482
rect 22430 36430 22482 36482
rect 22766 36430 22818 36482
rect 23102 36430 23154 36482
rect 23998 36430 24050 36482
rect 26574 36430 26626 36482
rect 26798 36430 26850 36482
rect 27358 36430 27410 36482
rect 30382 36430 30434 36482
rect 30942 36430 30994 36482
rect 32958 36430 33010 36482
rect 33630 36430 33682 36482
rect 34190 36430 34242 36482
rect 36206 36430 36258 36482
rect 39230 36430 39282 36482
rect 39342 36430 39394 36482
rect 39678 36430 39730 36482
rect 41582 36430 41634 36482
rect 42142 36430 42194 36482
rect 42254 36430 42306 36482
rect 44830 36430 44882 36482
rect 45502 36430 45554 36482
rect 46062 36430 46114 36482
rect 46622 36430 46674 36482
rect 47406 36430 47458 36482
rect 4958 36318 5010 36370
rect 5070 36318 5122 36370
rect 5854 36318 5906 36370
rect 5966 36318 6018 36370
rect 6302 36318 6354 36370
rect 6862 36318 6914 36370
rect 7422 36318 7474 36370
rect 9550 36318 9602 36370
rect 13582 36318 13634 36370
rect 19182 36318 19234 36370
rect 1822 36206 1874 36258
rect 2270 36206 2322 36258
rect 2718 36206 2770 36258
rect 3166 36206 3218 36258
rect 4734 36206 4786 36258
rect 6414 36206 6466 36258
rect 7646 36206 7698 36258
rect 12126 36206 12178 36258
rect 13694 36206 13746 36258
rect 14254 36206 14306 36258
rect 14478 36206 14530 36258
rect 19070 36206 19122 36258
rect 19406 36206 19458 36258
rect 19630 36262 19682 36314
rect 19742 36318 19794 36370
rect 23214 36318 23266 36370
rect 27022 36318 27074 36370
rect 29150 36318 29202 36370
rect 31054 36318 31106 36370
rect 31838 36318 31890 36370
rect 32398 36318 32450 36370
rect 34302 36318 34354 36370
rect 34638 36318 34690 36370
rect 35758 36318 35810 36370
rect 36990 36318 37042 36370
rect 38558 36318 38610 36370
rect 42366 36318 42418 36370
rect 42702 36318 42754 36370
rect 43486 36318 43538 36370
rect 20638 36206 20690 36258
rect 24670 36206 24722 36258
rect 25118 36206 25170 36258
rect 27918 36206 27970 36258
rect 28590 36206 28642 36258
rect 29262 36206 29314 36258
rect 29374 36206 29426 36258
rect 29598 36206 29650 36258
rect 31950 36206 32002 36258
rect 32174 36206 32226 36258
rect 35982 36206 36034 36258
rect 36318 36206 36370 36258
rect 38782 36206 38834 36258
rect 39566 36206 39618 36258
rect 40126 36206 40178 36258
rect 41134 36206 41186 36258
rect 41246 36206 41298 36258
rect 41358 36206 41410 36258
rect 41470 36206 41522 36258
rect 42478 36206 42530 36258
rect 43598 36206 43650 36258
rect 43934 36206 43986 36258
rect 44270 36206 44322 36258
rect 45166 36206 45218 36258
rect 45726 36206 45778 36258
rect 45950 36206 46002 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 5742 35870 5794 35922
rect 7534 35870 7586 35922
rect 7646 35870 7698 35922
rect 8542 35870 8594 35922
rect 9774 35870 9826 35922
rect 10222 35870 10274 35922
rect 12686 35870 12738 35922
rect 13694 35870 13746 35922
rect 15150 35870 15202 35922
rect 23662 35870 23714 35922
rect 28142 35870 28194 35922
rect 34974 35870 35026 35922
rect 39342 35870 39394 35922
rect 43150 35870 43202 35922
rect 44158 35870 44210 35922
rect 44830 35870 44882 35922
rect 2494 35758 2546 35810
rect 7086 35758 7138 35810
rect 7422 35758 7474 35810
rect 9998 35758 10050 35810
rect 11790 35758 11842 35810
rect 14030 35758 14082 35810
rect 15710 35758 15762 35810
rect 16494 35758 16546 35810
rect 16830 35758 16882 35810
rect 18174 35758 18226 35810
rect 23326 35758 23378 35810
rect 26238 35758 26290 35810
rect 27694 35758 27746 35810
rect 29150 35758 29202 35810
rect 30046 35758 30098 35810
rect 30158 35758 30210 35810
rect 32286 35758 32338 35810
rect 33518 35758 33570 35810
rect 38894 35758 38946 35810
rect 39902 35758 39954 35810
rect 42142 35758 42194 35810
rect 44718 35758 44770 35810
rect 46062 35758 46114 35810
rect 1710 35646 1762 35698
rect 6190 35646 6242 35698
rect 6638 35646 6690 35698
rect 7982 35646 8034 35698
rect 8878 35646 8930 35698
rect 9886 35646 9938 35698
rect 10670 35646 10722 35698
rect 11230 35646 11282 35698
rect 12126 35646 12178 35698
rect 12574 35646 12626 35698
rect 12798 35646 12850 35698
rect 13134 35646 13186 35698
rect 14366 35646 14418 35698
rect 16046 35646 16098 35698
rect 17390 35646 17442 35698
rect 20750 35646 20802 35698
rect 21086 35646 21138 35698
rect 22878 35646 22930 35698
rect 23214 35646 23266 35698
rect 23998 35646 24050 35698
rect 26462 35646 26514 35698
rect 27022 35646 27074 35698
rect 27470 35646 27522 35698
rect 28030 35646 28082 35698
rect 28590 35646 28642 35698
rect 30382 35646 30434 35698
rect 31166 35646 31218 35698
rect 31950 35646 32002 35698
rect 34638 35646 34690 35698
rect 38446 35646 38498 35698
rect 39118 35646 39170 35698
rect 41470 35646 41522 35698
rect 41694 35646 41746 35698
rect 41806 35646 41858 35698
rect 42478 35646 42530 35698
rect 43598 35646 43650 35698
rect 45390 35646 45442 35698
rect 4622 35534 4674 35586
rect 5294 35534 5346 35586
rect 11902 35534 11954 35586
rect 15262 35534 15314 35586
rect 20302 35534 20354 35586
rect 20638 35534 20690 35586
rect 24446 35534 24498 35586
rect 25342 35534 25394 35586
rect 25790 35534 25842 35586
rect 26798 35534 26850 35586
rect 27246 35534 27298 35586
rect 29710 35534 29762 35586
rect 30830 35534 30882 35586
rect 31614 35534 31666 35586
rect 33182 35534 33234 35586
rect 35646 35534 35698 35586
rect 37774 35534 37826 35586
rect 39006 35534 39058 35586
rect 40350 35534 40402 35586
rect 41246 35534 41298 35586
rect 42590 35534 42642 35586
rect 42702 35534 42754 35586
rect 48190 35534 48242 35586
rect 11566 35422 11618 35474
rect 13358 35422 13410 35474
rect 15374 35422 15426 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 13358 35086 13410 35138
rect 14814 35086 14866 35138
rect 19518 35086 19570 35138
rect 28478 35086 28530 35138
rect 29710 35086 29762 35138
rect 30494 35086 30546 35138
rect 36990 35086 37042 35138
rect 37326 35086 37378 35138
rect 3726 34974 3778 35026
rect 5742 34974 5794 35026
rect 9886 34974 9938 35026
rect 10894 34974 10946 35026
rect 14254 34974 14306 35026
rect 15150 34974 15202 35026
rect 15934 34974 15986 35026
rect 17838 34974 17890 35026
rect 18734 34974 18786 35026
rect 21310 34974 21362 35026
rect 24334 34974 24386 35026
rect 26462 34974 26514 35026
rect 30942 34974 30994 35026
rect 35982 34974 36034 35026
rect 38670 34974 38722 35026
rect 40798 34974 40850 35026
rect 41246 34974 41298 35026
rect 42478 34974 42530 35026
rect 44158 34974 44210 35026
rect 48190 34974 48242 35026
rect 2606 34862 2658 34914
rect 5630 34862 5682 34914
rect 6190 34862 6242 34914
rect 6414 34862 6466 34914
rect 6750 34862 6802 34914
rect 7646 34862 7698 34914
rect 9662 34862 9714 34914
rect 11678 34862 11730 34914
rect 13806 34862 13858 34914
rect 14030 34862 14082 34914
rect 16270 34862 16322 34914
rect 16606 34862 16658 34914
rect 18174 34862 18226 34914
rect 18622 34862 18674 34914
rect 18846 34862 18898 34914
rect 2942 34750 2994 34802
rect 3166 34750 3218 34802
rect 4174 34750 4226 34802
rect 7310 34750 7362 34802
rect 7870 34750 7922 34802
rect 8766 34750 8818 34802
rect 10334 34750 10386 34802
rect 11006 34750 11058 34802
rect 19406 34806 19458 34858
rect 22318 34862 22370 34914
rect 22878 34862 22930 34914
rect 23550 34862 23602 34914
rect 27358 34862 27410 34914
rect 27582 34862 27634 34914
rect 28254 34862 28306 34914
rect 29150 34862 29202 34914
rect 29374 34862 29426 34914
rect 30382 34862 30434 34914
rect 31390 34862 31442 34914
rect 32398 34862 32450 34914
rect 32734 34862 32786 34914
rect 34302 34862 34354 34914
rect 35198 34862 35250 34914
rect 35310 34862 35362 34914
rect 35870 34862 35922 34914
rect 36206 34862 36258 34914
rect 37998 34862 38050 34914
rect 41806 34862 41858 34914
rect 45278 34862 45330 34914
rect 11230 34750 11282 34802
rect 11902 34750 11954 34802
rect 12574 34750 12626 34802
rect 15374 34750 15426 34802
rect 15710 34750 15762 34802
rect 19966 34750 20018 34802
rect 20078 34750 20130 34802
rect 20526 34750 20578 34802
rect 21422 34750 21474 34802
rect 21646 34750 21698 34802
rect 21982 34750 22034 34802
rect 22654 34750 22706 34802
rect 33406 34750 33458 34802
rect 34414 34750 34466 34802
rect 34974 34750 35026 34802
rect 36318 34750 36370 34802
rect 42926 34750 42978 34802
rect 44046 34750 44098 34802
rect 44270 34750 44322 34802
rect 46062 34750 46114 34802
rect 1822 34638 1874 34690
rect 2382 34638 2434 34690
rect 2718 34638 2770 34690
rect 4622 34638 4674 34690
rect 5182 34638 5234 34690
rect 5854 34638 5906 34690
rect 6638 34638 6690 34690
rect 7422 34638 7474 34690
rect 8206 34638 8258 34690
rect 8878 34638 8930 34690
rect 9102 34638 9154 34690
rect 12238 34638 12290 34690
rect 17390 34638 17442 34690
rect 19518 34638 19570 34690
rect 20302 34638 20354 34690
rect 20638 34638 20690 34690
rect 20862 34638 20914 34690
rect 32846 34638 32898 34690
rect 32958 34638 33010 34690
rect 33854 34638 33906 34690
rect 35422 34638 35474 34690
rect 37214 34638 37266 34690
rect 41246 34638 41298 34690
rect 41358 34638 41410 34690
rect 41582 34638 41634 34690
rect 42590 34638 42642 34690
rect 43262 34638 43314 34690
rect 44942 34638 44994 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 6862 34302 6914 34354
rect 12350 34302 12402 34354
rect 19182 34302 19234 34354
rect 19294 34302 19346 34354
rect 42030 34302 42082 34354
rect 45726 34302 45778 34354
rect 45838 34302 45890 34354
rect 47854 34302 47906 34354
rect 2494 34190 2546 34242
rect 6526 34190 6578 34242
rect 7086 34190 7138 34242
rect 7198 34190 7250 34242
rect 7870 34190 7922 34242
rect 9998 34190 10050 34242
rect 11678 34190 11730 34242
rect 15710 34190 15762 34242
rect 17726 34190 17778 34242
rect 20974 34190 21026 34242
rect 23550 34190 23602 34242
rect 23662 34190 23714 34242
rect 23886 34190 23938 34242
rect 28814 34190 28866 34242
rect 30830 34190 30882 34242
rect 32174 34190 32226 34242
rect 37326 34190 37378 34242
rect 38670 34190 38722 34242
rect 41022 34190 41074 34242
rect 44382 34190 44434 34242
rect 1710 34078 1762 34130
rect 4958 34078 5010 34130
rect 5182 34078 5234 34130
rect 5630 34078 5682 34130
rect 6302 34078 6354 34130
rect 6638 34078 6690 34130
rect 7758 34078 7810 34130
rect 8094 34078 8146 34130
rect 8878 34078 8930 34130
rect 10334 34078 10386 34130
rect 11118 34078 11170 34130
rect 13246 34078 13298 34130
rect 13582 34078 13634 34130
rect 13918 34078 13970 34130
rect 14366 34078 14418 34130
rect 14814 34078 14866 34130
rect 15150 34078 15202 34130
rect 16718 34078 16770 34130
rect 17390 34078 17442 34130
rect 17838 34078 17890 34130
rect 18286 34078 18338 34130
rect 19406 34078 19458 34130
rect 19742 34078 19794 34130
rect 20190 34078 20242 34130
rect 24110 34078 24162 34130
rect 24558 34078 24610 34130
rect 25230 34078 25282 34130
rect 25342 34078 25394 34130
rect 25454 34078 25506 34130
rect 25790 34078 25842 34130
rect 26574 34078 26626 34130
rect 27470 34078 27522 34130
rect 27918 34078 27970 34130
rect 28142 34078 28194 34130
rect 29598 34078 29650 34130
rect 31278 34078 31330 34130
rect 31502 34078 31554 34130
rect 32958 34078 33010 34130
rect 33294 34078 33346 34130
rect 33518 34078 33570 34130
rect 34190 34078 34242 34130
rect 38446 34078 38498 34130
rect 39678 34078 39730 34130
rect 40014 34078 40066 34130
rect 40238 34078 40290 34130
rect 41470 34078 41522 34130
rect 45166 34078 45218 34130
rect 45950 34078 46002 34130
rect 46286 34078 46338 34130
rect 47182 34078 47234 34130
rect 4622 33966 4674 34018
rect 8318 33966 8370 34018
rect 10110 33966 10162 34018
rect 11006 33966 11058 34018
rect 12686 33966 12738 34018
rect 16158 33966 16210 34018
rect 17502 33966 17554 34018
rect 18734 33966 18786 34018
rect 23102 33966 23154 34018
rect 26798 33966 26850 34018
rect 29710 33966 29762 34018
rect 33182 33966 33234 34018
rect 35534 33966 35586 34018
rect 37102 33966 37154 34018
rect 40126 33966 40178 34018
rect 42254 33966 42306 34018
rect 46622 33966 46674 34018
rect 9774 33854 9826 33906
rect 40910 33854 40962 33906
rect 41246 33854 41298 33906
rect 42030 33854 42082 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 4510 33518 4562 33570
rect 6078 33518 6130 33570
rect 7422 33518 7474 33570
rect 12910 33518 12962 33570
rect 28254 33518 28306 33570
rect 31054 33518 31106 33570
rect 36094 33518 36146 33570
rect 46846 33518 46898 33570
rect 3054 33406 3106 33458
rect 4398 33406 4450 33458
rect 7982 33406 8034 33458
rect 10110 33406 10162 33458
rect 14030 33406 14082 33458
rect 15486 33406 15538 33458
rect 17614 33406 17666 33458
rect 18958 33406 19010 33458
rect 27358 33406 27410 33458
rect 27694 33406 27746 33458
rect 29710 33406 29762 33458
rect 30830 33406 30882 33458
rect 32734 33406 32786 33458
rect 34862 33406 34914 33458
rect 35422 33406 35474 33458
rect 37326 33406 37378 33458
rect 40126 33406 40178 33458
rect 42254 33406 42306 33458
rect 44942 33406 44994 33458
rect 3614 33294 3666 33346
rect 7422 33294 7474 33346
rect 10894 33294 10946 33346
rect 11678 33294 11730 33346
rect 12014 33294 12066 33346
rect 12910 33294 12962 33346
rect 14254 33294 14306 33346
rect 18398 33294 18450 33346
rect 19294 33294 19346 33346
rect 19742 33294 19794 33346
rect 22094 33294 22146 33346
rect 22878 33294 22930 33346
rect 24894 33294 24946 33346
rect 25678 33294 25730 33346
rect 27918 33294 27970 33346
rect 29374 33294 29426 33346
rect 30158 33294 30210 33346
rect 30942 33294 30994 33346
rect 32062 33294 32114 33346
rect 36094 33294 36146 33346
rect 37662 33294 37714 33346
rect 38334 33294 38386 33346
rect 38782 33294 38834 33346
rect 39342 33294 39394 33346
rect 43710 33294 43762 33346
rect 45838 33294 45890 33346
rect 47070 33294 47122 33346
rect 47630 33294 47682 33346
rect 47854 33294 47906 33346
rect 1710 33182 1762 33234
rect 1822 33182 1874 33234
rect 2270 33182 2322 33234
rect 3166 33182 3218 33234
rect 4062 33182 4114 33234
rect 5070 33182 5122 33234
rect 2046 33070 2098 33122
rect 2382 33070 2434 33122
rect 2606 33070 2658 33122
rect 2942 33070 2994 33122
rect 3726 33070 3778 33122
rect 3950 33070 4002 33122
rect 4734 33070 4786 33122
rect 4958 33070 5010 33122
rect 5854 33070 5906 33122
rect 5966 33070 6018 33122
rect 6302 33070 6354 33122
rect 6526 33070 6578 33122
rect 6638 33126 6690 33178
rect 7086 33182 7138 33234
rect 12574 33182 12626 33234
rect 14926 33182 14978 33234
rect 23102 33182 23154 33234
rect 24446 33182 24498 33234
rect 26350 33182 26402 33234
rect 29150 33182 29202 33234
rect 35758 33182 35810 33234
rect 36990 33182 37042 33234
rect 37998 33182 38050 33234
rect 43374 33182 43426 33234
rect 43934 33182 43986 33234
rect 44830 33182 44882 33234
rect 46174 33182 46226 33234
rect 47406 33182 47458 33234
rect 47518 33182 47570 33234
rect 11454 33070 11506 33122
rect 11566 33070 11618 33122
rect 13694 33070 13746 33122
rect 20414 33070 20466 33122
rect 20750 33070 20802 33122
rect 21646 33070 21698 33122
rect 26798 33070 26850 33122
rect 37214 33070 37266 33122
rect 37438 33070 37490 33122
rect 38110 33070 38162 33122
rect 38446 33070 38498 33122
rect 38670 33070 38722 33122
rect 43038 33070 43090 33122
rect 43822 33070 43874 33122
rect 45390 33070 45442 33122
rect 46062 33070 46114 33122
rect 46510 33070 46562 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 11902 32734 11954 32786
rect 15374 32734 15426 32786
rect 23214 32734 23266 32786
rect 24110 32734 24162 32786
rect 31502 32734 31554 32786
rect 32510 32734 32562 32786
rect 34974 32734 35026 32786
rect 36318 32734 36370 32786
rect 3054 32622 3106 32674
rect 3838 32622 3890 32674
rect 8206 32622 8258 32674
rect 10110 32622 10162 32674
rect 23438 32622 23490 32674
rect 24446 32622 24498 32674
rect 24558 32622 24610 32674
rect 25230 32622 25282 32674
rect 27022 32622 27074 32674
rect 29598 32622 29650 32674
rect 33518 32622 33570 32674
rect 36430 32622 36482 32674
rect 40910 32622 40962 32674
rect 41470 32622 41522 32674
rect 46062 32622 46114 32674
rect 2046 32510 2098 32562
rect 2270 32510 2322 32562
rect 2494 32510 2546 32562
rect 2830 32510 2882 32562
rect 3390 32510 3442 32562
rect 3614 32510 3666 32562
rect 3950 32510 4002 32562
rect 4958 32510 5010 32562
rect 5742 32510 5794 32562
rect 8990 32510 9042 32562
rect 11342 32510 11394 32562
rect 14478 32510 14530 32562
rect 15262 32510 15314 32562
rect 15598 32510 15650 32562
rect 16382 32510 16434 32562
rect 16830 32510 16882 32562
rect 19742 32510 19794 32562
rect 21310 32510 21362 32562
rect 22430 32510 22482 32562
rect 22654 32510 22706 32562
rect 23774 32510 23826 32562
rect 25678 32510 25730 32562
rect 27246 32510 27298 32562
rect 28702 32510 28754 32562
rect 30606 32510 30658 32562
rect 34862 32510 34914 32562
rect 37102 32510 37154 32562
rect 41134 32510 41186 32562
rect 44718 32510 44770 32562
rect 45390 32510 45442 32562
rect 2382 32398 2434 32450
rect 2942 32398 2994 32450
rect 5070 32398 5122 32450
rect 5630 32398 5682 32450
rect 9998 32398 10050 32450
rect 12574 32398 12626 32450
rect 16046 32398 16098 32450
rect 19182 32398 19234 32450
rect 20638 32398 20690 32450
rect 20862 32398 20914 32450
rect 21646 32398 21698 32450
rect 23102 32398 23154 32450
rect 25566 32398 25618 32450
rect 27806 32398 27858 32450
rect 29262 32398 29314 32450
rect 30718 32398 30770 32450
rect 33182 32398 33234 32450
rect 35982 32398 36034 32450
rect 38222 32398 38274 32450
rect 40238 32398 40290 32450
rect 6078 32342 6130 32394
rect 41358 32398 41410 32450
rect 41918 32398 41970 32450
rect 44046 32398 44098 32450
rect 48190 32398 48242 32450
rect 24558 32286 24610 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 3054 31950 3106 32002
rect 8542 31950 8594 32002
rect 8878 31950 8930 32002
rect 11790 31950 11842 32002
rect 12238 31950 12290 32002
rect 22094 31950 22146 32002
rect 43934 31950 43986 32002
rect 45726 31950 45778 32002
rect 8318 31838 8370 31890
rect 9774 31838 9826 31890
rect 10222 31838 10274 31890
rect 13806 31838 13858 31890
rect 16158 31838 16210 31890
rect 20302 31838 20354 31890
rect 23102 31838 23154 31890
rect 23998 31838 24050 31890
rect 32622 31838 32674 31890
rect 33518 31838 33570 31890
rect 37326 31838 37378 31890
rect 38110 31838 38162 31890
rect 39342 31838 39394 31890
rect 41470 31838 41522 31890
rect 44158 31838 44210 31890
rect 44382 31838 44434 31890
rect 1934 31726 1986 31778
rect 2830 31726 2882 31778
rect 6974 31726 7026 31778
rect 9438 31726 9490 31778
rect 10334 31726 10386 31778
rect 12462 31726 12514 31778
rect 13694 31726 13746 31778
rect 14590 31726 14642 31778
rect 15822 31726 15874 31778
rect 16606 31726 16658 31778
rect 17502 31726 17554 31778
rect 21198 31726 21250 31778
rect 22766 31726 22818 31778
rect 23326 31726 23378 31778
rect 24110 31726 24162 31778
rect 25454 31726 25506 31778
rect 25790 31726 25842 31778
rect 26462 31726 26514 31778
rect 27134 31726 27186 31778
rect 28030 31726 28082 31778
rect 30494 31726 30546 31778
rect 31614 31726 31666 31778
rect 36430 31726 36482 31778
rect 37998 31726 38050 31778
rect 38558 31726 38610 31778
rect 42254 31726 42306 31778
rect 43598 31726 43650 31778
rect 43934 31726 43986 31778
rect 45950 31726 46002 31778
rect 46174 31726 46226 31778
rect 46734 31726 46786 31778
rect 47630 31726 47682 31778
rect 48078 31726 48130 31778
rect 3726 31614 3778 31666
rect 5854 31614 5906 31666
rect 7198 31614 7250 31666
rect 9214 31614 9266 31666
rect 11678 31614 11730 31666
rect 11902 31614 11954 31666
rect 16270 31614 16322 31666
rect 16942 31614 16994 31666
rect 18174 31614 18226 31666
rect 20750 31614 20802 31666
rect 21422 31614 21474 31666
rect 21646 31614 21698 31666
rect 21870 31614 21922 31666
rect 24782 31614 24834 31666
rect 28590 31614 28642 31666
rect 29150 31614 29202 31666
rect 30382 31614 30434 31666
rect 33070 31614 33122 31666
rect 33182 31614 33234 31666
rect 35646 31614 35698 31666
rect 45166 31614 45218 31666
rect 45614 31614 45666 31666
rect 46510 31614 46562 31666
rect 46958 31614 47010 31666
rect 2046 31502 2098 31554
rect 2158 31502 2210 31554
rect 2382 31502 2434 31554
rect 3390 31502 3442 31554
rect 3838 31502 3890 31554
rect 3950 31502 4002 31554
rect 4174 31502 4226 31554
rect 4734 31502 4786 31554
rect 5070 31502 5122 31554
rect 5966 31502 6018 31554
rect 11342 31502 11394 31554
rect 15262 31502 15314 31554
rect 20638 31502 20690 31554
rect 22206 31502 22258 31554
rect 22430 31502 22482 31554
rect 25566 31502 25618 31554
rect 29262 31502 29314 31554
rect 29486 31502 29538 31554
rect 32846 31502 32898 31554
rect 37438 31502 37490 31554
rect 37550 31502 37602 31554
rect 38222 31502 38274 31554
rect 39006 31502 39058 31554
rect 42702 31502 42754 31554
rect 44830 31502 44882 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 6862 31166 6914 31218
rect 7198 31166 7250 31218
rect 8766 31166 8818 31218
rect 17390 31166 17442 31218
rect 22766 31166 22818 31218
rect 25678 31166 25730 31218
rect 28254 31166 28306 31218
rect 30606 31166 30658 31218
rect 33966 31166 34018 31218
rect 34526 31166 34578 31218
rect 34638 31166 34690 31218
rect 44270 31166 44322 31218
rect 46174 31166 46226 31218
rect 48302 31166 48354 31218
rect 2494 31054 2546 31106
rect 7870 31054 7922 31106
rect 8206 31054 8258 31106
rect 16158 31054 16210 31106
rect 22094 31054 22146 31106
rect 22430 31054 22482 31106
rect 28030 31054 28082 31106
rect 30158 31054 30210 31106
rect 31166 31054 31218 31106
rect 33070 31054 33122 31106
rect 33294 31054 33346 31106
rect 34750 31054 34802 31106
rect 37214 31054 37266 31106
rect 38558 31054 38610 31106
rect 40238 31054 40290 31106
rect 44718 31054 44770 31106
rect 45614 31054 45666 31106
rect 45950 31054 46002 31106
rect 46398 31054 46450 31106
rect 47406 31054 47458 31106
rect 1710 30942 1762 30994
rect 5182 30942 5234 30994
rect 6078 30942 6130 30994
rect 6526 30942 6578 30994
rect 9662 30942 9714 30994
rect 15374 30942 15426 30994
rect 15822 30942 15874 30994
rect 16606 30942 16658 30994
rect 17614 30942 17666 30994
rect 17950 30942 18002 30994
rect 18734 30942 18786 30994
rect 21534 30942 21586 30994
rect 24110 30942 24162 30994
rect 26014 30942 26066 30994
rect 26798 30942 26850 30994
rect 27470 30942 27522 30994
rect 28254 30942 28306 30994
rect 28478 30942 28530 30994
rect 29710 30942 29762 30994
rect 30830 30942 30882 30994
rect 31726 30942 31778 30994
rect 32622 30942 32674 30994
rect 33182 30942 33234 30994
rect 33742 30942 33794 30994
rect 37886 30942 37938 30994
rect 38334 30942 38386 30994
rect 38894 30942 38946 30994
rect 39342 30942 39394 30994
rect 39566 30942 39618 30994
rect 41470 30942 41522 30994
rect 44158 30942 44210 30994
rect 44382 30942 44434 30994
rect 45054 30942 45106 30994
rect 45278 30942 45330 30994
rect 46510 30942 46562 30994
rect 4622 30830 4674 30882
rect 5294 30830 5346 30882
rect 10334 30830 10386 30882
rect 12462 30830 12514 30882
rect 13246 30830 13298 30882
rect 20078 30830 20130 30882
rect 21198 30830 21250 30882
rect 23214 30830 23266 30882
rect 23774 30830 23826 30882
rect 25342 30830 25394 30882
rect 26686 30830 26738 30882
rect 29486 30830 29538 30882
rect 31838 30830 31890 30882
rect 33854 30830 33906 30882
rect 35086 30830 35138 30882
rect 38446 30830 38498 30882
rect 42366 30830 42418 30882
rect 44830 30830 44882 30882
rect 46958 30830 47010 30882
rect 8430 30718 8482 30770
rect 17278 30718 17330 30770
rect 24334 30718 24386 30770
rect 43934 30718 43986 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 7646 30382 7698 30434
rect 7982 30382 8034 30434
rect 17166 30382 17218 30434
rect 20414 30382 20466 30434
rect 20750 30382 20802 30434
rect 22094 30382 22146 30434
rect 22318 30382 22370 30434
rect 24446 30382 24498 30434
rect 25230 30382 25282 30434
rect 43262 30382 43314 30434
rect 46062 30382 46114 30434
rect 46398 30382 46450 30434
rect 1934 30270 1986 30322
rect 3054 30270 3106 30322
rect 3390 30270 3442 30322
rect 4958 30270 5010 30322
rect 12350 30270 12402 30322
rect 13582 30270 13634 30322
rect 16606 30270 16658 30322
rect 19854 30270 19906 30322
rect 20302 30270 20354 30322
rect 21422 30270 21474 30322
rect 24782 30270 24834 30322
rect 28030 30270 28082 30322
rect 31390 30270 31442 30322
rect 31950 30270 32002 30322
rect 39902 30270 39954 30322
rect 42254 30270 42306 30322
rect 45278 30270 45330 30322
rect 2942 30158 2994 30210
rect 7086 30158 7138 30210
rect 7310 30158 7362 30210
rect 8654 30158 8706 30210
rect 9214 30158 9266 30210
rect 9662 30158 9714 30210
rect 9886 30158 9938 30210
rect 10334 30158 10386 30210
rect 10782 30158 10834 30210
rect 12126 30158 12178 30210
rect 12910 30158 12962 30210
rect 14478 30158 14530 30210
rect 15934 30158 15986 30210
rect 16494 30158 16546 30210
rect 17838 30158 17890 30210
rect 18062 30158 18114 30210
rect 20638 30158 20690 30210
rect 21310 30158 21362 30210
rect 21534 30158 21586 30210
rect 21982 30158 22034 30210
rect 23214 30158 23266 30210
rect 23550 30158 23602 30210
rect 25566 30158 25618 30210
rect 25790 30158 25842 30210
rect 26014 30158 26066 30210
rect 27134 30158 27186 30210
rect 27470 30158 27522 30210
rect 30382 30158 30434 30210
rect 30942 30158 30994 30210
rect 32062 30158 32114 30210
rect 32734 30158 32786 30210
rect 33294 30158 33346 30210
rect 34750 30158 34802 30210
rect 34974 30158 35026 30210
rect 35758 30158 35810 30210
rect 37102 30158 37154 30210
rect 40798 30158 40850 30210
rect 43486 30158 43538 30210
rect 43934 30158 43986 30210
rect 45166 30158 45218 30210
rect 45614 30158 45666 30210
rect 46286 30158 46338 30210
rect 46846 30158 46898 30210
rect 47070 30158 47122 30210
rect 47630 30158 47682 30210
rect 1822 30046 1874 30098
rect 2046 30046 2098 30098
rect 3838 30046 3890 30098
rect 4062 30046 4114 30098
rect 6414 30046 6466 30098
rect 6974 30046 7026 30098
rect 8766 30046 8818 30098
rect 10222 30046 10274 30098
rect 10670 30046 10722 30098
rect 11902 30046 11954 30098
rect 14926 30046 14978 30098
rect 15710 30046 15762 30098
rect 17726 30046 17778 30098
rect 18846 30046 18898 30098
rect 19406 30046 19458 30098
rect 22766 30046 22818 30098
rect 24558 30046 24610 30098
rect 26350 30046 26402 30098
rect 29934 30046 29986 30098
rect 31054 30046 31106 30098
rect 31950 30046 32002 30098
rect 37774 30046 37826 30098
rect 45054 30046 45106 30098
rect 45950 30046 46002 30098
rect 47182 30046 47234 30098
rect 3950 29934 4002 29986
rect 4510 29934 4562 29986
rect 5854 29934 5906 29986
rect 9550 29934 9602 29986
rect 11230 29934 11282 29986
rect 14142 29934 14194 29986
rect 15598 29934 15650 29986
rect 22430 29934 22482 29986
rect 23774 29934 23826 29986
rect 23998 29934 24050 29986
rect 26238 29934 26290 29986
rect 28590 29934 28642 29986
rect 29374 29934 29426 29986
rect 29598 29934 29650 29986
rect 29822 29934 29874 29986
rect 33630 29934 33682 29986
rect 35310 29934 35362 29986
rect 36542 29934 36594 29986
rect 45390 29934 45442 29986
rect 48078 29934 48130 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 6526 29598 6578 29650
rect 11790 29598 11842 29650
rect 16606 29598 16658 29650
rect 18062 29598 18114 29650
rect 20862 29598 20914 29650
rect 23326 29598 23378 29650
rect 23438 29598 23490 29650
rect 24110 29598 24162 29650
rect 24222 29598 24274 29650
rect 24334 29598 24386 29650
rect 25790 29598 25842 29650
rect 27134 29598 27186 29650
rect 28478 29598 28530 29650
rect 32286 29598 32338 29650
rect 35870 29598 35922 29650
rect 37438 29598 37490 29650
rect 46846 29598 46898 29650
rect 2494 29486 2546 29538
rect 4174 29486 4226 29538
rect 4846 29486 4898 29538
rect 5070 29486 5122 29538
rect 5294 29486 5346 29538
rect 6974 29486 7026 29538
rect 8430 29486 8482 29538
rect 9886 29486 9938 29538
rect 10222 29486 10274 29538
rect 13582 29486 13634 29538
rect 17950 29486 18002 29538
rect 18846 29486 18898 29538
rect 21198 29486 21250 29538
rect 29150 29486 29202 29538
rect 30158 29486 30210 29538
rect 31614 29486 31666 29538
rect 34078 29486 34130 29538
rect 36766 29486 36818 29538
rect 37774 29486 37826 29538
rect 40014 29486 40066 29538
rect 41134 29486 41186 29538
rect 42814 29486 42866 29538
rect 44158 29486 44210 29538
rect 2046 29374 2098 29426
rect 2158 29374 2210 29426
rect 2830 29374 2882 29426
rect 3614 29374 3666 29426
rect 6078 29374 6130 29426
rect 6302 29374 6354 29426
rect 6750 29374 6802 29426
rect 7982 29374 8034 29426
rect 8878 29374 8930 29426
rect 9550 29374 9602 29426
rect 10558 29374 10610 29426
rect 12350 29374 12402 29426
rect 12686 29374 12738 29426
rect 14366 29374 14418 29426
rect 15374 29374 15426 29426
rect 16382 29374 16434 29426
rect 17390 29374 17442 29426
rect 17838 29374 17890 29426
rect 18958 29374 19010 29426
rect 19070 29374 19122 29426
rect 19854 29374 19906 29426
rect 20190 29374 20242 29426
rect 21310 29374 21362 29426
rect 22318 29374 22370 29426
rect 23214 29374 23266 29426
rect 23774 29374 23826 29426
rect 24782 29374 24834 29426
rect 25678 29374 25730 29426
rect 25902 29374 25954 29426
rect 26238 29374 26290 29426
rect 27918 29374 27970 29426
rect 28814 29374 28866 29426
rect 33182 29374 33234 29426
rect 33630 29374 33682 29426
rect 34526 29374 34578 29426
rect 34750 29374 34802 29426
rect 35758 29374 35810 29426
rect 36318 29374 36370 29426
rect 37214 29374 37266 29426
rect 37438 29374 37490 29426
rect 38782 29374 38834 29426
rect 41246 29374 41298 29426
rect 41918 29374 41970 29426
rect 43374 29374 43426 29426
rect 46622 29374 46674 29426
rect 47070 29374 47122 29426
rect 47294 29374 47346 29426
rect 2382 29262 2434 29314
rect 3726 29262 3778 29314
rect 20414 29262 20466 29314
rect 21758 29262 21810 29314
rect 21870 29262 21922 29314
rect 25342 29262 25394 29314
rect 26574 29262 26626 29314
rect 27582 29262 27634 29314
rect 28142 29262 28194 29314
rect 29710 29262 29762 29314
rect 31838 29262 31890 29314
rect 35422 29262 35474 29314
rect 38110 29262 38162 29314
rect 40238 29262 40290 29314
rect 41694 29262 41746 29314
rect 42702 29262 42754 29314
rect 46286 29262 46338 29314
rect 47854 29262 47906 29314
rect 48190 29262 48242 29314
rect 5630 29150 5682 29202
rect 7198 29150 7250 29202
rect 18398 29150 18450 29202
rect 42590 29150 42642 29202
rect 47406 29150 47458 29202
rect 48078 29150 48130 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 4510 28814 4562 28866
rect 4846 28814 4898 28866
rect 9438 28814 9490 28866
rect 12910 28814 12962 28866
rect 20862 28814 20914 28866
rect 21982 28814 22034 28866
rect 22318 28814 22370 28866
rect 29374 28814 29426 28866
rect 30830 28814 30882 28866
rect 34750 28814 34802 28866
rect 1822 28702 1874 28754
rect 8430 28702 8482 28754
rect 10110 28702 10162 28754
rect 13582 28702 13634 28754
rect 16270 28702 16322 28754
rect 18062 28702 18114 28754
rect 19966 28702 20018 28754
rect 21422 28702 21474 28754
rect 26238 28702 26290 28754
rect 28478 28702 28530 28754
rect 29486 28702 29538 28754
rect 31614 28702 31666 28754
rect 32846 28702 32898 28754
rect 33742 28702 33794 28754
rect 34190 28702 34242 28754
rect 34414 28702 34466 28754
rect 36430 28702 36482 28754
rect 38110 28702 38162 28754
rect 41358 28702 41410 28754
rect 43934 28702 43986 28754
rect 46062 28702 46114 28754
rect 48190 28702 48242 28754
rect 3502 28590 3554 28642
rect 5070 28590 5122 28642
rect 5854 28590 5906 28642
rect 6078 28590 6130 28642
rect 6974 28590 7026 28642
rect 8542 28590 8594 28642
rect 9214 28590 9266 28642
rect 11678 28590 11730 28642
rect 13918 28590 13970 28642
rect 14366 28590 14418 28642
rect 17390 28590 17442 28642
rect 18398 28590 18450 28642
rect 21758 28590 21810 28642
rect 22654 28590 22706 28642
rect 23438 28590 23490 28642
rect 24110 28590 24162 28642
rect 26462 28590 26514 28642
rect 26686 28590 26738 28642
rect 27022 28590 27074 28642
rect 27806 28590 27858 28642
rect 28142 28590 28194 28642
rect 31054 28590 31106 28642
rect 31502 28590 31554 28642
rect 32398 28590 32450 28642
rect 33070 28590 33122 28642
rect 35310 28590 35362 28642
rect 35646 28590 35698 28642
rect 35870 28590 35922 28642
rect 37102 28590 37154 28642
rect 37662 28590 37714 28642
rect 38446 28590 38498 28642
rect 41694 28590 41746 28642
rect 43262 28590 43314 28642
rect 44046 28590 44098 28642
rect 44942 28590 44994 28642
rect 45390 28590 45442 28642
rect 2382 28478 2434 28530
rect 7086 28478 7138 28530
rect 10670 28478 10722 28530
rect 17054 28478 17106 28530
rect 19406 28478 19458 28530
rect 20302 28478 20354 28530
rect 22990 28478 23042 28530
rect 26910 28478 26962 28530
rect 29150 28478 29202 28530
rect 36990 28478 37042 28530
rect 39230 28478 39282 28530
rect 41918 28478 41970 28530
rect 42030 28478 42082 28530
rect 42702 28478 42754 28530
rect 42926 28478 42978 28530
rect 43598 28478 43650 28530
rect 3838 28366 3890 28418
rect 6190 28366 6242 28418
rect 6974 28366 7026 28418
rect 19070 28366 19122 28418
rect 20526 28366 20578 28418
rect 20750 28366 20802 28418
rect 28366 28366 28418 28418
rect 35534 28366 35586 28418
rect 37214 28366 37266 28418
rect 42814 28366 42866 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 5294 28030 5346 28082
rect 5966 28030 6018 28082
rect 9886 28030 9938 28082
rect 10222 28030 10274 28082
rect 11230 28030 11282 28082
rect 13806 28030 13858 28082
rect 18286 28030 18338 28082
rect 18510 28030 18562 28082
rect 20526 28030 20578 28082
rect 24558 28030 24610 28082
rect 24782 28030 24834 28082
rect 37998 28030 38050 28082
rect 38558 28030 38610 28082
rect 39118 28030 39170 28082
rect 39566 28030 39618 28082
rect 39790 28030 39842 28082
rect 40350 28030 40402 28082
rect 41022 28030 41074 28082
rect 41470 28030 41522 28082
rect 47518 28030 47570 28082
rect 3838 27918 3890 27970
rect 5182 27918 5234 27970
rect 6078 27918 6130 27970
rect 6750 27918 6802 27970
rect 8654 27918 8706 27970
rect 9662 27918 9714 27970
rect 11342 27918 11394 27970
rect 14254 27918 14306 27970
rect 17726 27918 17778 27970
rect 21422 27918 21474 27970
rect 24110 27918 24162 27970
rect 26350 27918 26402 27970
rect 27246 27918 27298 27970
rect 28702 27918 28754 27970
rect 29710 27918 29762 27970
rect 32062 27918 32114 27970
rect 34078 27918 34130 27970
rect 34190 27918 34242 27970
rect 36766 27918 36818 27970
rect 39006 27918 39058 27970
rect 39902 27918 39954 27970
rect 47854 27918 47906 27970
rect 4510 27806 4562 27858
rect 6862 27806 6914 27858
rect 7534 27806 7586 27858
rect 8542 27806 8594 27858
rect 8878 27806 8930 27858
rect 9550 27806 9602 27858
rect 10110 27806 10162 27858
rect 11006 27806 11058 27858
rect 12014 27806 12066 27858
rect 12574 27806 12626 27858
rect 12910 27806 12962 27858
rect 15150 27806 15202 27858
rect 17502 27806 17554 27858
rect 18622 27806 18674 27858
rect 19518 27806 19570 27858
rect 22430 27806 22482 27858
rect 22766 27806 22818 27858
rect 23550 27806 23602 27858
rect 24446 27806 24498 27858
rect 25902 27806 25954 27858
rect 26798 27806 26850 27858
rect 27358 27806 27410 27858
rect 27582 27806 27634 27858
rect 27806 27806 27858 27858
rect 28142 27806 28194 27858
rect 29822 27806 29874 27858
rect 31838 27806 31890 27858
rect 33182 27806 33234 27858
rect 33406 27806 33458 27858
rect 33630 27806 33682 27858
rect 33854 27806 33906 27858
rect 37438 27806 37490 27858
rect 38110 27806 38162 27858
rect 39342 27806 39394 27858
rect 41806 27806 41858 27858
rect 45838 27806 45890 27858
rect 46398 27806 46450 27858
rect 46510 27806 46562 27858
rect 46622 27806 46674 27858
rect 48190 27806 48242 27858
rect 1710 27694 1762 27746
rect 7422 27694 7474 27746
rect 13134 27694 13186 27746
rect 15486 27694 15538 27746
rect 16830 27694 16882 27746
rect 17950 27694 18002 27746
rect 19070 27694 19122 27746
rect 20638 27694 20690 27746
rect 23326 27694 23378 27746
rect 25566 27694 25618 27746
rect 27246 27694 27298 27746
rect 31054 27694 31106 27746
rect 33518 27694 33570 27746
rect 34638 27694 34690 27746
rect 42590 27694 42642 27746
rect 44718 27694 44770 27746
rect 5406 27582 5458 27634
rect 26574 27582 26626 27634
rect 26910 27582 26962 27634
rect 37998 27582 38050 27634
rect 45502 27582 45554 27634
rect 45614 27582 45666 27634
rect 45950 27582 46002 27634
rect 47070 27582 47122 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 20414 27246 20466 27298
rect 29374 27246 29426 27298
rect 30382 27246 30434 27298
rect 2046 27134 2098 27186
rect 6526 27134 6578 27186
rect 8318 27134 8370 27186
rect 13582 27134 13634 27186
rect 18398 27134 18450 27186
rect 19966 27134 20018 27186
rect 23326 27134 23378 27186
rect 25118 27134 25170 27186
rect 26462 27134 26514 27186
rect 27470 27134 27522 27186
rect 28030 27134 28082 27186
rect 29150 27134 29202 27186
rect 30942 27134 30994 27186
rect 32174 27134 32226 27186
rect 34302 27134 34354 27186
rect 40014 27134 40066 27186
rect 40462 27134 40514 27186
rect 42142 27134 42194 27186
rect 44270 27134 44322 27186
rect 46062 27134 46114 27186
rect 48190 27134 48242 27186
rect 3614 27022 3666 27074
rect 5070 27022 5122 27074
rect 5854 27022 5906 27074
rect 6974 27022 7026 27074
rect 7534 27022 7586 27074
rect 10446 27022 10498 27074
rect 10894 27022 10946 27074
rect 11790 27022 11842 27074
rect 12350 27022 12402 27074
rect 12686 27022 12738 27074
rect 13022 27022 13074 27074
rect 13694 27022 13746 27074
rect 15822 27022 15874 27074
rect 16494 27022 16546 27074
rect 17166 27022 17218 27074
rect 18062 27022 18114 27074
rect 18958 27022 19010 27074
rect 19182 27022 19234 27074
rect 19854 27022 19906 27074
rect 20078 27022 20130 27074
rect 22094 27022 22146 27074
rect 22542 27022 22594 27074
rect 23214 27022 23266 27074
rect 25342 27022 25394 27074
rect 26350 27022 26402 27074
rect 26574 27022 26626 27074
rect 28254 27022 28306 27074
rect 30606 27022 30658 27074
rect 35086 27022 35138 27074
rect 37214 27022 37266 27074
rect 40798 27022 40850 27074
rect 41470 27022 41522 27074
rect 45390 27022 45442 27074
rect 3166 26910 3218 26962
rect 4174 26910 4226 26962
rect 4846 26910 4898 26962
rect 5966 26910 6018 26962
rect 7646 26910 7698 26962
rect 12014 26910 12066 26962
rect 12798 26910 12850 26962
rect 15150 26910 15202 26962
rect 15598 26910 15650 26962
rect 17838 26910 17890 26962
rect 26798 26910 26850 26962
rect 27246 26910 27298 26962
rect 37886 26910 37938 26962
rect 44942 26910 44994 26962
rect 2494 26798 2546 26850
rect 4510 26798 4562 26850
rect 16382 26798 16434 26850
rect 17054 26798 17106 26850
rect 21534 26798 21586 26850
rect 27470 26798 27522 26850
rect 28590 26798 28642 26850
rect 29710 26798 29762 26850
rect 31838 26798 31890 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 4734 26462 4786 26514
rect 11118 26462 11170 26514
rect 24334 26462 24386 26514
rect 26686 26462 26738 26514
rect 33406 26462 33458 26514
rect 37662 26462 37714 26514
rect 38670 26462 38722 26514
rect 46734 26462 46786 26514
rect 6302 26350 6354 26402
rect 10222 26350 10274 26402
rect 10558 26350 10610 26402
rect 14254 26350 14306 26402
rect 16382 26350 16434 26402
rect 17278 26350 17330 26402
rect 19518 26350 19570 26402
rect 26238 26350 26290 26402
rect 31390 26350 31442 26402
rect 35758 26350 35810 26402
rect 37550 26350 37602 26402
rect 37774 26350 37826 26402
rect 38222 26350 38274 26402
rect 38894 26350 38946 26402
rect 39566 26350 39618 26402
rect 42366 26350 42418 26402
rect 42814 26350 42866 26402
rect 45614 26350 45666 26402
rect 47070 26350 47122 26402
rect 2270 26238 2322 26290
rect 3054 26238 3106 26290
rect 4174 26238 4226 26290
rect 4622 26238 4674 26290
rect 6078 26238 6130 26290
rect 6414 26238 6466 26290
rect 8206 26238 8258 26290
rect 8990 26238 9042 26290
rect 11566 26238 11618 26290
rect 12126 26238 12178 26290
rect 15150 26238 15202 26290
rect 15710 26238 15762 26290
rect 16046 26238 16098 26290
rect 17614 26238 17666 26290
rect 19070 26238 19122 26290
rect 19406 26238 19458 26290
rect 19742 26238 19794 26290
rect 20302 26238 20354 26290
rect 20526 26238 20578 26290
rect 20638 26238 20690 26290
rect 21534 26238 21586 26290
rect 22318 26238 22370 26290
rect 22766 26238 22818 26290
rect 23214 26238 23266 26290
rect 23998 26238 24050 26290
rect 26574 26238 26626 26290
rect 26798 26238 26850 26290
rect 27246 26238 27298 26290
rect 27470 26238 27522 26290
rect 28590 26238 28642 26290
rect 30270 26238 30322 26290
rect 30606 26238 30658 26290
rect 31838 26238 31890 26290
rect 32958 26238 33010 26290
rect 33518 26238 33570 26290
rect 33630 26238 33682 26290
rect 34974 26238 35026 26290
rect 35422 26238 35474 26290
rect 35870 26238 35922 26290
rect 36430 26238 36482 26290
rect 37214 26238 37266 26290
rect 38446 26238 38498 26290
rect 39006 26238 39058 26290
rect 43262 26238 43314 26290
rect 46174 26238 46226 26290
rect 48190 26238 48242 26290
rect 2942 26126 2994 26178
rect 12462 26126 12514 26178
rect 16494 26126 16546 26178
rect 21422 26126 21474 26178
rect 23774 26126 23826 26178
rect 25454 26126 25506 26178
rect 25790 26126 25842 26178
rect 27582 26126 27634 26178
rect 32174 26126 32226 26178
rect 34078 26126 34130 26178
rect 34526 26126 34578 26178
rect 38110 26126 38162 26178
rect 39454 26126 39506 26178
rect 40014 26126 40066 26178
rect 41918 26126 41970 26178
rect 42142 26126 42194 26178
rect 42478 26126 42530 26178
rect 43710 26126 43762 26178
rect 4734 26014 4786 26066
rect 10782 26014 10834 26066
rect 20078 26014 20130 26066
rect 20862 26014 20914 26066
rect 22878 26014 22930 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 6974 25678 7026 25730
rect 12798 25678 12850 25730
rect 13918 25678 13970 25730
rect 17726 25678 17778 25730
rect 23214 25678 23266 25730
rect 26238 25678 26290 25730
rect 29486 25678 29538 25730
rect 47630 25678 47682 25730
rect 2494 25566 2546 25618
rect 4622 25566 4674 25618
rect 8654 25566 8706 25618
rect 14254 25566 14306 25618
rect 21870 25566 21922 25618
rect 24558 25566 24610 25618
rect 27582 25566 27634 25618
rect 29598 25566 29650 25618
rect 31166 25566 31218 25618
rect 35982 25566 36034 25618
rect 39230 25566 39282 25618
rect 43486 25566 43538 25618
rect 43934 25566 43986 25618
rect 44382 25566 44434 25618
rect 46398 25566 46450 25618
rect 47294 25566 47346 25618
rect 48190 25566 48242 25618
rect 1822 25454 1874 25506
rect 5742 25454 5794 25506
rect 6302 25454 6354 25506
rect 6638 25454 6690 25506
rect 7758 25454 7810 25506
rect 8542 25454 8594 25506
rect 11118 25454 11170 25506
rect 12910 25454 12962 25506
rect 14702 25454 14754 25506
rect 17502 25454 17554 25506
rect 18174 25454 18226 25506
rect 19966 25454 20018 25506
rect 21758 25454 21810 25506
rect 23438 25454 23490 25506
rect 24670 25454 24722 25506
rect 25006 25454 25058 25506
rect 26014 25454 26066 25506
rect 26686 25454 26738 25506
rect 29486 25454 29538 25506
rect 30494 25454 30546 25506
rect 30718 25454 30770 25506
rect 32286 25454 32338 25506
rect 34526 25454 34578 25506
rect 34974 25454 35026 25506
rect 36990 25454 37042 25506
rect 40238 25454 40290 25506
rect 40910 25454 40962 25506
rect 45054 25454 45106 25506
rect 45166 25454 45218 25506
rect 45614 25454 45666 25506
rect 46510 25454 46562 25506
rect 46846 25454 46898 25506
rect 47406 25454 47458 25506
rect 5966 25342 6018 25394
rect 9438 25342 9490 25394
rect 12238 25342 12290 25394
rect 13694 25342 13746 25394
rect 16270 25342 16322 25394
rect 16942 25342 16994 25394
rect 19182 25342 19234 25394
rect 27918 25342 27970 25394
rect 28590 25342 28642 25394
rect 31278 25342 31330 25394
rect 32174 25342 32226 25394
rect 33630 25342 33682 25394
rect 35422 25342 35474 25394
rect 35534 25342 35586 25394
rect 41918 25342 41970 25394
rect 44942 25342 44994 25394
rect 45838 25342 45890 25394
rect 46286 25342 46338 25394
rect 5070 25230 5122 25282
rect 18286 25230 18338 25282
rect 28254 25230 28306 25282
rect 31054 25230 31106 25282
rect 33518 25230 33570 25282
rect 35198 25230 35250 25282
rect 36542 25230 36594 25282
rect 37102 25230 37154 25282
rect 37214 25230 37266 25282
rect 37438 25230 37490 25282
rect 39790 25230 39842 25282
rect 40462 25230 40514 25282
rect 41134 25230 41186 25282
rect 41582 25230 41634 25282
rect 47294 25230 47346 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 2158 24894 2210 24946
rect 2606 24894 2658 24946
rect 5630 24894 5682 24946
rect 6526 24894 6578 24946
rect 9774 24894 9826 24946
rect 13022 24894 13074 24946
rect 16830 24894 16882 24946
rect 17502 24894 17554 24946
rect 19518 24894 19570 24946
rect 31838 24894 31890 24946
rect 34862 24894 34914 24946
rect 46958 24894 47010 24946
rect 2942 24782 2994 24834
rect 3838 24782 3890 24834
rect 6974 24782 7026 24834
rect 12574 24782 12626 24834
rect 16494 24782 16546 24834
rect 17614 24782 17666 24834
rect 18286 24782 18338 24834
rect 18958 24782 19010 24834
rect 19966 24782 20018 24834
rect 23662 24782 23714 24834
rect 28814 24782 28866 24834
rect 31166 24782 31218 24834
rect 31502 24782 31554 24834
rect 33742 24782 33794 24834
rect 40350 24782 40402 24834
rect 2270 24670 2322 24722
rect 2718 24670 2770 24722
rect 3390 24670 3442 24722
rect 5070 24670 5122 24722
rect 6526 24670 6578 24722
rect 8206 24670 8258 24722
rect 9438 24670 9490 24722
rect 9886 24670 9938 24722
rect 10110 24670 10162 24722
rect 13134 24670 13186 24722
rect 14030 24670 14082 24722
rect 15934 24670 15986 24722
rect 17502 24670 17554 24722
rect 19070 24670 19122 24722
rect 20862 24670 20914 24722
rect 22654 24670 22706 24722
rect 23102 24670 23154 24722
rect 23550 24670 23602 24722
rect 24446 24670 24498 24722
rect 25230 24670 25282 24722
rect 30942 24670 30994 24722
rect 33630 24670 33682 24722
rect 34302 24670 34354 24722
rect 35086 24670 35138 24722
rect 38782 24670 38834 24722
rect 39118 24670 39170 24722
rect 39678 24670 39730 24722
rect 40014 24670 40066 24722
rect 40910 24670 40962 24722
rect 41470 24670 41522 24722
rect 42254 24670 42306 24722
rect 45950 24670 46002 24722
rect 47294 24670 47346 24722
rect 47518 24670 47570 24722
rect 47966 24670 48018 24722
rect 11342 24558 11394 24610
rect 14142 24558 14194 24610
rect 15598 24558 15650 24610
rect 21198 24558 21250 24610
rect 23886 24558 23938 24610
rect 32510 24558 32562 24610
rect 33854 24558 33906 24610
rect 34750 24558 34802 24610
rect 35870 24558 35922 24610
rect 37998 24558 38050 24610
rect 43038 24558 43090 24610
rect 45166 24558 45218 24610
rect 46398 24558 46450 24610
rect 18958 24446 19010 24498
rect 45614 24446 45666 24498
rect 47854 24446 47906 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 2382 24110 2434 24162
rect 6190 24110 6242 24162
rect 8990 24110 9042 24162
rect 11566 24110 11618 24162
rect 19630 24110 19682 24162
rect 29934 24110 29986 24162
rect 37214 24110 37266 24162
rect 37886 24110 37938 24162
rect 43150 24110 43202 24162
rect 43486 24110 43538 24162
rect 4958 23998 5010 24050
rect 8094 23998 8146 24050
rect 12014 23998 12066 24050
rect 14142 23998 14194 24050
rect 18846 23998 18898 24050
rect 20190 23998 20242 24050
rect 24446 23998 24498 24050
rect 24558 23998 24610 24050
rect 29150 23998 29202 24050
rect 30942 23998 30994 24050
rect 31390 23998 31442 24050
rect 32286 23998 32338 24050
rect 32734 23998 32786 24050
rect 33070 23998 33122 24050
rect 36990 23998 37042 24050
rect 37998 23998 38050 24050
rect 40574 23998 40626 24050
rect 42142 23998 42194 24050
rect 45054 23998 45106 24050
rect 46062 23998 46114 24050
rect 48190 23998 48242 24050
rect 4286 23886 4338 23938
rect 4510 23886 4562 23938
rect 7758 23886 7810 23938
rect 9662 23886 9714 23938
rect 10558 23886 10610 23938
rect 11678 23886 11730 23938
rect 12462 23886 12514 23938
rect 13470 23886 13522 23938
rect 14702 23886 14754 23938
rect 15038 23886 15090 23938
rect 16046 23886 16098 23938
rect 19742 23886 19794 23938
rect 20078 23886 20130 23938
rect 21422 23886 21474 23938
rect 21870 23886 21922 23938
rect 22654 23886 22706 23938
rect 23102 23886 23154 23938
rect 23774 23886 23826 23938
rect 25006 23886 25058 23938
rect 26798 23886 26850 23938
rect 27134 23886 27186 23938
rect 30270 23886 30322 23938
rect 30606 23886 30658 23938
rect 31726 23886 31778 23938
rect 35870 23886 35922 23938
rect 38222 23886 38274 23938
rect 41582 23886 41634 23938
rect 42702 23886 42754 23938
rect 43150 23886 43202 23938
rect 45390 23886 45442 23938
rect 5630 23774 5682 23826
rect 10894 23774 10946 23826
rect 13582 23774 13634 23826
rect 15374 23774 15426 23826
rect 15486 23774 15538 23826
rect 16718 23774 16770 23826
rect 21310 23774 21362 23826
rect 23438 23774 23490 23826
rect 24222 23774 24274 23826
rect 27582 23774 27634 23826
rect 30830 23774 30882 23826
rect 35198 23774 35250 23826
rect 37550 23774 37602 23826
rect 4846 23662 4898 23714
rect 5070 23662 5122 23714
rect 15710 23662 15762 23714
rect 23326 23662 23378 23714
rect 27022 23662 27074 23714
rect 29710 23662 29762 23714
rect 40126 23662 40178 23714
rect 41134 23662 41186 23714
rect 42478 23662 42530 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 8318 23326 8370 23378
rect 12350 23326 12402 23378
rect 22766 23326 22818 23378
rect 23214 23326 23266 23378
rect 35758 23326 35810 23378
rect 44382 23326 44434 23378
rect 46062 23326 46114 23378
rect 7422 23214 7474 23266
rect 9550 23214 9602 23266
rect 12798 23214 12850 23266
rect 18398 23214 18450 23266
rect 22430 23214 22482 23266
rect 22878 23214 22930 23266
rect 24670 23214 24722 23266
rect 26014 23214 26066 23266
rect 26574 23214 26626 23266
rect 28478 23214 28530 23266
rect 30046 23214 30098 23266
rect 31278 23214 31330 23266
rect 31726 23214 31778 23266
rect 38110 23214 38162 23266
rect 44942 23214 44994 23266
rect 45838 23214 45890 23266
rect 47182 23214 47234 23266
rect 47966 23214 48018 23266
rect 1822 23102 1874 23154
rect 6190 23102 6242 23154
rect 7982 23102 8034 23154
rect 12238 23102 12290 23154
rect 14142 23102 14194 23154
rect 16606 23102 16658 23154
rect 17838 23102 17890 23154
rect 18846 23102 18898 23154
rect 22654 23102 22706 23154
rect 24110 23102 24162 23154
rect 24334 23102 24386 23154
rect 25566 23102 25618 23154
rect 25902 23102 25954 23154
rect 27134 23102 27186 23154
rect 28254 23102 28306 23154
rect 30270 23102 30322 23154
rect 30942 23102 30994 23154
rect 32510 23102 32562 23154
rect 32958 23102 33010 23154
rect 33406 23102 33458 23154
rect 33630 23102 33682 23154
rect 34414 23102 34466 23154
rect 38334 23102 38386 23154
rect 38558 23102 38610 23154
rect 38894 23102 38946 23154
rect 41022 23102 41074 23154
rect 45166 23102 45218 23154
rect 45502 23102 45554 23154
rect 46398 23102 46450 23154
rect 46734 23102 46786 23154
rect 47630 23102 47682 23154
rect 2494 22990 2546 23042
rect 4734 22990 4786 23042
rect 8206 22990 8258 23042
rect 12014 22990 12066 23042
rect 14478 22990 14530 23042
rect 16382 22990 16434 23042
rect 17950 22990 18002 23042
rect 19518 22990 19570 23042
rect 21646 22990 21698 23042
rect 23774 22990 23826 23042
rect 30830 22990 30882 23042
rect 33518 22990 33570 23042
rect 33966 22990 34018 23042
rect 35310 22990 35362 23042
rect 35982 22990 36034 23042
rect 36206 22990 36258 23042
rect 10110 22878 10162 22930
rect 23550 22878 23602 22930
rect 24558 22878 24610 22930
rect 36654 22990 36706 23042
rect 37102 22990 37154 23042
rect 38446 22990 38498 23042
rect 39118 22990 39170 23042
rect 41694 22990 41746 23042
rect 43822 22990 43874 23042
rect 44270 22990 44322 23042
rect 45054 22990 45106 23042
rect 47406 22990 47458 23042
rect 36654 22878 36706 22930
rect 39230 22878 39282 22930
rect 44158 22878 44210 22930
rect 45726 22878 45778 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 3390 22542 3442 22594
rect 11118 22542 11170 22594
rect 15150 22542 15202 22594
rect 29598 22542 29650 22594
rect 34974 22542 35026 22594
rect 40574 22542 40626 22594
rect 45950 22542 46002 22594
rect 46622 22542 46674 22594
rect 1822 22430 1874 22482
rect 2830 22430 2882 22482
rect 3950 22430 4002 22482
rect 6078 22430 6130 22482
rect 7758 22430 7810 22482
rect 9998 22430 10050 22482
rect 12910 22430 12962 22482
rect 15262 22430 15314 22482
rect 18734 22430 18786 22482
rect 19966 22430 20018 22482
rect 24446 22430 24498 22482
rect 31390 22430 31442 22482
rect 31726 22430 31778 22482
rect 35086 22430 35138 22482
rect 37214 22430 37266 22482
rect 39342 22430 39394 22482
rect 41134 22430 41186 22482
rect 42254 22430 42306 22482
rect 43598 22430 43650 22482
rect 46958 22430 47010 22482
rect 2382 22318 2434 22370
rect 2942 22318 2994 22370
rect 4510 22318 4562 22370
rect 4846 22318 4898 22370
rect 5630 22318 5682 22370
rect 10670 22318 10722 22370
rect 11678 22318 11730 22370
rect 13470 22318 13522 22370
rect 15934 22318 15986 22370
rect 19742 22318 19794 22370
rect 20078 22318 20130 22370
rect 20414 22318 20466 22370
rect 21534 22318 21586 22370
rect 26350 22318 26402 22370
rect 28142 22318 28194 22370
rect 29262 22318 29314 22370
rect 29710 22318 29762 22370
rect 30606 22318 30658 22370
rect 30830 22318 30882 22370
rect 34526 22318 34578 22370
rect 35310 22318 35362 22370
rect 35758 22318 35810 22370
rect 40126 22318 40178 22370
rect 43150 22318 43202 22370
rect 43374 22318 43426 22370
rect 43934 22318 43986 22370
rect 45502 22318 45554 22370
rect 45726 22318 45778 22370
rect 47182 22318 47234 22370
rect 47518 22318 47570 22370
rect 47742 22318 47794 22370
rect 14254 22206 14306 22258
rect 16606 22206 16658 22258
rect 19070 22206 19122 22258
rect 22318 22206 22370 22258
rect 25230 22206 25282 22258
rect 27582 22206 27634 22258
rect 33854 22206 33906 22258
rect 40462 22206 40514 22258
rect 40574 22206 40626 22258
rect 44270 22206 44322 22258
rect 44830 22206 44882 22258
rect 45054 22206 45106 22258
rect 46846 22206 46898 22258
rect 3838 22094 3890 22146
rect 12350 22094 12402 22146
rect 15374 22094 15426 22146
rect 19406 22094 19458 22146
rect 24894 22094 24946 22146
rect 25118 22094 25170 22146
rect 26686 22094 26738 22146
rect 28702 22094 28754 22146
rect 36206 22094 36258 22146
rect 36318 22094 36370 22146
rect 36430 22094 36482 22146
rect 44046 22094 44098 22146
rect 44942 22094 44994 22146
rect 46398 22094 46450 22146
rect 47518 22094 47570 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 8318 21758 8370 21810
rect 9774 21758 9826 21810
rect 10782 21758 10834 21810
rect 17390 21758 17442 21810
rect 17502 21758 17554 21810
rect 18398 21758 18450 21810
rect 18734 21758 18786 21810
rect 24334 21758 24386 21810
rect 25342 21758 25394 21810
rect 27358 21758 27410 21810
rect 30382 21758 30434 21810
rect 32174 21758 32226 21810
rect 33518 21758 33570 21810
rect 42254 21758 42306 21810
rect 46622 21758 46674 21810
rect 6974 21646 7026 21698
rect 11118 21646 11170 21698
rect 17614 21646 17666 21698
rect 17726 21646 17778 21698
rect 18510 21646 18562 21698
rect 19406 21646 19458 21698
rect 19518 21646 19570 21698
rect 20526 21646 20578 21698
rect 21198 21646 21250 21698
rect 21646 21646 21698 21698
rect 22094 21646 22146 21698
rect 22206 21646 22258 21698
rect 23662 21646 23714 21698
rect 23998 21646 24050 21698
rect 25118 21646 25170 21698
rect 26686 21646 26738 21698
rect 29038 21646 29090 21698
rect 30494 21646 30546 21698
rect 32398 21646 32450 21698
rect 37326 21646 37378 21698
rect 37886 21646 37938 21698
rect 41134 21646 41186 21698
rect 44046 21646 44098 21698
rect 47518 21646 47570 21698
rect 47854 21646 47906 21698
rect 4734 21534 4786 21586
rect 5294 21534 5346 21586
rect 5518 21534 5570 21586
rect 7870 21534 7922 21586
rect 8206 21534 8258 21586
rect 9662 21534 9714 21586
rect 9886 21534 9938 21586
rect 10222 21534 10274 21586
rect 11678 21534 11730 21586
rect 12014 21534 12066 21586
rect 15710 21534 15762 21586
rect 18062 21534 18114 21586
rect 18958 21534 19010 21586
rect 19294 21534 19346 21586
rect 19742 21534 19794 21586
rect 20078 21534 20130 21586
rect 21422 21534 21474 21586
rect 21870 21534 21922 21586
rect 22542 21534 22594 21586
rect 23886 21534 23938 21586
rect 24558 21534 24610 21586
rect 25454 21534 25506 21586
rect 26014 21534 26066 21586
rect 27582 21534 27634 21586
rect 29598 21534 29650 21586
rect 30718 21534 30770 21586
rect 31054 21534 31106 21586
rect 31838 21534 31890 21586
rect 32510 21534 32562 21586
rect 33182 21534 33234 21586
rect 33294 21534 33346 21586
rect 33742 21534 33794 21586
rect 34190 21534 34242 21586
rect 37662 21534 37714 21586
rect 39230 21534 39282 21586
rect 43262 21534 43314 21586
rect 46958 21534 47010 21586
rect 47182 21534 47234 21586
rect 48078 21534 48130 21586
rect 1934 21422 1986 21474
rect 4062 21422 4114 21474
rect 12798 21422 12850 21474
rect 14926 21422 14978 21474
rect 22206 21422 22258 21474
rect 31502 21422 31554 21474
rect 34862 21422 34914 21474
rect 36990 21422 37042 21474
rect 37774 21422 37826 21474
rect 39006 21422 39058 21474
rect 39790 21422 39842 21474
rect 40910 21422 40962 21474
rect 41694 21422 41746 21474
rect 46174 21422 46226 21474
rect 47070 21422 47122 21474
rect 5854 21310 5906 21362
rect 16494 21310 16546 21362
rect 41246 21310 41298 21362
rect 41806 21310 41858 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 6302 20974 6354 21026
rect 10334 20974 10386 21026
rect 20526 20974 20578 21026
rect 42814 20974 42866 21026
rect 4846 20862 4898 20914
rect 10222 20862 10274 20914
rect 13022 20862 13074 20914
rect 15710 20862 15762 20914
rect 21758 20862 21810 20914
rect 22766 20862 22818 20914
rect 23326 20862 23378 20914
rect 27694 20862 27746 20914
rect 30158 20862 30210 20914
rect 32062 20862 32114 20914
rect 33182 20862 33234 20914
rect 38334 20862 38386 20914
rect 39230 20862 39282 20914
rect 41358 20862 41410 20914
rect 42478 20862 42530 20914
rect 44382 20862 44434 20914
rect 45054 20862 45106 20914
rect 48190 20862 48242 20914
rect 2046 20750 2098 20802
rect 6078 20750 6130 20802
rect 6302 20750 6354 20802
rect 6750 20750 6802 20802
rect 7758 20750 7810 20802
rect 8654 20750 8706 20802
rect 9774 20750 9826 20802
rect 12910 20750 12962 20802
rect 18622 20750 18674 20802
rect 18958 20750 19010 20802
rect 20190 20750 20242 20802
rect 21534 20750 21586 20802
rect 22206 20750 22258 20802
rect 23774 20750 23826 20802
rect 25342 20750 25394 20802
rect 25566 20750 25618 20802
rect 28030 20750 28082 20802
rect 28478 20750 28530 20802
rect 29374 20750 29426 20802
rect 31614 20750 31666 20802
rect 32286 20750 32338 20802
rect 32622 20750 32674 20802
rect 33630 20750 33682 20802
rect 33966 20750 34018 20802
rect 35422 20750 35474 20802
rect 36318 20750 36370 20802
rect 36990 20750 37042 20802
rect 38110 20750 38162 20802
rect 38446 20750 38498 20802
rect 42030 20750 42082 20802
rect 45390 20750 45442 20802
rect 2718 20638 2770 20690
rect 11902 20638 11954 20690
rect 12350 20638 12402 20690
rect 13470 20638 13522 20690
rect 15374 20638 15426 20690
rect 17838 20638 17890 20690
rect 19070 20638 19122 20690
rect 24110 20638 24162 20690
rect 24222 20638 24274 20690
rect 26126 20638 26178 20690
rect 30606 20638 30658 20690
rect 31166 20638 31218 20690
rect 34190 20638 34242 20690
rect 34638 20638 34690 20690
rect 37326 20638 37378 20690
rect 37886 20638 37938 20690
rect 42590 20638 42642 20690
rect 46062 20638 46114 20690
rect 14030 20526 14082 20578
rect 15038 20526 15090 20578
rect 19518 20526 19570 20578
rect 27022 20526 27074 20578
rect 32062 20526 32114 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 2494 20190 2546 20242
rect 3278 20190 3330 20242
rect 7758 20190 7810 20242
rect 9886 20190 9938 20242
rect 15710 20190 15762 20242
rect 6862 20078 6914 20130
rect 11118 20078 11170 20130
rect 11566 20078 11618 20130
rect 11902 20078 11954 20130
rect 17950 20078 18002 20130
rect 18622 20078 18674 20130
rect 18734 20078 18786 20130
rect 19182 20078 19234 20130
rect 19294 20134 19346 20186
rect 20302 20190 20354 20242
rect 26238 20190 26290 20242
rect 30494 20190 30546 20242
rect 46398 20190 46450 20242
rect 47294 20190 47346 20242
rect 19406 20078 19458 20130
rect 24110 20078 24162 20130
rect 24446 20078 24498 20130
rect 25230 20078 25282 20130
rect 25342 20078 25394 20130
rect 31838 20078 31890 20130
rect 34078 20078 34130 20130
rect 34414 20078 34466 20130
rect 34526 20078 34578 20130
rect 34638 20078 34690 20130
rect 35310 20078 35362 20130
rect 36094 20078 36146 20130
rect 38446 20078 38498 20130
rect 38782 20078 38834 20130
rect 42478 20078 42530 20130
rect 46734 20078 46786 20130
rect 47182 20078 47234 20130
rect 47518 20078 47570 20130
rect 47854 20078 47906 20130
rect 4398 19966 4450 20018
rect 5742 19966 5794 20018
rect 7870 19966 7922 20018
rect 9886 19966 9938 20018
rect 10558 19966 10610 20018
rect 10894 19966 10946 20018
rect 12126 19966 12178 20018
rect 16270 19966 16322 20018
rect 16830 19966 16882 20018
rect 17390 19966 17442 20018
rect 17726 19966 17778 20018
rect 18174 19966 18226 20018
rect 18398 19966 18450 20018
rect 19070 19966 19122 20018
rect 19854 19966 19906 20018
rect 20190 19966 20242 20018
rect 20750 19966 20802 20018
rect 23886 19966 23938 20018
rect 24334 19966 24386 20018
rect 26462 19966 26514 20018
rect 26798 19966 26850 20018
rect 27470 19966 27522 20018
rect 27694 19966 27746 20018
rect 30158 19966 30210 20018
rect 31390 19966 31442 20018
rect 32062 19966 32114 20018
rect 33518 19966 33570 20018
rect 37214 19966 37266 20018
rect 39006 19966 39058 20018
rect 41806 19966 41858 20018
rect 45054 19966 45106 20018
rect 45278 19966 45330 20018
rect 46510 19966 46562 20018
rect 46846 19966 46898 20018
rect 47742 19966 47794 20018
rect 2158 19854 2210 19906
rect 3838 19854 3890 19906
rect 5294 19854 5346 19906
rect 8094 19854 8146 19906
rect 13022 19854 13074 19906
rect 17838 19854 17890 19906
rect 21422 19854 21474 19906
rect 23550 19854 23602 19906
rect 24670 19854 24722 19906
rect 26910 19854 26962 19906
rect 28590 19854 28642 19906
rect 28926 19854 28978 19906
rect 31054 19854 31106 19906
rect 31950 19854 32002 19906
rect 32510 19854 32562 19906
rect 33182 19854 33234 19906
rect 35646 19854 35698 19906
rect 36542 19854 36594 19906
rect 37438 19854 37490 19906
rect 37886 19854 37938 19906
rect 39566 19854 39618 19906
rect 40014 19854 40066 19906
rect 41022 19854 41074 19906
rect 44606 19854 44658 19906
rect 25342 19742 25394 19794
rect 28030 19742 28082 19794
rect 32398 19742 32450 19794
rect 37550 19742 37602 19794
rect 38110 19742 38162 19794
rect 45054 19742 45106 19794
rect 47854 19742 47906 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 15934 19406 15986 19458
rect 27358 19406 27410 19458
rect 29150 19406 29202 19458
rect 43934 19406 43986 19458
rect 1710 19294 1762 19346
rect 5182 19294 5234 19346
rect 5630 19294 5682 19346
rect 11230 19294 11282 19346
rect 12910 19294 12962 19346
rect 17166 19294 17218 19346
rect 18846 19294 18898 19346
rect 19294 19294 19346 19346
rect 20526 19294 20578 19346
rect 21310 19294 21362 19346
rect 24558 19294 24610 19346
rect 26686 19294 26738 19346
rect 28142 19294 28194 19346
rect 29710 19294 29762 19346
rect 30158 19294 30210 19346
rect 30942 19294 30994 19346
rect 35422 19294 35474 19346
rect 37774 19294 37826 19346
rect 39902 19294 39954 19346
rect 40238 19294 40290 19346
rect 43710 19294 43762 19346
rect 48190 19294 48242 19346
rect 4510 19182 4562 19234
rect 7086 19182 7138 19234
rect 8430 19182 8482 19234
rect 13694 19182 13746 19234
rect 15262 19182 15314 19234
rect 16382 19182 16434 19234
rect 16718 19182 16770 19234
rect 16942 19182 16994 19234
rect 18622 19182 18674 19234
rect 19742 19182 19794 19234
rect 20190 19182 20242 19234
rect 21422 19182 21474 19234
rect 22094 19182 22146 19234
rect 23326 19182 23378 19234
rect 23886 19182 23938 19234
rect 27582 19182 27634 19234
rect 27918 19182 27970 19234
rect 29486 19182 29538 19234
rect 30494 19182 30546 19234
rect 33854 19182 33906 19234
rect 36990 19182 37042 19234
rect 43038 19182 43090 19234
rect 45390 19182 45442 19234
rect 3838 19070 3890 19122
rect 5966 19070 6018 19122
rect 6078 19070 6130 19122
rect 6190 19070 6242 19122
rect 7534 19070 7586 19122
rect 7646 19070 7698 19122
rect 7758 19070 7810 19122
rect 9102 19070 9154 19122
rect 11678 19070 11730 19122
rect 12462 19070 12514 19122
rect 12574 19070 12626 19122
rect 15486 19070 15538 19122
rect 21758 19070 21810 19122
rect 22766 19070 22818 19122
rect 23102 19070 23154 19122
rect 33070 19070 33122 19122
rect 34190 19070 34242 19122
rect 34526 19070 34578 19122
rect 34974 19070 35026 19122
rect 42366 19070 42418 19122
rect 46062 19070 46114 19122
rect 6414 18958 6466 19010
rect 7870 18958 7922 19010
rect 11790 18958 11842 19010
rect 12126 18958 12178 19010
rect 12350 18958 12402 19010
rect 16494 18958 16546 19010
rect 17502 18958 17554 19010
rect 18174 18958 18226 19010
rect 18286 18958 18338 19010
rect 18398 18958 18450 19010
rect 21870 18958 21922 19010
rect 22430 18958 22482 19010
rect 34862 18958 34914 19010
rect 35870 18958 35922 19010
rect 36318 18958 36370 19010
rect 44270 18958 44322 19010
rect 45054 18958 45106 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 5854 18622 5906 18674
rect 6526 18622 6578 18674
rect 7086 18622 7138 18674
rect 18510 18622 18562 18674
rect 24110 18622 24162 18674
rect 31502 18622 31554 18674
rect 33070 18622 33122 18674
rect 38110 18622 38162 18674
rect 38894 18622 38946 18674
rect 45166 18622 45218 18674
rect 46174 18622 46226 18674
rect 7310 18510 7362 18562
rect 7422 18510 7474 18562
rect 7646 18510 7698 18562
rect 20862 18510 20914 18562
rect 21198 18510 21250 18562
rect 22878 18510 22930 18562
rect 23550 18510 23602 18562
rect 24446 18510 24498 18562
rect 31838 18510 31890 18562
rect 32510 18510 32562 18562
rect 33406 18510 33458 18562
rect 38334 18510 38386 18562
rect 39006 18510 39058 18562
rect 44494 18510 44546 18562
rect 45502 18510 45554 18562
rect 47070 18510 47122 18562
rect 47854 18510 47906 18562
rect 2046 18398 2098 18450
rect 2494 18398 2546 18450
rect 6526 18398 6578 18450
rect 8654 18398 8706 18450
rect 9662 18398 9714 18450
rect 12574 18398 12626 18450
rect 12798 18398 12850 18450
rect 13918 18398 13970 18450
rect 14590 18398 14642 18450
rect 17614 18398 17666 18450
rect 18062 18398 18114 18450
rect 18846 18398 18898 18450
rect 19630 18398 19682 18450
rect 19854 18398 19906 18450
rect 20302 18398 20354 18450
rect 21422 18398 21474 18450
rect 22766 18398 22818 18450
rect 23326 18398 23378 18450
rect 23886 18398 23938 18450
rect 24334 18398 24386 18450
rect 25342 18398 25394 18450
rect 29038 18398 29090 18450
rect 29598 18398 29650 18450
rect 30382 18398 30434 18450
rect 30830 18398 30882 18450
rect 31166 18398 31218 18450
rect 31502 18398 31554 18450
rect 32174 18398 32226 18450
rect 33854 18398 33906 18450
rect 37662 18398 37714 18450
rect 38222 18398 38274 18450
rect 39678 18398 39730 18450
rect 40910 18398 40962 18450
rect 43822 18398 43874 18450
rect 44718 18398 44770 18450
rect 45950 18398 46002 18450
rect 46174 18398 46226 18450
rect 46398 18398 46450 18450
rect 46734 18398 46786 18450
rect 46846 18398 46898 18450
rect 47182 18398 47234 18450
rect 48078 18398 48130 18450
rect 3166 18286 3218 18338
rect 7198 18286 7250 18338
rect 10894 18286 10946 18338
rect 16718 18286 16770 18338
rect 19406 18286 19458 18338
rect 19742 18286 19794 18338
rect 22542 18286 22594 18338
rect 24670 18286 24722 18338
rect 26014 18286 26066 18338
rect 28142 18286 28194 18338
rect 28590 18286 28642 18338
rect 29934 18286 29986 18338
rect 34526 18286 34578 18338
rect 36654 18286 36706 18338
rect 37102 18286 37154 18338
rect 39454 18286 39506 18338
rect 40350 18286 40402 18338
rect 42030 18286 42082 18338
rect 8430 18174 8482 18226
rect 13246 18174 13298 18226
rect 18062 18174 18114 18226
rect 19182 18174 19234 18226
rect 38894 18174 38946 18226
rect 43822 18174 43874 18226
rect 44158 18174 44210 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 20638 17838 20690 17890
rect 23774 17838 23826 17890
rect 43374 17838 43426 17890
rect 46398 17838 46450 17890
rect 1934 17726 1986 17778
rect 4622 17726 4674 17778
rect 6302 17726 6354 17778
rect 11118 17726 11170 17778
rect 12910 17726 12962 17778
rect 14142 17726 14194 17778
rect 25566 17726 25618 17778
rect 27134 17726 27186 17778
rect 32958 17726 33010 17778
rect 34638 17726 34690 17778
rect 35086 17726 35138 17778
rect 38446 17726 38498 17778
rect 42926 17726 42978 17778
rect 44046 17726 44098 17778
rect 47854 17726 47906 17778
rect 2270 17614 2322 17666
rect 3726 17614 3778 17666
rect 5070 17614 5122 17666
rect 6638 17614 6690 17666
rect 8206 17614 8258 17666
rect 14926 17614 14978 17666
rect 17054 17614 17106 17666
rect 17390 17614 17442 17666
rect 19406 17614 19458 17666
rect 19630 17614 19682 17666
rect 19966 17614 20018 17666
rect 20526 17614 20578 17666
rect 21646 17614 21698 17666
rect 22430 17614 22482 17666
rect 23102 17614 23154 17666
rect 23886 17614 23938 17666
rect 24670 17614 24722 17666
rect 25006 17614 25058 17666
rect 25902 17614 25954 17666
rect 28030 17614 28082 17666
rect 28590 17614 28642 17666
rect 29150 17614 29202 17666
rect 30158 17614 30210 17666
rect 33294 17614 33346 17666
rect 33854 17614 33906 17666
rect 34526 17614 34578 17666
rect 35646 17614 35698 17666
rect 35758 17614 35810 17666
rect 35982 17614 36034 17666
rect 39006 17614 39058 17666
rect 41918 17614 41970 17666
rect 43038 17614 43090 17666
rect 43374 17614 43426 17666
rect 44718 17614 44770 17666
rect 45390 17614 45442 17666
rect 46734 17614 46786 17666
rect 3950 17502 4002 17554
rect 6302 17502 6354 17554
rect 7310 17502 7362 17554
rect 7534 17502 7586 17554
rect 7758 17502 7810 17554
rect 7870 17502 7922 17554
rect 8990 17502 9042 17554
rect 11790 17502 11842 17554
rect 12462 17502 12514 17554
rect 12574 17502 12626 17554
rect 14366 17502 14418 17554
rect 14590 17502 14642 17554
rect 14702 17502 14754 17554
rect 15374 17502 15426 17554
rect 17950 17502 18002 17554
rect 19854 17502 19906 17554
rect 21870 17502 21922 17554
rect 22206 17502 22258 17554
rect 23326 17502 23378 17554
rect 26014 17502 26066 17554
rect 27358 17502 27410 17554
rect 27694 17502 27746 17554
rect 28478 17502 28530 17554
rect 29486 17502 29538 17554
rect 30830 17502 30882 17554
rect 33406 17502 33458 17554
rect 33630 17502 33682 17554
rect 34078 17502 34130 17554
rect 34190 17502 34242 17554
rect 36094 17502 36146 17554
rect 40686 17502 40738 17554
rect 42814 17502 42866 17554
rect 45166 17502 45218 17554
rect 45614 17502 45666 17554
rect 45950 17502 46002 17554
rect 46286 17502 46338 17554
rect 46958 17502 47010 17554
rect 47070 17502 47122 17554
rect 47518 17502 47570 17554
rect 3278 17390 3330 17442
rect 3502 17390 3554 17442
rect 3614 17390 3666 17442
rect 5966 17390 6018 17442
rect 6190 17390 6242 17442
rect 7646 17390 7698 17442
rect 11454 17390 11506 17442
rect 12126 17390 12178 17442
rect 12350 17390 12402 17442
rect 13470 17390 13522 17442
rect 13806 17390 13858 17442
rect 16942 17390 16994 17442
rect 20078 17390 20130 17442
rect 20638 17390 20690 17442
rect 23774 17390 23826 17442
rect 24334 17390 24386 17442
rect 26350 17390 26402 17442
rect 26686 17390 26738 17442
rect 28254 17390 28306 17442
rect 44942 17390 44994 17442
rect 45838 17390 45890 17442
rect 46398 17390 46450 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 1710 17054 1762 17106
rect 2718 17054 2770 17106
rect 3726 17054 3778 17106
rect 3166 16942 3218 16994
rect 4062 16998 4114 17050
rect 4510 17054 4562 17106
rect 5518 17054 5570 17106
rect 10558 17054 10610 17106
rect 10782 17054 10834 17106
rect 17390 17054 17442 17106
rect 18622 17054 18674 17106
rect 22430 17054 22482 17106
rect 24334 17054 24386 17106
rect 24558 17054 24610 17106
rect 29150 17054 29202 17106
rect 29486 17054 29538 17106
rect 29822 17054 29874 17106
rect 30830 17054 30882 17106
rect 31950 17054 32002 17106
rect 32174 17054 32226 17106
rect 40238 17054 40290 17106
rect 24670 16942 24722 16994
rect 26238 16942 26290 16994
rect 27022 16942 27074 16994
rect 28366 16942 28418 16994
rect 30718 16942 30770 16994
rect 44942 16942 44994 16994
rect 47966 16942 48018 16994
rect 2270 16830 2322 16882
rect 2606 16830 2658 16882
rect 2830 16830 2882 16882
rect 4174 16830 4226 16882
rect 5854 16830 5906 16882
rect 6638 16830 6690 16882
rect 9550 16830 9602 16882
rect 9998 16830 10050 16882
rect 10446 16830 10498 16882
rect 13806 16830 13858 16882
rect 14814 16830 14866 16882
rect 17614 16830 17666 16882
rect 18062 16830 18114 16882
rect 18398 16830 18450 16882
rect 19070 16830 19122 16882
rect 20078 16830 20130 16882
rect 22542 16830 22594 16882
rect 23438 16830 23490 16882
rect 23774 16830 23826 16882
rect 25790 16830 25842 16882
rect 26574 16830 26626 16882
rect 26910 16830 26962 16882
rect 27246 16830 27298 16882
rect 28702 16830 28754 16882
rect 30942 16830 30994 16882
rect 31278 16830 31330 16882
rect 31502 16830 31554 16882
rect 32062 16830 32114 16882
rect 33070 16830 33122 16882
rect 36094 16830 36146 16882
rect 36542 16830 36594 16882
rect 40910 16830 40962 16882
rect 44158 16830 44210 16882
rect 47294 16830 47346 16882
rect 47518 16830 47570 16882
rect 47742 16830 47794 16882
rect 4958 16718 5010 16770
rect 8766 16718 8818 16770
rect 11006 16718 11058 16770
rect 13134 16718 13186 16770
rect 15374 16718 15426 16770
rect 17502 16718 17554 16770
rect 18510 16718 18562 16770
rect 18846 16718 18898 16770
rect 20974 16718 21026 16770
rect 23214 16718 23266 16770
rect 25230 16718 25282 16770
rect 27582 16718 27634 16770
rect 27694 16718 27746 16770
rect 30382 16718 30434 16770
rect 35422 16718 35474 16770
rect 37214 16718 37266 16770
rect 39342 16718 39394 16770
rect 39678 16718 39730 16770
rect 41694 16718 41746 16770
rect 43822 16718 43874 16770
rect 47070 16718 47122 16770
rect 4062 16606 4114 16658
rect 22990 16606 23042 16658
rect 27918 16606 27970 16658
rect 28030 16606 28082 16658
rect 39902 16606 39954 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 4398 16270 4450 16322
rect 12686 16270 12738 16322
rect 16494 16270 16546 16322
rect 21422 16270 21474 16322
rect 27022 16270 27074 16322
rect 2158 16158 2210 16210
rect 3166 16158 3218 16210
rect 4062 16158 4114 16210
rect 6078 16158 6130 16210
rect 7870 16158 7922 16210
rect 8318 16158 8370 16210
rect 13918 16158 13970 16210
rect 23438 16158 23490 16210
rect 23886 16158 23938 16210
rect 26686 16158 26738 16210
rect 31390 16158 31442 16210
rect 33070 16158 33122 16210
rect 36430 16158 36482 16210
rect 37102 16158 37154 16210
rect 39230 16158 39282 16210
rect 41358 16158 41410 16210
rect 41806 16158 41858 16210
rect 42702 16158 42754 16210
rect 46062 16158 46114 16210
rect 48190 16158 48242 16210
rect 5182 16046 5234 16098
rect 6750 16046 6802 16098
rect 7310 16046 7362 16098
rect 11230 16046 11282 16098
rect 11902 16046 11954 16098
rect 16046 16046 16098 16098
rect 17054 16046 17106 16098
rect 20750 16046 20802 16098
rect 23102 16046 23154 16098
rect 24222 16046 24274 16098
rect 24558 16046 24610 16098
rect 25566 16046 25618 16098
rect 27694 16046 27746 16098
rect 28254 16046 28306 16098
rect 29598 16046 29650 16098
rect 30270 16046 30322 16098
rect 30830 16046 30882 16098
rect 33630 16046 33682 16098
rect 37886 16046 37938 16098
rect 38446 16046 38498 16098
rect 42366 16046 42418 16098
rect 42926 16046 42978 16098
rect 43150 16046 43202 16098
rect 43486 16046 43538 16098
rect 43822 16046 43874 16098
rect 45390 16046 45442 16098
rect 4286 15934 4338 15986
rect 4398 15934 4450 15986
rect 4846 15934 4898 15986
rect 6302 15934 6354 15986
rect 10446 15934 10498 15986
rect 16382 15934 16434 15986
rect 16494 15934 16546 15986
rect 17614 15934 17666 15986
rect 19630 15934 19682 15986
rect 21310 15934 21362 15986
rect 21758 15934 21810 15986
rect 22094 15934 22146 15986
rect 22318 15934 22370 15986
rect 23998 15934 24050 15986
rect 24446 15934 24498 15986
rect 25230 15934 25282 15986
rect 25902 15934 25954 15986
rect 26126 15934 26178 15986
rect 26798 15934 26850 15986
rect 29374 15934 29426 15986
rect 32622 15934 32674 15986
rect 34302 15934 34354 15986
rect 37662 15934 37714 15986
rect 38110 15934 38162 15986
rect 41694 15934 41746 15986
rect 42590 15934 42642 15986
rect 43710 15934 43762 15986
rect 2718 15822 2770 15874
rect 3502 15822 3554 15874
rect 4958 15822 5010 15874
rect 5966 15822 6018 15874
rect 6190 15822 6242 15874
rect 19742 15822 19794 15874
rect 21982 15822 22034 15874
rect 24894 15822 24946 15874
rect 25790 15822 25842 15874
rect 27918 15822 27970 15874
rect 28590 15822 28642 15874
rect 30382 15822 30434 15874
rect 30494 15822 30546 15874
rect 31726 15822 31778 15874
rect 31950 15822 32002 15874
rect 32062 15822 32114 15874
rect 32174 15822 32226 15874
rect 37998 15822 38050 15874
rect 41918 15822 41970 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 2158 15486 2210 15538
rect 3502 15486 3554 15538
rect 7646 15486 7698 15538
rect 8430 15486 8482 15538
rect 12238 15486 12290 15538
rect 16270 15486 16322 15538
rect 17502 15486 17554 15538
rect 33182 15486 33234 15538
rect 33294 15486 33346 15538
rect 35310 15486 35362 15538
rect 35422 15486 35474 15538
rect 37326 15486 37378 15538
rect 37774 15486 37826 15538
rect 38222 15486 38274 15538
rect 38670 15486 38722 15538
rect 39790 15486 39842 15538
rect 39902 15486 39954 15538
rect 41134 15486 41186 15538
rect 42478 15486 42530 15538
rect 43486 15486 43538 15538
rect 43934 15486 43986 15538
rect 45054 15486 45106 15538
rect 46174 15486 46226 15538
rect 46958 15486 47010 15538
rect 47182 15486 47234 15538
rect 47742 15486 47794 15538
rect 48078 15486 48130 15538
rect 4174 15374 4226 15426
rect 4846 15374 4898 15426
rect 5518 15374 5570 15426
rect 5854 15374 5906 15426
rect 8318 15374 8370 15426
rect 17950 15374 18002 15426
rect 20526 15374 20578 15426
rect 26014 15374 26066 15426
rect 33406 15374 33458 15426
rect 39678 15374 39730 15426
rect 41246 15374 41298 15426
rect 41582 15374 41634 15426
rect 44270 15374 44322 15426
rect 45390 15374 45442 15426
rect 47406 15374 47458 15426
rect 47518 15374 47570 15426
rect 2606 15262 2658 15314
rect 3950 15262 4002 15314
rect 4622 15262 4674 15314
rect 5294 15262 5346 15314
rect 6414 15262 6466 15314
rect 6862 15262 6914 15314
rect 7982 15262 8034 15314
rect 8654 15262 8706 15314
rect 8766 15262 8818 15314
rect 9886 15262 9938 15314
rect 10334 15262 10386 15314
rect 11454 15262 11506 15314
rect 12574 15262 12626 15314
rect 15822 15262 15874 15314
rect 19070 15262 19122 15314
rect 19406 15262 19458 15314
rect 24446 15262 24498 15314
rect 25230 15262 25282 15314
rect 28590 15262 28642 15314
rect 31614 15262 31666 15314
rect 32062 15262 32114 15314
rect 32174 15262 32226 15314
rect 33966 15262 34018 15314
rect 34862 15262 34914 15314
rect 35198 15262 35250 15314
rect 36430 15262 36482 15314
rect 36878 15262 36930 15314
rect 40910 15262 40962 15314
rect 41806 15262 41858 15314
rect 42814 15262 42866 15314
rect 43150 15262 43202 15314
rect 45838 15262 45890 15314
rect 46846 15262 46898 15314
rect 47966 15262 48018 15314
rect 3166 15150 3218 15202
rect 7198 15150 7250 15202
rect 11230 15150 11282 15202
rect 11790 15150 11842 15202
rect 13022 15150 13074 15202
rect 15150 15150 15202 15202
rect 16718 15150 16770 15202
rect 21646 15150 21698 15202
rect 23774 15150 23826 15202
rect 28142 15150 28194 15202
rect 29262 15150 29314 15202
rect 31390 15150 31442 15202
rect 31838 15150 31890 15202
rect 34078 15150 34130 15202
rect 35982 15150 36034 15202
rect 42142 15150 42194 15202
rect 48078 15038 48130 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 2382 14702 2434 14754
rect 2718 14702 2770 14754
rect 13470 14702 13522 14754
rect 16494 14702 16546 14754
rect 21422 14702 21474 14754
rect 23662 14702 23714 14754
rect 28478 14702 28530 14754
rect 39790 14702 39842 14754
rect 2382 14590 2434 14642
rect 2830 14590 2882 14642
rect 3278 14590 3330 14642
rect 7870 14590 7922 14642
rect 9438 14590 9490 14642
rect 10446 14590 10498 14642
rect 11566 14590 11618 14642
rect 13582 14590 13634 14642
rect 15262 14590 15314 14642
rect 20750 14590 20802 14642
rect 22206 14590 22258 14642
rect 26574 14590 26626 14642
rect 27134 14590 27186 14642
rect 27582 14590 27634 14642
rect 28030 14590 28082 14642
rect 28590 14590 28642 14642
rect 29262 14590 29314 14642
rect 31502 14590 31554 14642
rect 33630 14590 33682 14642
rect 34078 14590 34130 14642
rect 41358 14590 41410 14642
rect 48190 14590 48242 14642
rect 5182 14478 5234 14530
rect 5518 14478 5570 14530
rect 7086 14478 7138 14530
rect 7758 14478 7810 14530
rect 8542 14478 8594 14530
rect 9102 14478 9154 14530
rect 9214 14478 9266 14530
rect 9662 14478 9714 14530
rect 9886 14478 9938 14530
rect 11118 14478 11170 14530
rect 11902 14478 11954 14530
rect 12238 14478 12290 14530
rect 12686 14478 12738 14530
rect 13806 14478 13858 14530
rect 15038 14478 15090 14530
rect 15710 14478 15762 14530
rect 16606 14478 16658 14530
rect 16942 14478 16994 14530
rect 17950 14478 18002 14530
rect 21310 14478 21362 14530
rect 22542 14478 22594 14530
rect 23886 14478 23938 14530
rect 24222 14478 24274 14530
rect 24894 14478 24946 14530
rect 25454 14478 25506 14530
rect 26126 14478 26178 14530
rect 26462 14478 26514 14530
rect 29038 14478 29090 14530
rect 29374 14478 29426 14530
rect 29710 14478 29762 14530
rect 30830 14478 30882 14530
rect 33854 14478 33906 14530
rect 34190 14478 34242 14530
rect 34526 14478 34578 14530
rect 35198 14478 35250 14530
rect 37326 14478 37378 14530
rect 38894 14478 38946 14530
rect 44158 14478 44210 14530
rect 45278 14478 45330 14530
rect 4846 14366 4898 14418
rect 4958 14366 5010 14418
rect 5966 14366 6018 14418
rect 6190 14366 6242 14418
rect 6638 14366 6690 14418
rect 8318 14366 8370 14418
rect 12798 14366 12850 14418
rect 14254 14366 14306 14418
rect 14478 14366 14530 14418
rect 14814 14366 14866 14418
rect 15486 14366 15538 14418
rect 18622 14366 18674 14418
rect 22990 14366 23042 14418
rect 23326 14366 23378 14418
rect 24110 14366 24162 14418
rect 25790 14366 25842 14418
rect 34862 14366 34914 14418
rect 35422 14366 35474 14418
rect 36318 14366 36370 14418
rect 37774 14366 37826 14418
rect 38222 14366 38274 14418
rect 39454 14366 39506 14418
rect 39678 14366 39730 14418
rect 43486 14366 43538 14418
rect 46062 14366 46114 14418
rect 1822 14254 1874 14306
rect 3614 14254 3666 14306
rect 4062 14254 4114 14306
rect 4622 14254 4674 14306
rect 5742 14254 5794 14306
rect 6526 14254 6578 14306
rect 6750 14254 6802 14306
rect 7534 14254 7586 14306
rect 7982 14254 8034 14306
rect 10782 14254 10834 14306
rect 12910 14254 12962 14306
rect 14590 14254 14642 14306
rect 16494 14254 16546 14306
rect 17278 14254 17330 14306
rect 21422 14254 21474 14306
rect 23550 14254 23602 14306
rect 25118 14254 25170 14306
rect 26686 14254 26738 14306
rect 30382 14254 30434 14306
rect 35310 14254 35362 14306
rect 35870 14254 35922 14306
rect 36990 14254 37042 14306
rect 39118 14254 39170 14306
rect 39342 14254 39394 14306
rect 40910 14254 40962 14306
rect 44942 14254 44994 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 2270 13918 2322 13970
rect 2718 13918 2770 13970
rect 6638 13918 6690 13970
rect 7086 13918 7138 13970
rect 7758 13918 7810 13970
rect 9662 13918 9714 13970
rect 15262 13918 15314 13970
rect 17726 13918 17778 13970
rect 23886 13918 23938 13970
rect 26574 13918 26626 13970
rect 28478 13918 28530 13970
rect 28814 13918 28866 13970
rect 29374 13918 29426 13970
rect 30830 13918 30882 13970
rect 31614 13918 31666 13970
rect 33630 13918 33682 13970
rect 41022 13918 41074 13970
rect 41582 13918 41634 13970
rect 43598 13918 43650 13970
rect 46958 13918 47010 13970
rect 47630 13918 47682 13970
rect 4174 13806 4226 13858
rect 8878 13806 8930 13858
rect 14926 13806 14978 13858
rect 15934 13806 15986 13858
rect 16270 13806 16322 13858
rect 16606 13806 16658 13858
rect 23662 13806 23714 13858
rect 24110 13806 24162 13858
rect 25566 13806 25618 13858
rect 45502 13806 45554 13858
rect 45838 13806 45890 13858
rect 46622 13806 46674 13858
rect 3502 13694 3554 13746
rect 6862 13694 6914 13746
rect 7422 13694 7474 13746
rect 7870 13694 7922 13746
rect 7982 13694 8034 13746
rect 8430 13694 8482 13746
rect 8542 13694 8594 13746
rect 8654 13694 8706 13746
rect 10222 13694 10274 13746
rect 10670 13694 10722 13746
rect 14366 13694 14418 13746
rect 15710 13694 15762 13746
rect 16830 13694 16882 13746
rect 17502 13694 17554 13746
rect 17950 13694 18002 13746
rect 18174 13694 18226 13746
rect 20638 13694 20690 13746
rect 21422 13694 21474 13746
rect 21534 13694 21586 13746
rect 21758 13694 21810 13746
rect 21982 13694 22034 13746
rect 23214 13694 23266 13746
rect 23438 13694 23490 13746
rect 24222 13694 24274 13746
rect 25902 13694 25954 13746
rect 26126 13694 26178 13746
rect 27470 13694 27522 13746
rect 30382 13694 30434 13746
rect 31278 13694 31330 13746
rect 33966 13694 34018 13746
rect 34190 13694 34242 13746
rect 34526 13694 34578 13746
rect 34974 13694 35026 13746
rect 38446 13694 38498 13746
rect 38670 13694 38722 13746
rect 38894 13694 38946 13746
rect 39230 13694 39282 13746
rect 39566 13694 39618 13746
rect 39790 13694 39842 13746
rect 40238 13694 40290 13746
rect 43486 13694 43538 13746
rect 43710 13694 43762 13746
rect 43934 13694 43986 13746
rect 46958 13694 47010 13746
rect 47294 13694 47346 13746
rect 47518 13694 47570 13746
rect 47854 13694 47906 13746
rect 3054 13582 3106 13634
rect 6302 13582 6354 13634
rect 6750 13582 6802 13634
rect 11342 13582 11394 13634
rect 13470 13582 13522 13634
rect 13806 13582 13858 13634
rect 16382 13582 16434 13634
rect 19406 13582 19458 13634
rect 22318 13582 22370 13634
rect 23326 13582 23378 13634
rect 24670 13582 24722 13634
rect 25678 13582 25730 13634
rect 27022 13582 27074 13634
rect 27918 13582 27970 13634
rect 29822 13582 29874 13634
rect 32062 13582 32114 13634
rect 33070 13582 33122 13634
rect 34078 13582 34130 13634
rect 35646 13582 35698 13634
rect 37774 13582 37826 13634
rect 39342 13582 39394 13634
rect 41694 13582 41746 13634
rect 9998 13470 10050 13522
rect 22542 13470 22594 13522
rect 22878 13470 22930 13522
rect 26238 13470 26290 13522
rect 27806 13470 27858 13522
rect 28030 13470 28082 13522
rect 29038 13470 29090 13522
rect 33294 13470 33346 13522
rect 38334 13470 38386 13522
rect 41806 13470 41858 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 2046 13134 2098 13186
rect 2494 13134 2546 13186
rect 3054 13134 3106 13186
rect 4622 13134 4674 13186
rect 34078 13134 34130 13186
rect 34526 13134 34578 13186
rect 2382 13022 2434 13074
rect 4622 13022 4674 13074
rect 7758 13022 7810 13074
rect 9886 13022 9938 13074
rect 11454 13022 11506 13074
rect 12126 13022 12178 13074
rect 16718 13022 16770 13074
rect 20750 13022 20802 13074
rect 27358 13022 27410 13074
rect 28142 13022 28194 13074
rect 29934 13022 29986 13074
rect 32062 13022 32114 13074
rect 32622 13022 32674 13074
rect 33518 13022 33570 13074
rect 35870 13022 35922 13074
rect 38558 13022 38610 13074
rect 40686 13022 40738 13074
rect 41022 13022 41074 13074
rect 43150 13022 43202 13074
rect 5966 12910 6018 12962
rect 6414 12910 6466 12962
rect 6638 12910 6690 12962
rect 7086 12910 7138 12962
rect 10334 12910 10386 12962
rect 10558 12910 10610 12962
rect 10782 12910 10834 12962
rect 11790 12910 11842 12962
rect 12238 12910 12290 12962
rect 13918 12910 13970 12962
rect 17054 12910 17106 12962
rect 17390 12910 17442 12962
rect 17838 12910 17890 12962
rect 18622 12910 18674 12962
rect 22430 12910 22482 12962
rect 22766 12910 22818 12962
rect 23438 12910 23490 12962
rect 23774 12910 23826 12962
rect 24558 12910 24610 12962
rect 25230 12910 25282 12962
rect 28030 12910 28082 12962
rect 28366 12910 28418 12962
rect 29150 12910 29202 12962
rect 33406 12910 33458 12962
rect 33742 12910 33794 12962
rect 34190 12910 34242 12962
rect 34414 12910 34466 12962
rect 35086 12910 35138 12962
rect 35534 12910 35586 12962
rect 36206 12910 36258 12962
rect 37886 12910 37938 12962
rect 43822 12910 43874 12962
rect 46510 12910 46562 12962
rect 46846 12910 46898 12962
rect 47182 12910 47234 12962
rect 12014 12798 12066 12850
rect 12574 12798 12626 12850
rect 14590 12798 14642 12850
rect 17166 12798 17218 12850
rect 21646 12798 21698 12850
rect 21758 12798 21810 12850
rect 21982 12798 22034 12850
rect 22206 12798 22258 12850
rect 23102 12798 23154 12850
rect 23550 12798 23602 12850
rect 28590 12798 28642 12850
rect 33182 12798 33234 12850
rect 34862 12798 34914 12850
rect 46062 12798 46114 12850
rect 47854 12798 47906 12850
rect 1934 12686 1986 12738
rect 2830 12686 2882 12738
rect 3278 12686 3330 12738
rect 3726 12686 3778 12738
rect 4174 12686 4226 12738
rect 5070 12686 5122 12738
rect 5742 12686 5794 12738
rect 6190 12686 6242 12738
rect 10558 12686 10610 12738
rect 11230 12686 11282 12738
rect 11454 12686 11506 12738
rect 22654 12686 22706 12738
rect 24110 12686 24162 12738
rect 35310 12686 35362 12738
rect 37102 12686 37154 12738
rect 44830 12686 44882 12738
rect 45166 12686 45218 12738
rect 45726 12686 45778 12738
rect 45950 12686 46002 12738
rect 46846 12686 46898 12738
rect 47630 12686 47682 12738
rect 48190 12686 48242 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 1934 12350 1986 12402
rect 6750 12350 6802 12402
rect 7646 12350 7698 12402
rect 7982 12350 8034 12402
rect 9550 12350 9602 12402
rect 10334 12350 10386 12402
rect 10670 12350 10722 12402
rect 10894 12350 10946 12402
rect 11678 12350 11730 12402
rect 12126 12350 12178 12402
rect 13022 12350 13074 12402
rect 14030 12350 14082 12402
rect 14254 12350 14306 12402
rect 14590 12350 14642 12402
rect 15150 12350 15202 12402
rect 16270 12350 16322 12402
rect 16494 12350 16546 12402
rect 16718 12350 16770 12402
rect 17838 12350 17890 12402
rect 18510 12350 18562 12402
rect 18622 12350 18674 12402
rect 18734 12350 18786 12402
rect 19854 12350 19906 12402
rect 19966 12350 20018 12402
rect 20302 12350 20354 12402
rect 20414 12350 20466 12402
rect 21310 12350 21362 12402
rect 21534 12350 21586 12402
rect 25342 12350 25394 12402
rect 26350 12350 26402 12402
rect 26462 12350 26514 12402
rect 26574 12350 26626 12402
rect 27806 12350 27858 12402
rect 28478 12350 28530 12402
rect 28590 12350 28642 12402
rect 28702 12350 28754 12402
rect 29374 12350 29426 12402
rect 31614 12350 31666 12402
rect 34078 12350 34130 12402
rect 34414 12350 34466 12402
rect 36654 12350 36706 12402
rect 40350 12350 40402 12402
rect 42814 12350 42866 12402
rect 44158 12350 44210 12402
rect 44942 12350 44994 12402
rect 3838 12238 3890 12290
rect 8654 12238 8706 12290
rect 10110 12238 10162 12290
rect 12574 12238 12626 12290
rect 13918 12238 13970 12290
rect 14478 12238 14530 12290
rect 16382 12238 16434 12290
rect 18174 12238 18226 12290
rect 21198 12238 21250 12290
rect 22542 12238 22594 12290
rect 26014 12238 26066 12290
rect 27582 12238 27634 12290
rect 29822 12238 29874 12290
rect 31278 12238 31330 12290
rect 31390 12238 31442 12290
rect 31838 12238 31890 12290
rect 32062 12238 32114 12290
rect 32174 12238 32226 12290
rect 39006 12238 39058 12290
rect 41918 12238 41970 12290
rect 46062 12238 46114 12290
rect 3054 12126 3106 12178
rect 6974 12126 7026 12178
rect 7310 12126 7362 12178
rect 8990 12126 9042 12178
rect 9886 12126 9938 12178
rect 10446 12126 10498 12178
rect 11006 12126 11058 12178
rect 11566 12126 11618 12178
rect 11902 12126 11954 12178
rect 12350 12126 12402 12178
rect 15038 12126 15090 12178
rect 15374 12126 15426 12178
rect 15598 12126 15650 12178
rect 17614 12126 17666 12178
rect 17838 12126 17890 12178
rect 19182 12126 19234 12178
rect 19294 12126 19346 12178
rect 19742 12126 19794 12178
rect 20526 12126 20578 12178
rect 20974 12126 21026 12178
rect 21870 12126 21922 12178
rect 25678 12126 25730 12178
rect 27022 12126 27074 12178
rect 27918 12126 27970 12178
rect 28142 12126 28194 12178
rect 29038 12126 29090 12178
rect 29486 12126 29538 12178
rect 29598 12126 29650 12178
rect 30830 12126 30882 12178
rect 33070 12126 33122 12178
rect 34750 12126 34802 12178
rect 34862 12126 34914 12178
rect 34974 12126 35026 12178
rect 35422 12126 35474 12178
rect 35534 12126 35586 12178
rect 35870 12126 35922 12178
rect 36094 12126 36146 12178
rect 36318 12126 36370 12178
rect 36542 12126 36594 12178
rect 39790 12126 39842 12178
rect 41246 12126 41298 12178
rect 45278 12126 45330 12178
rect 2270 12014 2322 12066
rect 2830 12014 2882 12066
rect 5966 12014 6018 12066
rect 6414 12014 6466 12066
rect 6862 12014 6914 12066
rect 24670 12014 24722 12066
rect 30494 12014 30546 12066
rect 31502 12014 31554 12066
rect 36878 12014 36930 12066
rect 41134 12014 41186 12066
rect 42366 12014 42418 12066
rect 48190 12014 48242 12066
rect 13022 11902 13074 11954
rect 13134 11902 13186 11954
rect 13358 11902 13410 11954
rect 14590 11902 14642 11954
rect 33294 11902 33346 11954
rect 33630 11902 33682 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 7758 11566 7810 11618
rect 22206 11566 22258 11618
rect 23102 11566 23154 11618
rect 34078 11566 34130 11618
rect 34862 11566 34914 11618
rect 37438 11566 37490 11618
rect 46398 11566 46450 11618
rect 1822 11454 1874 11506
rect 5070 11454 5122 11506
rect 7534 11454 7586 11506
rect 12462 11454 12514 11506
rect 14366 11454 14418 11506
rect 16494 11454 16546 11506
rect 20526 11454 20578 11506
rect 21310 11454 21362 11506
rect 21534 11454 21586 11506
rect 22542 11454 22594 11506
rect 23886 11454 23938 11506
rect 24446 11454 24498 11506
rect 24782 11454 24834 11506
rect 25902 11454 25954 11506
rect 26350 11454 26402 11506
rect 31614 11454 31666 11506
rect 33742 11454 33794 11506
rect 35870 11454 35922 11506
rect 37102 11454 37154 11506
rect 37550 11454 37602 11506
rect 39006 11454 39058 11506
rect 40574 11454 40626 11506
rect 41470 11454 41522 11506
rect 43038 11454 43090 11506
rect 43486 11454 43538 11506
rect 2270 11342 2322 11394
rect 5630 11342 5682 11394
rect 6302 11342 6354 11394
rect 6750 11342 6802 11394
rect 8094 11342 8146 11394
rect 8990 11342 9042 11394
rect 9438 11342 9490 11394
rect 9662 11342 9714 11394
rect 9886 11342 9938 11394
rect 10670 11342 10722 11394
rect 11118 11342 11170 11394
rect 12238 11342 12290 11394
rect 13582 11342 13634 11394
rect 17614 11342 17666 11394
rect 18398 11342 18450 11394
rect 22318 11342 22370 11394
rect 22766 11342 22818 11394
rect 25342 11342 25394 11394
rect 26798 11342 26850 11394
rect 27470 11342 27522 11394
rect 29710 11342 29762 11394
rect 30942 11342 30994 11394
rect 34526 11342 34578 11394
rect 35086 11342 35138 11394
rect 35534 11342 35586 11394
rect 35758 11342 35810 11394
rect 37998 11342 38050 11394
rect 40238 11342 40290 11394
rect 41134 11342 41186 11394
rect 42030 11342 42082 11394
rect 42366 11342 42418 11394
rect 45390 11342 45442 11394
rect 45726 11342 45778 11394
rect 45838 11342 45890 11394
rect 46510 11342 46562 11394
rect 47182 11342 47234 11394
rect 47630 11342 47682 11394
rect 2942 11230 2994 11282
rect 6078 11230 6130 11282
rect 7086 11230 7138 11282
rect 8542 11230 8594 11282
rect 11230 11230 11282 11282
rect 11790 11230 11842 11282
rect 12014 11230 12066 11282
rect 12686 11230 12738 11282
rect 16830 11230 16882 11282
rect 17166 11230 17218 11282
rect 23326 11230 23378 11282
rect 25118 11230 25170 11282
rect 34190 11230 34242 11282
rect 44830 11230 44882 11282
rect 44942 11230 44994 11282
rect 46398 11230 46450 11282
rect 46846 11230 46898 11282
rect 47518 11230 47570 11282
rect 5854 11118 5906 11170
rect 6638 11118 6690 11170
rect 6862 11118 6914 11170
rect 8766 11118 8818 11170
rect 8878 11118 8930 11170
rect 11342 11118 11394 11170
rect 12126 11118 12178 11170
rect 21870 11118 21922 11170
rect 23214 11118 23266 11170
rect 26910 11118 26962 11170
rect 27022 11118 27074 11170
rect 27806 11118 27858 11170
rect 28254 11118 28306 11170
rect 29262 11118 29314 11170
rect 30494 11118 30546 11170
rect 34750 11118 34802 11170
rect 38446 11118 38498 11170
rect 42478 11118 42530 11170
rect 42702 11118 42754 11170
rect 45166 11118 45218 11170
rect 45502 11118 45554 11170
rect 46958 11118 47010 11170
rect 47294 11118 47346 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 3054 10782 3106 10834
rect 3502 10782 3554 10834
rect 7198 10782 7250 10834
rect 8094 10782 8146 10834
rect 8654 10782 8706 10834
rect 14030 10782 14082 10834
rect 15038 10782 15090 10834
rect 16046 10782 16098 10834
rect 16270 10782 16322 10834
rect 17726 10782 17778 10834
rect 18174 10782 18226 10834
rect 20414 10782 20466 10834
rect 32398 10782 32450 10834
rect 34862 10782 34914 10834
rect 35534 10782 35586 10834
rect 36990 10782 37042 10834
rect 40014 10782 40066 10834
rect 46958 10782 47010 10834
rect 4510 10670 4562 10722
rect 6974 10670 7026 10722
rect 11902 10670 11954 10722
rect 13246 10670 13298 10722
rect 13358 10670 13410 10722
rect 13806 10670 13858 10722
rect 14254 10670 14306 10722
rect 14926 10670 14978 10722
rect 15486 10670 15538 10722
rect 18958 10670 19010 10722
rect 19854 10670 19906 10722
rect 20750 10670 20802 10722
rect 23326 10670 23378 10722
rect 26126 10670 26178 10722
rect 26462 10670 26514 10722
rect 26686 10670 26738 10722
rect 28030 10670 28082 10722
rect 30606 10670 30658 10722
rect 34190 10670 34242 10722
rect 34302 10670 34354 10722
rect 35310 10670 35362 10722
rect 36206 10670 36258 10722
rect 37550 10670 37602 10722
rect 38894 10670 38946 10722
rect 41022 10670 41074 10722
rect 43150 10670 43202 10722
rect 46510 10670 46562 10722
rect 47182 10670 47234 10722
rect 47294 10670 47346 10722
rect 3838 10558 3890 10610
rect 7310 10558 7362 10610
rect 7422 10558 7474 10610
rect 12686 10558 12738 10610
rect 13694 10558 13746 10610
rect 14478 10558 14530 10610
rect 15262 10558 15314 10610
rect 16382 10558 16434 10610
rect 16494 10558 16546 10610
rect 16942 10558 16994 10610
rect 17838 10558 17890 10610
rect 17950 10558 18002 10610
rect 18510 10558 18562 10610
rect 19182 10558 19234 10610
rect 19518 10558 19570 10610
rect 20974 10558 21026 10610
rect 21086 10558 21138 10610
rect 21198 10558 21250 10610
rect 21870 10558 21922 10610
rect 22094 10558 22146 10610
rect 22990 10558 23042 10610
rect 23774 10558 23826 10610
rect 23998 10558 24050 10610
rect 25678 10558 25730 10610
rect 27358 10558 27410 10610
rect 30830 10558 30882 10610
rect 31166 10558 31218 10610
rect 34526 10558 34578 10610
rect 35646 10558 35698 10610
rect 35870 10558 35922 10610
rect 36542 10558 36594 10610
rect 37998 10558 38050 10610
rect 39230 10558 39282 10610
rect 39678 10558 39730 10610
rect 40014 10558 40066 10610
rect 40350 10558 40402 10610
rect 40910 10558 40962 10610
rect 41806 10558 41858 10610
rect 42478 10558 42530 10610
rect 46062 10558 46114 10610
rect 46734 10558 46786 10610
rect 2158 10446 2210 10498
rect 2494 10446 2546 10498
rect 6638 10446 6690 10498
rect 9102 10446 9154 10498
rect 9774 10446 9826 10498
rect 18734 10446 18786 10498
rect 21982 10446 22034 10498
rect 23886 10446 23938 10498
rect 24446 10446 24498 10498
rect 25230 10446 25282 10498
rect 26238 10446 26290 10498
rect 30158 10446 30210 10498
rect 30718 10446 30770 10498
rect 31950 10446 32002 10498
rect 33182 10446 33234 10498
rect 33630 10446 33682 10498
rect 41022 10446 41074 10498
rect 45278 10446 45330 10498
rect 46286 10446 46338 10498
rect 21646 10334 21698 10386
rect 21870 10334 21922 10386
rect 22542 10334 22594 10386
rect 23550 10334 23602 10386
rect 37774 10334 37826 10386
rect 38222 10334 38274 10386
rect 38670 10334 38722 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 2942 9998 2994 10050
rect 3614 9998 3666 10050
rect 10222 9998 10274 10050
rect 11566 9998 11618 10050
rect 12798 9998 12850 10050
rect 42814 9998 42866 10050
rect 2942 9886 2994 9938
rect 4622 9886 4674 9938
rect 6190 9886 6242 9938
rect 10110 9886 10162 9938
rect 11006 9886 11058 9938
rect 12014 9886 12066 9938
rect 12574 9886 12626 9938
rect 12910 9886 12962 9938
rect 15374 9886 15426 9938
rect 16382 9886 16434 9938
rect 18510 9886 18562 9938
rect 19070 9886 19122 9938
rect 21646 9886 21698 9938
rect 23774 9886 23826 9938
rect 25678 9886 25730 9938
rect 27806 9886 27858 9938
rect 32062 9886 32114 9938
rect 35310 9886 35362 9938
rect 46062 9886 46114 9938
rect 48190 9886 48242 9938
rect 3838 9774 3890 9826
rect 7870 9774 7922 9826
rect 8206 9774 8258 9826
rect 8542 9774 8594 9826
rect 9326 9774 9378 9826
rect 11678 9774 11730 9826
rect 15710 9774 15762 9826
rect 24558 9774 24610 9826
rect 24894 9774 24946 9826
rect 28254 9774 28306 9826
rect 29262 9774 29314 9826
rect 32510 9774 32562 9826
rect 36094 9774 36146 9826
rect 36990 9774 37042 9826
rect 37214 9774 37266 9826
rect 37998 9774 38050 9826
rect 40014 9774 40066 9826
rect 42142 9774 42194 9826
rect 42366 9774 42418 9826
rect 43038 9774 43090 9826
rect 43262 9774 43314 9826
rect 44046 9774 44098 9826
rect 45278 9774 45330 9826
rect 2046 9662 2098 9714
rect 7310 9662 7362 9714
rect 7534 9662 7586 9714
rect 13806 9662 13858 9714
rect 14814 9662 14866 9714
rect 20750 9662 20802 9714
rect 29934 9662 29986 9714
rect 33182 9662 33234 9714
rect 37550 9662 37602 9714
rect 39566 9662 39618 9714
rect 41022 9662 41074 9714
rect 43486 9662 43538 9714
rect 44270 9662 44322 9714
rect 2382 9550 2434 9602
rect 3390 9550 3442 9602
rect 4286 9550 4338 9602
rect 5070 9550 5122 9602
rect 6638 9550 6690 9602
rect 6974 9550 7026 9602
rect 7646 9550 7698 9602
rect 8318 9550 8370 9602
rect 8990 9550 9042 9602
rect 9214 9550 9266 9602
rect 10446 9550 10498 9602
rect 13918 9550 13970 9602
rect 14142 9550 14194 9602
rect 19406 9550 19458 9602
rect 19854 9550 19906 9602
rect 20190 9550 20242 9602
rect 28478 9550 28530 9602
rect 35758 9550 35810 9602
rect 36430 9550 36482 9602
rect 37102 9550 37154 9602
rect 39678 9550 39730 9602
rect 44942 9550 44994 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 2942 9214 2994 9266
rect 3390 9214 3442 9266
rect 7310 9214 7362 9266
rect 9662 9214 9714 9266
rect 10446 9214 10498 9266
rect 16046 9214 16098 9266
rect 17726 9214 17778 9266
rect 18286 9214 18338 9266
rect 23326 9214 23378 9266
rect 24558 9214 24610 9266
rect 25454 9214 25506 9266
rect 26014 9214 26066 9266
rect 26462 9214 26514 9266
rect 27806 9214 27858 9266
rect 28142 9214 28194 9266
rect 28590 9214 28642 9266
rect 29710 9214 29762 9266
rect 30830 9214 30882 9266
rect 32062 9214 32114 9266
rect 36654 9214 36706 9266
rect 37102 9214 37154 9266
rect 37886 9214 37938 9266
rect 38782 9214 38834 9266
rect 40014 9214 40066 9266
rect 44942 9214 44994 9266
rect 46734 9214 46786 9266
rect 47406 9214 47458 9266
rect 7534 9102 7586 9154
rect 8430 9102 8482 9154
rect 14254 9102 14306 9154
rect 15038 9102 15090 9154
rect 16942 9102 16994 9154
rect 17390 9102 17442 9154
rect 22094 9102 22146 9154
rect 23214 9102 23266 9154
rect 27246 9102 27298 9154
rect 29150 9102 29202 9154
rect 29486 9102 29538 9154
rect 29822 9102 29874 9154
rect 30046 9102 30098 9154
rect 30606 9102 30658 9154
rect 31166 9102 31218 9154
rect 31950 9102 32002 9154
rect 37662 9102 37714 9154
rect 38558 9102 38610 9154
rect 38894 9102 38946 9154
rect 39118 9102 39170 9154
rect 40126 9102 40178 9154
rect 40910 9102 40962 9154
rect 41022 9102 41074 9154
rect 45278 9102 45330 9154
rect 46398 9102 46450 9154
rect 47294 9102 47346 9154
rect 2046 8990 2098 9042
rect 3726 8990 3778 9042
rect 7982 8990 8034 9042
rect 8206 8990 8258 9042
rect 8878 8990 8930 9042
rect 9998 8990 10050 9042
rect 13582 8990 13634 9042
rect 14030 8990 14082 9042
rect 14702 8990 14754 9042
rect 14926 8990 14978 9042
rect 15262 8990 15314 9042
rect 18622 8990 18674 9042
rect 21758 8990 21810 9042
rect 22206 8990 22258 9042
rect 27022 8990 27074 9042
rect 30830 8990 30882 9042
rect 31390 8990 31442 9042
rect 31838 8990 31890 9042
rect 36094 8990 36146 9042
rect 37886 8990 37938 9042
rect 38222 8990 38274 9042
rect 39678 8990 39730 9042
rect 40350 8990 40402 9042
rect 41246 8990 41298 9042
rect 44494 8990 44546 9042
rect 46622 8990 46674 9042
rect 47070 8990 47122 9042
rect 47854 8990 47906 9042
rect 2494 8878 2546 8930
rect 4398 8878 4450 8930
rect 6526 8878 6578 8930
rect 7422 8878 7474 8930
rect 7870 8878 7922 8930
rect 10782 8878 10834 8930
rect 12910 8878 12962 8930
rect 14478 8878 14530 8930
rect 16494 8878 16546 8930
rect 19294 8878 19346 8930
rect 21422 8878 21474 8930
rect 21870 8878 21922 8930
rect 22766 8878 22818 8930
rect 23886 8878 23938 8930
rect 32510 8878 32562 8930
rect 33294 8878 33346 8930
rect 35422 8878 35474 8930
rect 41694 8878 41746 8930
rect 43822 8878 43874 8930
rect 45726 8878 45778 8930
rect 47966 8878 48018 8930
rect 2494 8766 2546 8818
rect 2718 8766 2770 8818
rect 3278 8766 3330 8818
rect 8766 8766 8818 8818
rect 15822 8766 15874 8818
rect 16494 8766 16546 8818
rect 23886 8766 23938 8818
rect 24670 8766 24722 8818
rect 27918 8766 27970 8818
rect 28478 8766 28530 8818
rect 47406 8766 47458 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 4846 8430 4898 8482
rect 7422 8430 7474 8482
rect 8878 8430 8930 8482
rect 36318 8430 36370 8482
rect 1934 8318 1986 8370
rect 3278 8318 3330 8370
rect 4174 8318 4226 8370
rect 4958 8318 5010 8370
rect 3726 8206 3778 8258
rect 2382 8094 2434 8146
rect 5742 8094 5794 8146
rect 5854 8094 5906 8146
rect 6414 8318 6466 8370
rect 8654 8318 8706 8370
rect 12798 8318 12850 8370
rect 13470 8318 13522 8370
rect 19182 8318 19234 8370
rect 22654 8318 22706 8370
rect 28590 8318 28642 8370
rect 32062 8318 32114 8370
rect 32510 8318 32562 8370
rect 37102 8318 37154 8370
rect 46062 8318 46114 8370
rect 48190 8318 48242 8370
rect 6414 8206 6466 8258
rect 6862 8206 6914 8258
rect 7310 8206 7362 8258
rect 7982 8206 8034 8258
rect 8206 8206 8258 8258
rect 9102 8206 9154 8258
rect 9326 8206 9378 8258
rect 10670 8206 10722 8258
rect 12014 8206 12066 8258
rect 12350 8206 12402 8258
rect 16270 8206 16322 8258
rect 17502 8206 17554 8258
rect 18174 8206 18226 8258
rect 19518 8206 19570 8258
rect 19854 8206 19906 8258
rect 20190 8206 20242 8258
rect 21534 8206 21586 8258
rect 23662 8206 23714 8258
rect 25902 8206 25954 8258
rect 27806 8206 27858 8258
rect 33854 8206 33906 8258
rect 34526 8206 34578 8258
rect 34750 8206 34802 8258
rect 35870 8206 35922 8258
rect 36206 8206 36258 8258
rect 37774 8206 37826 8258
rect 37998 8206 38050 8258
rect 38894 8206 38946 8258
rect 39566 8206 39618 8258
rect 39790 8206 39842 8258
rect 40910 8206 40962 8258
rect 41022 8206 41074 8258
rect 41918 8206 41970 8258
rect 42142 8206 42194 8258
rect 42590 8206 42642 8258
rect 42814 8206 42866 8258
rect 43822 8206 43874 8258
rect 44158 8206 44210 8258
rect 45390 8206 45442 8258
rect 8094 8094 8146 8146
rect 10446 8094 10498 8146
rect 12798 8094 12850 8146
rect 15598 8094 15650 8146
rect 16830 8094 16882 8146
rect 17054 8094 17106 8146
rect 18510 8094 18562 8146
rect 18846 8094 18898 8146
rect 19070 8094 19122 8146
rect 20414 8094 20466 8146
rect 21422 8094 21474 8146
rect 23774 8094 23826 8146
rect 26350 8094 26402 8146
rect 29486 8094 29538 8146
rect 29598 8094 29650 8146
rect 30382 8094 30434 8146
rect 31278 8094 31330 8146
rect 34190 8094 34242 8146
rect 35086 8094 35138 8146
rect 35422 8094 35474 8146
rect 35758 8094 35810 8146
rect 41358 8094 41410 8146
rect 41582 8094 41634 8146
rect 43150 8094 43202 8146
rect 2830 7982 2882 8034
rect 4622 7982 4674 8034
rect 5630 7982 5682 8034
rect 6750 7982 6802 8034
rect 6974 7982 7026 8034
rect 7758 7982 7810 8034
rect 9774 7982 9826 8034
rect 10222 7982 10274 8034
rect 11118 7982 11170 8034
rect 11454 7982 11506 8034
rect 16718 7982 16770 8034
rect 16942 7982 16994 8034
rect 17838 7982 17890 8034
rect 18622 7982 18674 8034
rect 19630 7982 19682 8034
rect 21198 7982 21250 8034
rect 21982 7982 22034 8034
rect 22990 7982 23042 8034
rect 23326 7982 23378 8034
rect 26462 7982 26514 8034
rect 28142 7982 28194 8034
rect 29150 7982 29202 8034
rect 29262 7982 29314 8034
rect 29374 7982 29426 8034
rect 30270 7982 30322 8034
rect 30830 7982 30882 8034
rect 32958 7982 33010 8034
rect 33294 7982 33346 8034
rect 34414 7982 34466 8034
rect 35198 7982 35250 8034
rect 35534 7982 35586 8034
rect 36318 7982 36370 8034
rect 37438 7982 37490 8034
rect 38446 7982 38498 8034
rect 38670 7982 38722 8034
rect 38782 7982 38834 8034
rect 39230 7982 39282 8034
rect 40238 7982 40290 8034
rect 41694 7982 41746 8034
rect 42478 7982 42530 8034
rect 43262 7982 43314 8034
rect 43374 7982 43426 8034
rect 44942 7982 44994 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 1822 7646 1874 7698
rect 6974 7646 7026 7698
rect 8094 7646 8146 7698
rect 8654 7646 8706 7698
rect 9102 7646 9154 7698
rect 9998 7646 10050 7698
rect 10334 7646 10386 7698
rect 10894 7646 10946 7698
rect 15150 7646 15202 7698
rect 15934 7646 15986 7698
rect 16382 7646 16434 7698
rect 16942 7646 16994 7698
rect 18846 7646 18898 7698
rect 19294 7646 19346 7698
rect 19854 7646 19906 7698
rect 23102 7646 23154 7698
rect 23438 7646 23490 7698
rect 23886 7646 23938 7698
rect 27582 7646 27634 7698
rect 27806 7646 27858 7698
rect 32286 7646 32338 7698
rect 33742 7646 33794 7698
rect 35870 7646 35922 7698
rect 38894 7646 38946 7698
rect 40126 7646 40178 7698
rect 40238 7646 40290 7698
rect 40350 7646 40402 7698
rect 41470 7646 41522 7698
rect 42814 7646 42866 7698
rect 43822 7646 43874 7698
rect 44270 7646 44322 7698
rect 45054 7646 45106 7698
rect 45614 7646 45666 7698
rect 46622 7646 46674 7698
rect 46846 7646 46898 7698
rect 47406 7646 47458 7698
rect 47854 7646 47906 7698
rect 4174 7534 4226 7586
rect 6638 7534 6690 7586
rect 10782 7534 10834 7586
rect 13806 7534 13858 7586
rect 14814 7534 14866 7586
rect 15822 7534 15874 7586
rect 20638 7534 20690 7586
rect 21086 7534 21138 7586
rect 21982 7534 22034 7586
rect 24222 7534 24274 7586
rect 25790 7534 25842 7586
rect 26574 7534 26626 7586
rect 27470 7534 27522 7586
rect 28814 7534 28866 7586
rect 31390 7534 31442 7586
rect 33070 7534 33122 7586
rect 33406 7534 33458 7586
rect 34750 7534 34802 7586
rect 35198 7534 35250 7586
rect 36766 7534 36818 7586
rect 37214 7534 37266 7586
rect 39118 7534 39170 7586
rect 41246 7534 41298 7586
rect 44606 7534 44658 7586
rect 48190 7534 48242 7586
rect 3502 7422 3554 7474
rect 6974 7422 7026 7474
rect 7310 7422 7362 7474
rect 7534 7422 7586 7474
rect 7758 7422 7810 7474
rect 12238 7422 12290 7474
rect 14366 7422 14418 7474
rect 17278 7422 17330 7474
rect 17726 7422 17778 7474
rect 17838 7422 17890 7474
rect 19630 7422 19682 7474
rect 20302 7422 20354 7474
rect 20974 7422 21026 7474
rect 21198 7422 21250 7474
rect 22206 7422 22258 7474
rect 24558 7422 24610 7474
rect 25566 7422 25618 7474
rect 26910 7422 26962 7474
rect 27134 7422 27186 7474
rect 28030 7422 28082 7474
rect 31278 7422 31330 7474
rect 32174 7422 32226 7474
rect 35534 7422 35586 7474
rect 36206 7422 36258 7474
rect 36990 7422 37042 7474
rect 38110 7422 38162 7474
rect 38670 7422 38722 7474
rect 39678 7422 39730 7474
rect 40910 7422 40962 7474
rect 41134 7422 41186 7474
rect 41806 7422 41858 7474
rect 41918 7422 41970 7474
rect 42254 7422 42306 7474
rect 42478 7422 42530 7474
rect 43710 7422 43762 7474
rect 44046 7422 44098 7474
rect 45166 7422 45218 7474
rect 46958 7422 47010 7474
rect 47294 7422 47346 7474
rect 2718 7310 2770 7362
rect 3166 7310 3218 7362
rect 6302 7310 6354 7362
rect 9774 7310 9826 7362
rect 17502 7310 17554 7362
rect 18510 7310 18562 7362
rect 26350 7310 26402 7362
rect 26686 7310 26738 7362
rect 30942 7310 30994 7362
rect 34302 7310 34354 7362
rect 36430 7310 36482 7362
rect 36878 7310 36930 7362
rect 38334 7310 38386 7362
rect 38782 7310 38834 7362
rect 43262 7310 43314 7362
rect 16158 7198 16210 7250
rect 16718 7198 16770 7250
rect 19966 7198 20018 7250
rect 20414 7198 20466 7250
rect 22430 7198 22482 7250
rect 22654 7198 22706 7250
rect 35534 7198 35586 7250
rect 37774 7198 37826 7250
rect 45054 7198 45106 7250
rect 47406 7198 47458 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 2830 6862 2882 6914
rect 3502 6862 3554 6914
rect 4622 6862 4674 6914
rect 11454 6862 11506 6914
rect 11678 6862 11730 6914
rect 35310 6862 35362 6914
rect 38110 6862 38162 6914
rect 38222 6862 38274 6914
rect 39454 6862 39506 6914
rect 39566 6862 39618 6914
rect 2830 6750 2882 6802
rect 4622 6750 4674 6802
rect 8430 6750 8482 6802
rect 13022 6750 13074 6802
rect 14142 6750 14194 6802
rect 17838 6750 17890 6802
rect 27022 6750 27074 6802
rect 27470 6750 27522 6802
rect 28366 6750 28418 6802
rect 32398 6750 32450 6802
rect 34862 6750 34914 6802
rect 39118 6750 39170 6802
rect 44270 6750 44322 6802
rect 48302 6750 48354 6802
rect 3838 6638 3890 6690
rect 5854 6638 5906 6690
rect 6750 6638 6802 6690
rect 6974 6638 7026 6690
rect 7422 6638 7474 6690
rect 8990 6638 9042 6690
rect 9214 6638 9266 6690
rect 9550 6638 9602 6690
rect 9662 6638 9714 6690
rect 10446 6638 10498 6690
rect 10670 6638 10722 6690
rect 11230 6638 11282 6690
rect 12126 6638 12178 6690
rect 13694 6638 13746 6690
rect 16270 6638 16322 6690
rect 17054 6638 17106 6690
rect 17950 6638 18002 6690
rect 18174 6638 18226 6690
rect 19518 6638 19570 6690
rect 19854 6638 19906 6690
rect 20078 6638 20130 6690
rect 21534 6638 21586 6690
rect 21870 6638 21922 6690
rect 22094 6638 22146 6690
rect 23550 6638 23602 6690
rect 24222 6638 24274 6690
rect 24894 6638 24946 6690
rect 27358 6638 27410 6690
rect 29934 6638 29986 6690
rect 30270 6638 30322 6690
rect 31278 6638 31330 6690
rect 31502 6638 31554 6690
rect 32174 6638 32226 6690
rect 32734 6638 32786 6690
rect 33070 6638 33122 6690
rect 33294 6638 33346 6690
rect 33630 6638 33682 6690
rect 34302 6638 34354 6690
rect 35422 6638 35474 6690
rect 36318 6638 36370 6690
rect 37102 6638 37154 6690
rect 38782 6638 38834 6690
rect 40126 6638 40178 6690
rect 40350 6638 40402 6690
rect 41358 6638 41410 6690
rect 44718 6638 44770 6690
rect 45054 6638 45106 6690
rect 46958 6638 47010 6690
rect 47294 6638 47346 6690
rect 47854 6638 47906 6690
rect 3390 6526 3442 6578
rect 4286 6526 4338 6578
rect 11006 6526 11058 6578
rect 12574 6526 12626 6578
rect 17502 6526 17554 6578
rect 18622 6526 18674 6578
rect 18846 6526 18898 6578
rect 22430 6526 22482 6578
rect 27582 6526 27634 6578
rect 27806 6526 27858 6578
rect 30606 6526 30658 6578
rect 30830 6526 30882 6578
rect 35758 6526 35810 6578
rect 35982 6526 36034 6578
rect 37774 6526 37826 6578
rect 38558 6526 38610 6578
rect 39006 6526 39058 6578
rect 39790 6526 39842 6578
rect 42142 6526 42194 6578
rect 44942 6526 44994 6578
rect 45390 6526 45442 6578
rect 46062 6526 46114 6578
rect 46622 6526 46674 6578
rect 47518 6526 47570 6578
rect 5182 6414 5234 6466
rect 6190 6414 6242 6466
rect 6302 6414 6354 6466
rect 6414 6414 6466 6466
rect 7086 6414 7138 6466
rect 8094 6414 8146 6466
rect 8318 6414 8370 6466
rect 8542 6414 8594 6466
rect 9326 6414 9378 6466
rect 10110 6414 10162 6466
rect 13470 6414 13522 6466
rect 17726 6414 17778 6466
rect 18398 6414 18450 6466
rect 19966 6414 20018 6466
rect 20414 6414 20466 6466
rect 20750 6414 20802 6466
rect 22094 6414 22146 6466
rect 22990 6414 23042 6466
rect 23774 6414 23826 6466
rect 29486 6414 29538 6466
rect 30494 6414 30546 6466
rect 31838 6414 31890 6466
rect 33182 6414 33234 6466
rect 34078 6414 34130 6466
rect 36094 6414 36146 6466
rect 37438 6414 37490 6466
rect 40238 6414 40290 6466
rect 40910 6414 40962 6466
rect 46174 6414 46226 6466
rect 46398 6414 46450 6466
rect 46958 6414 47010 6466
rect 47630 6414 47682 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 3502 6078 3554 6130
rect 7086 6078 7138 6130
rect 9774 6078 9826 6130
rect 13470 6078 13522 6130
rect 14478 6078 14530 6130
rect 16382 6078 16434 6130
rect 16718 6078 16770 6130
rect 16830 6078 16882 6130
rect 17502 6078 17554 6130
rect 19294 6078 19346 6130
rect 20974 6078 21026 6130
rect 22094 6078 22146 6130
rect 22990 6078 23042 6130
rect 23886 6078 23938 6130
rect 24334 6078 24386 6130
rect 26126 6078 26178 6130
rect 28366 6078 28418 6130
rect 29934 6078 29986 6130
rect 31726 6078 31778 6130
rect 34750 6078 34802 6130
rect 35198 6078 35250 6130
rect 36206 6078 36258 6130
rect 37214 6078 37266 6130
rect 37662 6078 37714 6130
rect 39342 6078 39394 6130
rect 40238 6078 40290 6130
rect 44718 6078 44770 6130
rect 8430 5966 8482 6018
rect 11006 5966 11058 6018
rect 11454 5966 11506 6018
rect 13694 5966 13746 6018
rect 22542 5966 22594 6018
rect 23326 5966 23378 6018
rect 24558 5966 24610 6018
rect 25566 5966 25618 6018
rect 27134 5966 27186 6018
rect 27694 5966 27746 6018
rect 28590 5966 28642 6018
rect 29262 5966 29314 6018
rect 31950 5966 32002 6018
rect 33518 5966 33570 6018
rect 33742 5966 33794 6018
rect 33966 5966 34018 6018
rect 36430 5966 36482 6018
rect 39566 5966 39618 6018
rect 44382 5966 44434 6018
rect 44494 5966 44546 6018
rect 46062 5966 46114 6018
rect 3838 5854 3890 5906
rect 7422 5854 7474 5906
rect 7646 5854 7698 5906
rect 7982 5854 8034 5906
rect 8094 5854 8146 5906
rect 8654 5854 8706 5906
rect 8766 5854 8818 5906
rect 8990 5854 9042 5906
rect 9998 5854 10050 5906
rect 10222 5854 10274 5906
rect 10670 5854 10722 5906
rect 11230 5854 11282 5906
rect 11342 5854 11394 5906
rect 12910 5854 12962 5906
rect 13134 5854 13186 5906
rect 14142 5854 14194 5906
rect 14254 5854 14306 5906
rect 14702 5854 14754 5906
rect 14926 5854 14978 5906
rect 15486 5854 15538 5906
rect 15598 5854 15650 5906
rect 16046 5854 16098 5906
rect 16606 5854 16658 5906
rect 17614 5854 17666 5906
rect 17726 5854 17778 5906
rect 18062 5854 18114 5906
rect 18622 5854 18674 5906
rect 19070 5854 19122 5906
rect 19966 5854 20018 5906
rect 20190 5854 20242 5906
rect 21534 5854 21586 5906
rect 22318 5854 22370 5906
rect 24110 5854 24162 5906
rect 25118 5854 25170 5906
rect 25342 5854 25394 5906
rect 25790 5854 25842 5906
rect 26350 5854 26402 5906
rect 27358 5854 27410 5906
rect 27918 5854 27970 5906
rect 28478 5854 28530 5906
rect 28814 5854 28866 5906
rect 29374 5854 29426 5906
rect 30382 5854 30434 5906
rect 30606 5854 30658 5906
rect 31054 5854 31106 5906
rect 31502 5854 31554 5906
rect 31614 5854 31666 5906
rect 33070 5854 33122 5906
rect 34414 5854 34466 5906
rect 35758 5854 35810 5906
rect 36654 5854 36706 5906
rect 41022 5854 41074 5906
rect 45278 5854 45330 5906
rect 4622 5742 4674 5794
rect 6750 5742 6802 5794
rect 10110 5742 10162 5794
rect 12350 5742 12402 5794
rect 13582 5742 13634 5794
rect 15822 5742 15874 5794
rect 19182 5742 19234 5794
rect 19630 5742 19682 5794
rect 21198 5742 21250 5794
rect 21758 5742 21810 5794
rect 22206 5742 22258 5794
rect 24222 5742 24274 5794
rect 27246 5742 27298 5794
rect 29038 5742 29090 5794
rect 30830 5742 30882 5794
rect 32510 5742 32562 5794
rect 34078 5742 34130 5794
rect 36766 5742 36818 5794
rect 41806 5742 41858 5794
rect 43934 5742 43986 5794
rect 48190 5742 48242 5794
rect 10558 5630 10610 5682
rect 12574 5630 12626 5682
rect 33182 5630 33234 5682
rect 35870 5630 35922 5682
rect 39678 5630 39730 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 5630 5294 5682 5346
rect 6638 5294 6690 5346
rect 7310 5294 7362 5346
rect 7422 5294 7474 5346
rect 13470 5294 13522 5346
rect 18734 5294 18786 5346
rect 19294 5294 19346 5346
rect 19630 5294 19682 5346
rect 19742 5294 19794 5346
rect 22094 5294 22146 5346
rect 23438 5294 23490 5346
rect 23774 5294 23826 5346
rect 24334 5294 24386 5346
rect 24446 5294 24498 5346
rect 33854 5294 33906 5346
rect 4622 5182 4674 5234
rect 5070 5182 5122 5234
rect 5742 5182 5794 5234
rect 6414 5182 6466 5234
rect 11678 5182 11730 5234
rect 12462 5182 12514 5234
rect 16158 5182 16210 5234
rect 18286 5182 18338 5234
rect 18846 5182 18898 5234
rect 19294 5182 19346 5234
rect 26462 5182 26514 5234
rect 28590 5182 28642 5234
rect 29262 5182 29314 5234
rect 30158 5182 30210 5234
rect 33406 5182 33458 5234
rect 34638 5182 34690 5234
rect 35086 5182 35138 5234
rect 35646 5182 35698 5234
rect 35982 5182 36034 5234
rect 37102 5182 37154 5234
rect 40014 5182 40066 5234
rect 42142 5182 42194 5234
rect 42478 5182 42530 5234
rect 45390 5182 45442 5234
rect 6974 5070 7026 5122
rect 7982 5070 8034 5122
rect 8094 5070 8146 5122
rect 8206 5070 8258 5122
rect 8766 5070 8818 5122
rect 9550 5070 9602 5122
rect 12014 5070 12066 5122
rect 12350 5070 12402 5122
rect 12574 5070 12626 5122
rect 13582 5070 13634 5122
rect 14366 5070 14418 5122
rect 15486 5070 15538 5122
rect 20414 5070 20466 5122
rect 20638 5070 20690 5122
rect 22206 5070 22258 5122
rect 23102 5070 23154 5122
rect 23998 5070 24050 5122
rect 25342 5070 25394 5122
rect 25790 5070 25842 5122
rect 29150 5070 29202 5122
rect 29710 5070 29762 5122
rect 30494 5070 30546 5122
rect 33742 5070 33794 5122
rect 34414 5070 34466 5122
rect 34750 5070 34802 5122
rect 36990 5070 37042 5122
rect 39230 5070 39282 5122
rect 46510 5070 46562 5122
rect 46958 5070 47010 5122
rect 47070 5070 47122 5122
rect 47518 5070 47570 5122
rect 47854 5070 47906 5122
rect 7758 4958 7810 5010
rect 13806 4958 13858 5010
rect 14142 4958 14194 5010
rect 19966 4958 20018 5010
rect 20302 4958 20354 5010
rect 22542 4958 22594 5010
rect 22766 4958 22818 5010
rect 24782 4958 24834 5010
rect 25006 4958 25058 5010
rect 29374 4958 29426 5010
rect 31278 4958 31330 5010
rect 34078 4958 34130 5010
rect 38894 4958 38946 5010
rect 47630 4958 47682 5010
rect 14254 4846 14306 4898
rect 15038 4846 15090 4898
rect 21422 4846 21474 4898
rect 22878 4846 22930 4898
rect 25118 4846 25170 4898
rect 35198 4846 35250 4898
rect 36094 4846 36146 4898
rect 42590 4846 42642 4898
rect 43038 4846 43090 4898
rect 44158 4846 44210 4898
rect 44942 4846 44994 4898
rect 46734 4846 46786 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 5294 4510 5346 4562
rect 5854 4510 5906 4562
rect 9886 4510 9938 4562
rect 10222 4510 10274 4562
rect 24110 4510 24162 4562
rect 24558 4510 24610 4562
rect 25790 4510 25842 4562
rect 26238 4510 26290 4562
rect 26798 4510 26850 4562
rect 30718 4510 30770 4562
rect 31278 4510 31330 4562
rect 31726 4510 31778 4562
rect 31838 4510 31890 4562
rect 40126 4510 40178 4562
rect 41246 4510 41298 4562
rect 44942 4510 44994 4562
rect 16046 4398 16098 4450
rect 25230 4398 25282 4450
rect 28142 4398 28194 4450
rect 31390 4398 31442 4450
rect 35198 4398 35250 4450
rect 38446 4398 38498 4450
rect 39566 4398 39618 4450
rect 41134 4398 41186 4450
rect 43710 4398 43762 4450
rect 46062 4398 46114 4450
rect 6190 4286 6242 4338
rect 13582 4286 13634 4338
rect 16830 4286 16882 4338
rect 17614 4286 17666 4338
rect 20750 4286 20802 4338
rect 27470 4286 27522 4338
rect 31950 4286 32002 4338
rect 32286 4286 32338 4338
rect 35982 4286 36034 4338
rect 39118 4286 39170 4338
rect 44382 4286 44434 4338
rect 45278 4286 45330 4338
rect 6862 4174 6914 4226
rect 8990 4174 9042 4226
rect 10334 4174 10386 4226
rect 10670 4174 10722 4226
rect 12798 4174 12850 4226
rect 13918 4174 13970 4226
rect 18286 4174 18338 4226
rect 20414 4174 20466 4226
rect 21534 4174 21586 4226
rect 23662 4174 23714 4226
rect 30270 4174 30322 4226
rect 33070 4174 33122 4226
rect 36318 4174 36370 4226
rect 41582 4174 41634 4226
rect 48190 4174 48242 4226
rect 25342 4062 25394 4114
rect 39678 4062 39730 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 7534 3726 7586 3778
rect 10334 3726 10386 3778
rect 11230 3726 11282 3778
rect 13134 3726 13186 3778
rect 17614 3726 17666 3778
rect 18846 3726 18898 3778
rect 19518 3726 19570 3778
rect 22094 3726 22146 3778
rect 22430 3726 22482 3778
rect 22878 3726 22930 3778
rect 6414 3614 6466 3666
rect 6862 3614 6914 3666
rect 7310 3614 7362 3666
rect 7646 3614 7698 3666
rect 8430 3614 8482 3666
rect 8878 3614 8930 3666
rect 9998 3614 10050 3666
rect 10446 3614 10498 3666
rect 11342 3614 11394 3666
rect 12238 3614 12290 3666
rect 13246 3614 13298 3666
rect 14142 3614 14194 3666
rect 14590 3614 14642 3666
rect 15038 3614 15090 3666
rect 15822 3614 15874 3666
rect 16494 3614 16546 3666
rect 17726 3614 17778 3666
rect 18398 3614 18450 3666
rect 18846 3614 18898 3666
rect 19294 3614 19346 3666
rect 19630 3614 19682 3666
rect 20078 3614 20130 3666
rect 20974 3614 21026 3666
rect 21422 3614 21474 3666
rect 21870 3614 21922 3666
rect 22206 3614 22258 3666
rect 22766 3614 22818 3666
rect 23214 3614 23266 3666
rect 24110 3614 24162 3666
rect 25342 3614 25394 3666
rect 27470 3614 27522 3666
rect 28590 3614 28642 3666
rect 35534 3614 35586 3666
rect 36766 3614 36818 3666
rect 38894 3614 38946 3666
rect 39790 3614 39842 3666
rect 41918 3614 41970 3666
rect 43822 3614 43874 3666
rect 45054 3614 45106 3666
rect 23662 3502 23714 3554
rect 24558 3502 24610 3554
rect 35982 3502 36034 3554
rect 42590 3502 42642 3554
rect 47630 3502 47682 3554
rect 9550 3390 9602 3442
rect 10894 3390 10946 3442
rect 11790 3390 11842 3442
rect 12686 3390 12738 3442
rect 17390 3390 17442 3442
rect 46958 3390 47010 3442
rect 48190 3390 48242 3442
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 3584 49200 3696 50000
rect 5152 49200 5264 50000
rect 6720 49200 6832 50000
rect 8288 49200 8400 50000
rect 9856 49200 9968 50000
rect 11424 49200 11536 50000
rect 12992 49200 13104 50000
rect 14560 49200 14672 50000
rect 16128 49200 16240 50000
rect 17696 49200 17808 50000
rect 19264 49200 19376 50000
rect 20832 49200 20944 50000
rect 22400 49200 22512 50000
rect 23968 49200 24080 50000
rect 25536 49200 25648 50000
rect 25900 49308 26740 49364
rect 3612 45780 3668 49200
rect 5180 47460 5236 49200
rect 5180 47404 5572 47460
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 3836 45780 3892 45790
rect 3612 45778 3892 45780
rect 3612 45726 3838 45778
rect 3890 45726 3892 45778
rect 3612 45724 3892 45726
rect 3836 45714 3892 45724
rect 5516 45778 5572 47404
rect 5516 45726 5518 45778
rect 5570 45726 5572 45778
rect 5516 45714 5572 45726
rect 6748 45780 6804 49200
rect 8316 47012 8372 49200
rect 8316 46956 8596 47012
rect 6972 45780 7028 45790
rect 6748 45778 7028 45780
rect 6748 45726 6974 45778
rect 7026 45726 7028 45778
rect 6748 45724 7028 45726
rect 6972 45714 7028 45724
rect 8540 45778 8596 46956
rect 9660 45890 9716 45902
rect 9660 45838 9662 45890
rect 9714 45838 9716 45890
rect 9324 45780 9380 45790
rect 8540 45726 8542 45778
rect 8594 45726 8596 45778
rect 8540 45714 8596 45726
rect 9100 45778 9380 45780
rect 9100 45726 9326 45778
rect 9378 45726 9380 45778
rect 9100 45724 9380 45726
rect 5628 45668 5684 45678
rect 2940 45220 2996 45230
rect 2940 45218 3220 45220
rect 2940 45166 2942 45218
rect 2994 45166 3220 45218
rect 2940 45164 3220 45166
rect 2940 45154 2996 45164
rect 3052 44994 3108 45006
rect 3052 44942 3054 44994
rect 3106 44942 3108 44994
rect 3052 44548 3108 44942
rect 2604 44492 3108 44548
rect 2604 44434 2660 44492
rect 2604 44382 2606 44434
rect 2658 44382 2660 44434
rect 2604 44370 2660 44382
rect 1932 44322 1988 44334
rect 1932 44270 1934 44322
rect 1986 44270 1988 44322
rect 1820 43426 1876 43438
rect 1820 43374 1822 43426
rect 1874 43374 1876 43426
rect 1820 42754 1876 43374
rect 1932 43316 1988 44270
rect 3164 44212 3220 45164
rect 5628 45218 5684 45612
rect 7980 45666 8036 45678
rect 7980 45614 7982 45666
rect 8034 45614 8036 45666
rect 7980 45444 8036 45614
rect 7980 45378 8036 45388
rect 8540 45444 8596 45454
rect 5628 45166 5630 45218
rect 5682 45166 5684 45218
rect 5628 45154 5684 45166
rect 8204 45218 8260 45230
rect 8204 45166 8206 45218
rect 8258 45166 8260 45218
rect 3276 45106 3332 45118
rect 3276 45054 3278 45106
rect 3330 45054 3332 45106
rect 3276 44436 3332 45054
rect 3276 44370 3332 44380
rect 3388 45106 3444 45118
rect 3388 45054 3390 45106
rect 3442 45054 3444 45106
rect 3164 44156 3332 44212
rect 3276 43762 3332 44156
rect 3276 43710 3278 43762
rect 3330 43710 3332 43762
rect 3276 43652 3332 43710
rect 3388 43762 3444 45054
rect 4956 45106 5012 45118
rect 4956 45054 4958 45106
rect 5010 45054 5012 45106
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4732 44436 4788 44446
rect 4732 44342 4788 44380
rect 3388 43710 3390 43762
rect 3442 43710 3444 43762
rect 3388 43698 3444 43710
rect 3500 43764 3556 43774
rect 3276 43586 3332 43596
rect 1932 43250 1988 43260
rect 3500 43538 3556 43708
rect 4844 43652 4900 43662
rect 4844 43558 4900 43596
rect 3500 43486 3502 43538
rect 3554 43486 3556 43538
rect 3164 42868 3220 42878
rect 3388 42868 3444 42878
rect 3164 42866 3388 42868
rect 3164 42814 3166 42866
rect 3218 42814 3388 42866
rect 3164 42812 3388 42814
rect 3164 42802 3220 42812
rect 3388 42802 3444 42812
rect 2268 42756 2324 42766
rect 1820 42702 1822 42754
rect 1874 42702 1876 42754
rect 1708 42532 1764 42542
rect 1708 41858 1764 42476
rect 1708 41806 1710 41858
rect 1762 41806 1764 41858
rect 1708 41794 1764 41806
rect 1708 41524 1764 41534
rect 1820 41524 1876 42702
rect 1764 41468 1876 41524
rect 2156 42754 2324 42756
rect 2156 42702 2270 42754
rect 2322 42702 2324 42754
rect 2156 42700 2324 42702
rect 1708 41458 1764 41468
rect 1372 41412 1428 41422
rect 1372 22148 1428 41356
rect 1820 39620 1876 39630
rect 1820 39618 1988 39620
rect 1820 39566 1822 39618
rect 1874 39566 1988 39618
rect 1820 39564 1988 39566
rect 1820 39554 1876 39564
rect 1932 39396 1988 39564
rect 1484 37492 1540 37502
rect 1484 26740 1540 37436
rect 1820 37266 1876 37278
rect 1820 37214 1822 37266
rect 1874 37214 1876 37266
rect 1820 36258 1876 37214
rect 1820 36206 1822 36258
rect 1874 36206 1876 36258
rect 1708 35700 1764 35710
rect 1820 35700 1876 36206
rect 1708 35698 1876 35700
rect 1708 35646 1710 35698
rect 1762 35646 1876 35698
rect 1708 35644 1876 35646
rect 1708 34692 1764 35644
rect 1708 34130 1764 34636
rect 1820 34804 1876 34814
rect 1820 34690 1876 34748
rect 1820 34638 1822 34690
rect 1874 34638 1876 34690
rect 1820 34468 1876 34638
rect 1932 34468 1988 39340
rect 2156 38276 2212 42700
rect 2268 42690 2324 42700
rect 2828 42642 2884 42654
rect 2828 42590 2830 42642
rect 2882 42590 2884 42642
rect 2268 42532 2324 42542
rect 2268 41074 2324 42476
rect 2828 42420 2884 42590
rect 3052 42644 3108 42654
rect 3500 42644 3556 43486
rect 3836 43538 3892 43550
rect 3836 43486 3838 43538
rect 3890 43486 3892 43538
rect 3052 42642 3220 42644
rect 3052 42590 3054 42642
rect 3106 42590 3220 42642
rect 3052 42588 3220 42590
rect 3052 42578 3108 42588
rect 3164 42532 3220 42588
rect 3500 42578 3556 42588
rect 3612 43316 3668 43326
rect 3164 42466 3220 42476
rect 2716 41188 2772 41198
rect 2828 41188 2884 42364
rect 2716 41186 2884 41188
rect 2716 41134 2718 41186
rect 2770 41134 2884 41186
rect 2716 41132 2884 41134
rect 2716 41122 2772 41132
rect 2268 41022 2270 41074
rect 2322 41022 2324 41074
rect 2268 41010 2324 41022
rect 2492 40626 2548 40638
rect 3276 40628 3332 40638
rect 2492 40574 2494 40626
rect 2546 40574 2548 40626
rect 2268 40514 2324 40526
rect 2268 40462 2270 40514
rect 2322 40462 2324 40514
rect 2268 40404 2324 40462
rect 2380 40404 2436 40414
rect 2268 40348 2380 40404
rect 2380 38948 2436 40348
rect 2492 39730 2548 40574
rect 2828 40626 3332 40628
rect 2828 40574 3278 40626
rect 3330 40574 3332 40626
rect 2828 40572 3332 40574
rect 2604 40516 2660 40526
rect 2604 40422 2660 40460
rect 2828 40514 2884 40572
rect 3276 40562 3332 40572
rect 2828 40462 2830 40514
rect 2882 40462 2884 40514
rect 2828 40450 2884 40462
rect 3388 40516 3444 40526
rect 3388 40422 3444 40460
rect 3164 40404 3220 40414
rect 3164 40310 3220 40348
rect 2492 39678 2494 39730
rect 2546 39678 2548 39730
rect 2492 39666 2548 39678
rect 3612 39396 3668 43260
rect 3724 42868 3780 42878
rect 3724 42774 3780 42812
rect 3836 42084 3892 43486
rect 4508 43426 4564 43438
rect 4508 43374 4510 43426
rect 4562 43374 4564 43426
rect 4508 43316 4564 43374
rect 4508 43250 4564 43260
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4844 42980 4900 42990
rect 4732 42866 4788 42878
rect 4732 42814 4734 42866
rect 4786 42814 4788 42866
rect 3612 39330 3668 39340
rect 3724 42028 3892 42084
rect 4060 42754 4116 42766
rect 4060 42702 4062 42754
rect 4114 42702 4116 42754
rect 3724 40402 3780 42028
rect 3836 41858 3892 41870
rect 3836 41806 3838 41858
rect 3890 41806 3892 41858
rect 3836 41300 3892 41806
rect 4060 41300 4116 42702
rect 4732 42644 4788 42814
rect 4844 42754 4900 42924
rect 4844 42702 4846 42754
rect 4898 42702 4900 42754
rect 4844 42690 4900 42702
rect 4732 42578 4788 42588
rect 4620 41972 4676 41982
rect 4956 41972 5012 45054
rect 7756 44996 7812 45006
rect 7420 44994 7812 44996
rect 7420 44942 7758 44994
rect 7810 44942 7812 44994
rect 7420 44940 7812 44942
rect 6188 44436 6244 44446
rect 5740 44380 6020 44436
rect 5740 44324 5796 44380
rect 5404 44268 5796 44324
rect 5404 43538 5460 44268
rect 5740 44210 5796 44268
rect 5740 44158 5742 44210
rect 5794 44158 5796 44210
rect 5740 44146 5796 44158
rect 5852 44210 5908 44222
rect 5852 44158 5854 44210
rect 5906 44158 5908 44210
rect 5404 43486 5406 43538
rect 5458 43486 5460 43538
rect 5404 43474 5460 43486
rect 5516 44098 5572 44110
rect 5516 44046 5518 44098
rect 5570 44046 5572 44098
rect 5516 42756 5572 44046
rect 5852 43876 5908 44158
rect 5964 44212 6020 44380
rect 6188 44342 6244 44380
rect 6300 44212 6356 44222
rect 7420 44212 7476 44940
rect 7756 44930 7812 44940
rect 8092 44884 8148 44894
rect 7868 44882 8148 44884
rect 7868 44830 8094 44882
rect 8146 44830 8148 44882
rect 7868 44828 8148 44830
rect 7756 44324 7812 44334
rect 7756 44230 7812 44268
rect 5964 44210 6580 44212
rect 5964 44158 6302 44210
rect 6354 44158 6580 44210
rect 5964 44156 6580 44158
rect 6300 44146 6356 44156
rect 5740 43820 5908 43876
rect 5740 43428 5796 43820
rect 6524 43762 6580 44156
rect 6524 43710 6526 43762
rect 6578 43710 6580 43762
rect 6524 43698 6580 43710
rect 7196 44210 7476 44212
rect 7196 44158 7422 44210
rect 7474 44158 7476 44210
rect 7196 44156 7476 44158
rect 7196 43650 7252 44156
rect 7420 44146 7476 44156
rect 7756 44100 7812 44110
rect 7308 43764 7364 43774
rect 7308 43670 7364 43708
rect 7756 43762 7812 44044
rect 7756 43710 7758 43762
rect 7810 43710 7812 43762
rect 7756 43698 7812 43710
rect 7196 43598 7198 43650
rect 7250 43598 7252 43650
rect 7196 43586 7252 43598
rect 5740 43334 5796 43372
rect 6076 43538 6132 43550
rect 6076 43486 6078 43538
rect 6130 43486 6132 43538
rect 5628 42756 5684 42766
rect 5516 42754 5684 42756
rect 5516 42702 5630 42754
rect 5682 42702 5684 42754
rect 5516 42700 5684 42702
rect 5628 42690 5684 42700
rect 5964 42756 6020 42766
rect 6076 42756 6132 43486
rect 6748 43538 6804 43550
rect 6748 43486 6750 43538
rect 6802 43486 6804 43538
rect 6636 43426 6692 43438
rect 6636 43374 6638 43426
rect 6690 43374 6692 43426
rect 6300 42980 6356 42990
rect 6300 42886 6356 42924
rect 6636 42980 6692 43374
rect 6636 42914 6692 42924
rect 6748 43428 6804 43486
rect 7868 43538 7924 44828
rect 8092 44818 8148 44828
rect 8204 44212 8260 45166
rect 8428 44882 8484 44894
rect 8428 44830 8430 44882
rect 8482 44830 8484 44882
rect 8428 44324 8484 44830
rect 8428 44258 8484 44268
rect 8092 43764 8148 43774
rect 8204 43764 8260 44156
rect 8148 43708 8260 43764
rect 8092 43698 8148 43708
rect 7868 43486 7870 43538
rect 7922 43486 7924 43538
rect 7868 43474 7924 43486
rect 5964 42754 6132 42756
rect 5964 42702 5966 42754
rect 6018 42702 6132 42754
rect 5964 42700 6132 42702
rect 5964 42690 6020 42700
rect 5740 42644 5796 42654
rect 5740 42550 5796 42588
rect 6412 42642 6468 42654
rect 6412 42590 6414 42642
rect 6466 42590 6468 42642
rect 6300 42532 6356 42542
rect 6300 42438 6356 42476
rect 6412 42420 6468 42590
rect 6748 42644 6804 43372
rect 7868 42868 7924 42878
rect 7868 42866 8036 42868
rect 7868 42814 7870 42866
rect 7922 42814 8036 42866
rect 7868 42812 8036 42814
rect 7868 42802 7924 42812
rect 6972 42756 7028 42766
rect 6972 42754 7476 42756
rect 6972 42702 6974 42754
rect 7026 42702 7476 42754
rect 6972 42700 7476 42702
rect 6972 42690 7028 42700
rect 7420 42644 7476 42700
rect 7532 42644 7588 42654
rect 7756 42644 7812 42654
rect 7420 42642 7588 42644
rect 7420 42590 7534 42642
rect 7586 42590 7588 42642
rect 7420 42588 7588 42590
rect 6748 42578 6804 42588
rect 7084 42532 7140 42542
rect 7196 42532 7252 42542
rect 7084 42530 7196 42532
rect 7084 42478 7086 42530
rect 7138 42478 7196 42530
rect 7084 42476 7196 42478
rect 7084 42466 7140 42476
rect 6412 42354 6468 42364
rect 4620 41970 5012 41972
rect 4620 41918 4622 41970
rect 4674 41918 4958 41970
rect 5010 41918 5012 41970
rect 4620 41916 5012 41918
rect 4620 41906 4676 41916
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 3836 41234 3892 41244
rect 3948 41244 4116 41300
rect 4620 41300 4676 41310
rect 3836 41076 3892 41086
rect 3948 41076 4004 41244
rect 4620 41206 4676 41244
rect 4732 41186 4788 41198
rect 4732 41134 4734 41186
rect 4786 41134 4788 41186
rect 3836 41074 4004 41076
rect 3836 41022 3838 41074
rect 3890 41022 4004 41074
rect 3836 41020 4004 41022
rect 3836 41010 3892 41020
rect 3948 40628 4004 41020
rect 4060 41076 4116 41086
rect 4396 41076 4452 41086
rect 4060 41074 4452 41076
rect 4060 41022 4062 41074
rect 4114 41022 4398 41074
rect 4450 41022 4452 41074
rect 4060 41020 4452 41022
rect 4060 41010 4116 41020
rect 4396 41010 4452 41020
rect 4732 40964 4788 41134
rect 4732 40898 4788 40908
rect 4060 40628 4116 40638
rect 3948 40626 4116 40628
rect 3948 40574 4062 40626
rect 4114 40574 4116 40626
rect 3948 40572 4116 40574
rect 4956 40628 5012 41916
rect 5740 42084 5796 42094
rect 5740 41970 5796 42028
rect 5740 41918 5742 41970
rect 5794 41918 5796 41970
rect 5740 41906 5796 41918
rect 7196 41074 7252 42476
rect 7308 42530 7364 42542
rect 7308 42478 7310 42530
rect 7362 42478 7364 42530
rect 7308 41860 7364 42478
rect 7308 41794 7364 41804
rect 7196 41022 7198 41074
rect 7250 41022 7252 41074
rect 7196 41010 7252 41022
rect 7532 41186 7588 42588
rect 7644 42642 7924 42644
rect 7644 42590 7758 42642
rect 7810 42590 7924 42642
rect 7644 42588 7924 42590
rect 7644 42532 7700 42588
rect 7756 42578 7812 42588
rect 7644 42466 7700 42476
rect 7868 41858 7924 42588
rect 7868 41806 7870 41858
rect 7922 41806 7924 41858
rect 7868 41794 7924 41806
rect 7980 41748 8036 42812
rect 8316 41972 8372 41982
rect 8540 41972 8596 45388
rect 8988 44994 9044 45006
rect 8988 44942 8990 44994
rect 9042 44942 9044 44994
rect 8652 44322 8708 44334
rect 8652 44270 8654 44322
rect 8706 44270 8708 44322
rect 8652 43650 8708 44270
rect 8988 44212 9044 44942
rect 9100 44434 9156 45724
rect 9324 45714 9380 45724
rect 9436 45668 9492 45678
rect 9436 45574 9492 45612
rect 9548 45444 9604 45454
rect 9548 45106 9604 45388
rect 9548 45054 9550 45106
rect 9602 45054 9604 45106
rect 9548 45042 9604 45054
rect 9660 44548 9716 45838
rect 9884 45780 9940 49200
rect 10108 45780 10164 45790
rect 9884 45778 10164 45780
rect 9884 45726 10110 45778
rect 10162 45726 10164 45778
rect 9884 45724 10164 45726
rect 11452 45780 11508 49200
rect 13020 47572 13076 49200
rect 12572 47516 13076 47572
rect 11676 45780 11732 45790
rect 11452 45778 11732 45780
rect 11452 45726 11678 45778
rect 11730 45726 11732 45778
rect 11452 45724 11732 45726
rect 10108 45714 10164 45724
rect 11676 45714 11732 45724
rect 12572 45778 12628 47516
rect 13132 45890 13188 45902
rect 13132 45838 13134 45890
rect 13186 45838 13188 45890
rect 12572 45726 12574 45778
rect 12626 45726 12628 45778
rect 12572 45714 12628 45726
rect 13020 45780 13076 45790
rect 10892 45668 10948 45678
rect 11340 45668 11396 45678
rect 10892 45666 11340 45668
rect 10892 45614 10894 45666
rect 10946 45614 11340 45666
rect 10892 45612 11340 45614
rect 10892 45444 10948 45612
rect 11340 45574 11396 45612
rect 10892 45378 10948 45388
rect 13020 45330 13076 45724
rect 13132 45668 13188 45838
rect 13916 45780 13972 45790
rect 13916 45686 13972 45724
rect 14588 45780 14644 49200
rect 14588 45714 14644 45724
rect 16044 46002 16100 46014
rect 16044 45950 16046 46002
rect 16098 45950 16100 46002
rect 13132 45602 13188 45612
rect 13020 45278 13022 45330
rect 13074 45278 13076 45330
rect 13020 45266 13076 45278
rect 14028 45332 14084 45342
rect 12684 45106 12740 45118
rect 13020 45108 13076 45118
rect 12684 45054 12686 45106
rect 12738 45054 12740 45106
rect 10332 44996 10388 45006
rect 9548 44492 9716 44548
rect 10220 44994 10388 44996
rect 10220 44942 10334 44994
rect 10386 44942 10388 44994
rect 10220 44940 10388 44942
rect 9548 44436 9604 44492
rect 9100 44382 9102 44434
rect 9154 44382 9156 44434
rect 9100 44370 9156 44382
rect 9436 44380 9604 44436
rect 10220 44434 10276 44940
rect 10332 44930 10388 44940
rect 12460 44994 12516 45006
rect 12460 44942 12462 44994
rect 12514 44942 12516 44994
rect 10220 44382 10222 44434
rect 10274 44382 10276 44434
rect 9436 44324 9492 44380
rect 10220 44370 10276 44382
rect 9212 44268 9492 44324
rect 9212 44212 9268 44268
rect 8988 44156 9268 44212
rect 9324 44100 9380 44110
rect 8988 44098 9380 44100
rect 8988 44046 9326 44098
rect 9378 44046 9380 44098
rect 8988 44044 9380 44046
rect 8988 43876 9044 44044
rect 9324 44034 9380 44044
rect 8652 43598 8654 43650
rect 8706 43598 8708 43650
rect 8652 43204 8708 43598
rect 8764 43820 9044 43876
rect 8764 43538 8820 43820
rect 8764 43486 8766 43538
rect 8818 43486 8820 43538
rect 8764 43474 8820 43486
rect 9436 43428 9492 44268
rect 9660 44324 9716 44334
rect 12236 44324 12292 44334
rect 9716 44268 10052 44324
rect 9660 44230 9716 44268
rect 9548 44212 9604 44222
rect 9548 44118 9604 44156
rect 9996 43762 10052 44268
rect 12236 44322 12404 44324
rect 12236 44270 12238 44322
rect 12290 44270 12404 44322
rect 12236 44268 12404 44270
rect 12236 44258 12292 44268
rect 10332 44212 10388 44222
rect 10668 44212 10724 44222
rect 10332 44210 10724 44212
rect 10332 44158 10334 44210
rect 10386 44158 10670 44210
rect 10722 44158 10724 44210
rect 10332 44156 10724 44158
rect 10332 44146 10388 44156
rect 10668 44146 10724 44156
rect 10892 44210 10948 44222
rect 10892 44158 10894 44210
rect 10946 44158 10948 44210
rect 9996 43710 9998 43762
rect 10050 43710 10052 43762
rect 9660 43428 9716 43438
rect 9436 43426 9716 43428
rect 9436 43374 9662 43426
rect 9714 43374 9716 43426
rect 9436 43372 9716 43374
rect 9660 43204 9716 43372
rect 8652 43148 9044 43204
rect 8652 42756 8708 42766
rect 8652 42642 8708 42700
rect 8652 42590 8654 42642
rect 8706 42590 8708 42642
rect 8652 42578 8708 42590
rect 8876 42642 8932 42654
rect 8876 42590 8878 42642
rect 8930 42590 8932 42642
rect 8764 42530 8820 42542
rect 8764 42478 8766 42530
rect 8818 42478 8820 42530
rect 8764 42084 8820 42478
rect 8764 42018 8820 42028
rect 8316 41970 8540 41972
rect 8316 41918 8318 41970
rect 8370 41918 8540 41970
rect 8316 41916 8540 41918
rect 8316 41906 8372 41916
rect 8540 41878 8596 41916
rect 8092 41748 8148 41758
rect 7980 41692 8092 41748
rect 8092 41682 8148 41692
rect 8876 41298 8932 42590
rect 8988 42420 9044 43148
rect 9548 42866 9604 42878
rect 9548 42814 9550 42866
rect 9602 42814 9604 42866
rect 9548 42532 9604 42814
rect 9660 42756 9716 43148
rect 9660 42690 9716 42700
rect 9996 42642 10052 43710
rect 10108 44098 10164 44110
rect 10108 44046 10110 44098
rect 10162 44046 10164 44098
rect 10108 43204 10164 44046
rect 10892 44100 10948 44158
rect 10892 44034 10948 44044
rect 12348 43652 12404 44268
rect 12460 44212 12516 44942
rect 12572 44212 12628 44222
rect 12460 44210 12628 44212
rect 12460 44158 12574 44210
rect 12626 44158 12628 44210
rect 12460 44156 12628 44158
rect 12572 43876 12628 44156
rect 12684 44100 12740 45054
rect 12684 44034 12740 44044
rect 12908 45106 13076 45108
rect 12908 45054 13022 45106
rect 13074 45054 13076 45106
rect 12908 45052 13076 45054
rect 12684 43876 12740 43886
rect 12572 43820 12684 43876
rect 12572 43762 12628 43820
rect 12684 43810 12740 43820
rect 12572 43710 12574 43762
rect 12626 43710 12628 43762
rect 12572 43698 12628 43710
rect 12796 43764 12852 43774
rect 12908 43764 12964 45052
rect 13020 45042 13076 45052
rect 13244 45106 13300 45118
rect 13244 45054 13246 45106
rect 13298 45054 13300 45106
rect 12796 43762 12964 43764
rect 12796 43710 12798 43762
rect 12850 43710 12964 43762
rect 12796 43708 12964 43710
rect 13020 43764 13076 43774
rect 12796 43698 12852 43708
rect 13020 43670 13076 43708
rect 13132 43764 13188 43774
rect 13244 43764 13300 45054
rect 14028 45106 14084 45276
rect 14588 45108 14644 45118
rect 14028 45054 14030 45106
rect 14082 45054 14084 45106
rect 14028 45042 14084 45054
rect 14476 45052 14588 45108
rect 13132 43762 13300 43764
rect 13132 43710 13134 43762
rect 13186 43710 13300 43762
rect 13132 43708 13300 43710
rect 13356 43876 13412 43886
rect 13132 43698 13188 43708
rect 12460 43652 12516 43662
rect 12348 43596 12460 43652
rect 10108 43138 10164 43148
rect 10332 43538 10388 43550
rect 10332 43486 10334 43538
rect 10386 43486 10388 43538
rect 10332 42980 10388 43486
rect 10780 43426 10836 43438
rect 10780 43374 10782 43426
rect 10834 43374 10836 43426
rect 10780 43204 10836 43374
rect 10780 43138 10836 43148
rect 11340 43426 11396 43438
rect 11340 43374 11342 43426
rect 11394 43374 11396 43426
rect 11340 43314 11396 43374
rect 11340 43262 11342 43314
rect 11394 43262 11396 43314
rect 10332 42924 10836 42980
rect 9996 42590 9998 42642
rect 10050 42590 10052 42642
rect 9996 42578 10052 42590
rect 10332 42644 10388 42654
rect 9548 42476 9940 42532
rect 8988 42364 9828 42420
rect 9548 42196 9604 42206
rect 9436 41970 9492 41982
rect 9436 41918 9438 41970
rect 9490 41918 9492 41970
rect 9436 41860 9492 41918
rect 9436 41794 9492 41804
rect 8876 41246 8878 41298
rect 8930 41246 8932 41298
rect 8876 41234 8932 41246
rect 8316 41188 8372 41198
rect 7532 41134 7534 41186
rect 7586 41134 7588 41186
rect 5852 40964 5908 40974
rect 5852 40870 5908 40908
rect 7084 40964 7140 40974
rect 5068 40628 5124 40638
rect 4956 40626 5236 40628
rect 4956 40574 5070 40626
rect 5122 40574 5236 40626
rect 4956 40572 5236 40574
rect 4060 40562 4116 40572
rect 5068 40562 5124 40572
rect 3724 40350 3726 40402
rect 3778 40350 3780 40402
rect 3724 39172 3780 40350
rect 3500 39116 3780 39172
rect 3836 40516 3892 40526
rect 2492 38948 2548 38958
rect 2380 38946 2548 38948
rect 2380 38894 2494 38946
rect 2546 38894 2548 38946
rect 2380 38892 2548 38894
rect 2492 38882 2548 38892
rect 3164 38836 3220 38846
rect 3164 38742 3220 38780
rect 3388 38724 3444 38762
rect 3388 38658 3444 38668
rect 2156 38210 2212 38220
rect 3164 38164 3220 38174
rect 3164 38070 3220 38108
rect 3388 38164 3444 38174
rect 2268 37828 2324 37838
rect 2156 37826 2324 37828
rect 2156 37774 2270 37826
rect 2322 37774 2324 37826
rect 2156 37772 2324 37774
rect 2156 37044 2212 37772
rect 2268 37762 2324 37772
rect 2492 37156 2548 37166
rect 2492 37062 2548 37100
rect 2156 35308 2212 36988
rect 1820 34412 1932 34468
rect 1932 34402 1988 34412
rect 2044 35252 2212 35308
rect 2268 36258 2324 36270
rect 2268 36206 2270 36258
rect 2322 36206 2324 36258
rect 2044 34244 2100 35252
rect 1708 34078 1710 34130
rect 1762 34078 1764 34130
rect 1708 34066 1764 34078
rect 1820 34188 2100 34244
rect 2268 35140 2324 36206
rect 2492 36260 2548 36270
rect 2492 35810 2548 36204
rect 2492 35758 2494 35810
rect 2546 35758 2548 35810
rect 2492 35746 2548 35758
rect 2716 36258 2772 36270
rect 3164 36260 3220 36270
rect 2716 36206 2718 36258
rect 2770 36206 2772 36258
rect 1708 33236 1764 33246
rect 1708 33142 1764 33180
rect 1820 33234 1876 34188
rect 1820 33182 1822 33234
rect 1874 33182 1876 33234
rect 1820 33170 1876 33182
rect 1932 34020 1988 34030
rect 1932 32900 1988 33964
rect 2268 33234 2324 35084
rect 2716 35140 2772 36206
rect 2716 35074 2772 35084
rect 3052 36258 3220 36260
rect 3052 36206 3166 36258
rect 3218 36206 3220 36258
rect 3052 36204 3220 36206
rect 2604 34916 2660 34926
rect 2604 34914 2884 34916
rect 2604 34862 2606 34914
rect 2658 34862 2884 34914
rect 2604 34860 2884 34862
rect 2604 34850 2660 34860
rect 2380 34690 2436 34702
rect 2380 34638 2382 34690
rect 2434 34638 2436 34690
rect 2380 33684 2436 34638
rect 2716 34690 2772 34702
rect 2716 34638 2718 34690
rect 2770 34638 2772 34690
rect 2716 34356 2772 34638
rect 2492 34300 2772 34356
rect 2492 34242 2548 34300
rect 2492 34190 2494 34242
rect 2546 34190 2548 34242
rect 2492 34178 2548 34190
rect 2828 34244 2884 34860
rect 2380 33618 2436 33628
rect 2268 33182 2270 33234
rect 2322 33182 2324 33234
rect 2044 33124 2100 33134
rect 2044 33030 2100 33068
rect 2268 33012 2324 33182
rect 2268 32946 2324 32956
rect 2380 33122 2436 33134
rect 2380 33070 2382 33122
rect 2434 33070 2436 33122
rect 1708 32844 1988 32900
rect 1708 31892 1764 32844
rect 2380 32788 2436 33070
rect 1708 30994 1764 31836
rect 1708 30942 1710 30994
rect 1762 30942 1764 30994
rect 1708 28532 1764 30942
rect 1820 32732 2436 32788
rect 2604 33122 2660 33134
rect 2604 33070 2606 33122
rect 2658 33070 2660 33122
rect 1820 30100 1876 32732
rect 2044 32562 2100 32574
rect 2044 32510 2046 32562
rect 2098 32510 2100 32562
rect 2044 32228 2100 32510
rect 2044 32162 2100 32172
rect 2268 32562 2324 32574
rect 2268 32510 2270 32562
rect 2322 32510 2324 32562
rect 2268 32116 2324 32510
rect 2492 32562 2548 32574
rect 2492 32510 2494 32562
rect 2546 32510 2548 32562
rect 2268 32050 2324 32060
rect 2380 32450 2436 32462
rect 2380 32398 2382 32450
rect 2434 32398 2436 32450
rect 1932 31780 1988 31790
rect 2380 31780 2436 32398
rect 2492 32004 2548 32510
rect 2492 31938 2548 31948
rect 1932 31778 2324 31780
rect 1932 31726 1934 31778
rect 1986 31726 2324 31778
rect 1932 31724 2324 31726
rect 2380 31724 2548 31780
rect 1932 31714 1988 31724
rect 2044 31554 2100 31566
rect 2044 31502 2046 31554
rect 2098 31502 2100 31554
rect 1932 30324 1988 30334
rect 2044 30324 2100 31502
rect 2156 31554 2212 31566
rect 2156 31502 2158 31554
rect 2210 31502 2212 31554
rect 2156 31220 2212 31502
rect 2156 30436 2212 31164
rect 2268 30772 2324 31724
rect 2380 31556 2436 31566
rect 2380 31462 2436 31500
rect 2492 31106 2548 31724
rect 2492 31054 2494 31106
rect 2546 31054 2548 31106
rect 2492 31042 2548 31054
rect 2268 30716 2548 30772
rect 2156 30380 2324 30436
rect 2044 30268 2212 30324
rect 1932 30230 1988 30268
rect 2044 30100 2100 30110
rect 1820 30098 1988 30100
rect 1820 30046 1822 30098
rect 1874 30046 1988 30098
rect 1820 30044 1988 30046
rect 1820 30034 1876 30044
rect 1820 29876 1876 29886
rect 1820 28754 1876 29820
rect 1820 28702 1822 28754
rect 1874 28702 1876 28754
rect 1820 28690 1876 28702
rect 1932 29092 1988 30044
rect 2044 30006 2100 30044
rect 2156 29876 2212 30268
rect 2044 29820 2212 29876
rect 2044 29426 2100 29820
rect 2044 29374 2046 29426
rect 2098 29374 2100 29426
rect 2044 29362 2100 29374
rect 2156 29428 2212 29438
rect 2268 29428 2324 30380
rect 2156 29426 2324 29428
rect 2156 29374 2158 29426
rect 2210 29374 2324 29426
rect 2156 29372 2324 29374
rect 2492 29538 2548 30716
rect 2492 29486 2494 29538
rect 2546 29486 2548 29538
rect 2156 29204 2212 29372
rect 2380 29316 2436 29326
rect 1820 28532 1876 28542
rect 1708 28476 1820 28532
rect 1820 28466 1876 28476
rect 1484 26674 1540 26684
rect 1596 28308 1652 28318
rect 1932 28308 1988 29036
rect 1596 25284 1652 28252
rect 1708 28252 1988 28308
rect 2044 29148 2212 29204
rect 2268 29314 2436 29316
rect 2268 29262 2382 29314
rect 2434 29262 2436 29314
rect 2268 29260 2436 29262
rect 1708 27746 1764 28252
rect 2044 28196 2100 29148
rect 1932 28140 2100 28196
rect 2156 28756 2212 28766
rect 1708 27694 1710 27746
rect 1762 27694 1764 27746
rect 1708 27682 1764 27694
rect 1820 28084 1876 28094
rect 1484 25228 1652 25284
rect 1708 26292 1764 26302
rect 1484 25172 1540 25228
rect 1484 25106 1540 25116
rect 1372 22082 1428 22092
rect 1596 24948 1652 24958
rect 1484 22036 1540 22046
rect 1148 21364 1204 21374
rect 1036 19908 1092 19918
rect 1036 15204 1092 19852
rect 1148 15428 1204 21308
rect 1260 18900 1316 18910
rect 1260 16996 1316 18844
rect 1484 17220 1540 21980
rect 1484 17154 1540 17164
rect 1596 17108 1652 24892
rect 1708 22484 1764 26236
rect 1820 25506 1876 28028
rect 1932 26908 1988 28140
rect 2044 27188 2100 27198
rect 2156 27188 2212 28700
rect 2044 27186 2212 27188
rect 2044 27134 2046 27186
rect 2098 27134 2212 27186
rect 2044 27132 2212 27134
rect 2044 27122 2100 27132
rect 2268 26908 2324 29260
rect 2380 29250 2436 29260
rect 2380 29092 2436 29102
rect 2380 28530 2436 29036
rect 2492 28868 2548 29486
rect 2604 29428 2660 33070
rect 2828 33124 2884 34188
rect 2940 34802 2996 34814
rect 2940 34750 2942 34802
rect 2994 34750 2996 34802
rect 2940 33572 2996 34750
rect 3052 34804 3108 36204
rect 3164 36194 3220 36204
rect 3052 34738 3108 34748
rect 3164 34802 3220 34814
rect 3164 34750 3166 34802
rect 3218 34750 3220 34802
rect 2940 33506 2996 33516
rect 3052 33460 3108 33470
rect 3164 33460 3220 34750
rect 3388 34692 3444 38108
rect 3388 34626 3444 34636
rect 3500 37492 3556 39116
rect 3836 38834 3892 40460
rect 4620 40292 4676 40302
rect 4620 40290 4900 40292
rect 4620 40238 4622 40290
rect 4674 40238 4900 40290
rect 4620 40236 4900 40238
rect 4620 40226 4676 40236
rect 4396 40180 4452 40190
rect 4284 40178 4452 40180
rect 4284 40126 4398 40178
rect 4450 40126 4452 40178
rect 4284 40124 4452 40126
rect 4284 39058 4340 40124
rect 4396 40114 4452 40124
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4620 39732 4676 39742
rect 4284 39006 4286 39058
rect 4338 39006 4340 39058
rect 4284 38994 4340 39006
rect 4508 39730 4676 39732
rect 4508 39678 4622 39730
rect 4674 39678 4676 39730
rect 4508 39676 4676 39678
rect 3836 38782 3838 38834
rect 3890 38782 3892 38834
rect 3836 38724 3892 38782
rect 4172 38836 4228 38846
rect 4172 38742 4228 38780
rect 4396 38834 4452 38846
rect 4396 38782 4398 38834
rect 4450 38782 4452 38834
rect 3612 38668 3892 38724
rect 4396 38724 4452 38782
rect 4508 38836 4564 39676
rect 4620 39666 4676 39676
rect 4844 39508 4900 40236
rect 4620 39452 4900 39508
rect 4620 39058 4676 39452
rect 5068 39396 5124 39406
rect 5068 39302 5124 39340
rect 4620 39006 4622 39058
rect 4674 39006 4676 39058
rect 4620 38994 4676 39006
rect 4508 38770 4564 38780
rect 4844 38946 4900 38958
rect 4844 38894 4846 38946
rect 4898 38894 4900 38946
rect 4844 38836 4900 38894
rect 4844 38770 4900 38780
rect 4956 38834 5012 38846
rect 4956 38782 4958 38834
rect 5010 38782 5012 38834
rect 3612 38274 3668 38668
rect 4396 38658 4452 38668
rect 4956 38724 5012 38782
rect 4956 38658 5012 38668
rect 5180 38612 5236 40572
rect 6972 40514 7028 40526
rect 6972 40462 6974 40514
rect 7026 40462 7028 40514
rect 6860 40402 6916 40414
rect 6860 40350 6862 40402
rect 6914 40350 6916 40402
rect 5628 39618 5684 39630
rect 5628 39566 5630 39618
rect 5682 39566 5684 39618
rect 5628 39396 5684 39566
rect 6412 39508 6468 39518
rect 5628 39330 5684 39340
rect 5964 39506 6468 39508
rect 5964 39454 6414 39506
rect 6466 39454 6468 39506
rect 5964 39452 6468 39454
rect 5964 39058 6020 39452
rect 6412 39442 6468 39452
rect 5964 39006 5966 39058
rect 6018 39006 6020 39058
rect 5964 38994 6020 39006
rect 6860 38948 6916 40350
rect 5068 38556 5180 38612
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 3612 38222 3614 38274
rect 3666 38222 3668 38274
rect 3612 38210 3668 38222
rect 5068 38164 5124 38556
rect 5180 38546 5236 38556
rect 5628 38834 5684 38846
rect 5628 38782 5630 38834
rect 5682 38782 5684 38834
rect 5628 38274 5684 38782
rect 5852 38834 5908 38846
rect 5852 38782 5854 38834
rect 5906 38782 5908 38834
rect 5852 38500 5908 38782
rect 6188 38836 6244 38846
rect 6188 38834 6468 38836
rect 6188 38782 6190 38834
rect 6242 38782 6468 38834
rect 6188 38780 6468 38782
rect 6188 38770 6244 38780
rect 5852 38434 5908 38444
rect 6412 38722 6468 38780
rect 6412 38670 6414 38722
rect 6466 38670 6468 38722
rect 5628 38222 5630 38274
rect 5682 38222 5684 38274
rect 5628 38210 5684 38222
rect 6188 38276 6244 38286
rect 6188 38274 6356 38276
rect 6188 38222 6190 38274
rect 6242 38222 6356 38274
rect 6188 38220 6356 38222
rect 6188 38210 6244 38220
rect 5068 38070 5124 38108
rect 3724 38052 3780 38062
rect 4172 38052 4228 38062
rect 3724 38050 4228 38052
rect 3724 37998 3726 38050
rect 3778 37998 4174 38050
rect 4226 37998 4228 38050
rect 3724 37996 4228 37998
rect 3724 37986 3780 37996
rect 4172 37986 4228 37996
rect 4732 38050 4788 38062
rect 4732 37998 4734 38050
rect 4786 37998 4788 38050
rect 3052 33458 3220 33460
rect 3052 33406 3054 33458
rect 3106 33406 3220 33458
rect 3052 33404 3220 33406
rect 3276 33572 3332 33582
rect 3052 33394 3108 33404
rect 3164 33236 3220 33246
rect 3276 33236 3332 33516
rect 3500 33236 3556 37436
rect 3612 37826 3668 37838
rect 4060 37828 4116 37838
rect 4284 37828 4340 37838
rect 4732 37828 4788 37998
rect 3612 37774 3614 37826
rect 3666 37774 3668 37826
rect 3612 36260 3668 37774
rect 3948 37826 4116 37828
rect 3948 37774 4062 37826
rect 4114 37774 4116 37826
rect 3948 37772 4116 37774
rect 3948 36484 4004 37772
rect 4060 37762 4116 37772
rect 4172 37826 4452 37828
rect 4172 37774 4286 37826
rect 4338 37774 4452 37826
rect 4172 37772 4452 37774
rect 3948 36418 4004 36428
rect 4060 36484 4116 36494
rect 4172 36484 4228 37772
rect 4284 37762 4340 37772
rect 4284 37268 4340 37278
rect 4284 36708 4340 37212
rect 4396 37156 4452 37772
rect 4732 37762 4788 37772
rect 5292 37828 5348 37838
rect 4732 37492 4788 37502
rect 5180 37492 5236 37502
rect 4788 37436 4900 37492
rect 4732 37426 4788 37436
rect 4844 37266 4900 37436
rect 4844 37214 4846 37266
rect 4898 37214 4900 37266
rect 4844 37202 4900 37214
rect 4620 37156 4676 37166
rect 4396 37154 4788 37156
rect 4396 37102 4622 37154
rect 4674 37102 4788 37154
rect 4396 37100 4788 37102
rect 4620 37090 4676 37100
rect 4732 37044 4788 37100
rect 4732 36988 5012 37044
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4284 36652 4564 36708
rect 4508 36594 4564 36652
rect 4508 36542 4510 36594
rect 4562 36542 4564 36594
rect 4508 36530 4564 36542
rect 4060 36482 4228 36484
rect 4060 36430 4062 36482
rect 4114 36430 4228 36482
rect 4060 36428 4228 36430
rect 4396 36484 4452 36494
rect 4060 36418 4116 36428
rect 4396 36390 4452 36428
rect 4844 36372 4900 36382
rect 4732 36260 4788 36270
rect 3612 36258 4788 36260
rect 3612 36206 4734 36258
rect 4786 36206 4788 36258
rect 3612 36204 4788 36206
rect 4732 36194 4788 36204
rect 4620 35588 4676 35598
rect 4844 35588 4900 36316
rect 4956 36370 5012 36988
rect 5180 36932 5236 37436
rect 5292 37266 5348 37772
rect 5516 37828 5572 37838
rect 5740 37828 5796 37838
rect 5572 37826 5796 37828
rect 5572 37774 5742 37826
rect 5794 37774 5796 37826
rect 5572 37772 5796 37774
rect 6300 37828 6356 38220
rect 6412 38050 6468 38670
rect 6860 38722 6916 38892
rect 6972 39060 7028 40462
rect 6972 38834 7028 39004
rect 6972 38782 6974 38834
rect 7026 38782 7028 38834
rect 6972 38770 7028 38782
rect 6860 38670 6862 38722
rect 6914 38670 6916 38722
rect 6860 38658 6916 38670
rect 7084 38668 7140 40908
rect 7196 40404 7252 40414
rect 7420 40404 7476 40414
rect 7196 40402 7476 40404
rect 7196 40350 7198 40402
rect 7250 40350 7422 40402
rect 7474 40350 7476 40402
rect 7196 40348 7476 40350
rect 7196 40338 7252 40348
rect 7420 40338 7476 40348
rect 7532 40180 7588 41134
rect 7980 41132 8316 41188
rect 7756 40964 7812 40974
rect 7532 40114 7588 40124
rect 7644 40178 7700 40190
rect 7644 40126 7646 40178
rect 7698 40126 7700 40178
rect 7644 39172 7700 40126
rect 7532 39116 7700 39172
rect 7532 38836 7588 39116
rect 7532 38770 7588 38780
rect 7644 38834 7700 38846
rect 7644 38782 7646 38834
rect 7698 38782 7700 38834
rect 7084 38612 7588 38668
rect 6412 37998 6414 38050
rect 6466 37998 6468 38050
rect 6412 37986 6468 37998
rect 6636 38500 6692 38510
rect 6636 38050 6692 38444
rect 6636 37998 6638 38050
rect 6690 37998 6692 38050
rect 6524 37828 6580 37838
rect 6300 37826 6580 37828
rect 6300 37774 6526 37826
rect 6578 37774 6580 37826
rect 6300 37772 6580 37774
rect 5516 37762 5572 37772
rect 5740 37762 5796 37772
rect 6524 37762 6580 37772
rect 5404 37492 5460 37502
rect 5404 37490 6356 37492
rect 5404 37438 5406 37490
rect 5458 37438 6356 37490
rect 5404 37436 6356 37438
rect 5404 37426 5460 37436
rect 5292 37214 5294 37266
rect 5346 37214 5348 37266
rect 5292 37044 5348 37214
rect 5516 37268 5572 37278
rect 5740 37268 5796 37278
rect 5572 37266 5796 37268
rect 5572 37214 5742 37266
rect 5794 37214 5796 37266
rect 5572 37212 5796 37214
rect 5516 37174 5572 37212
rect 5740 37202 5796 37212
rect 5852 37268 5908 37278
rect 5292 36978 5348 36988
rect 5180 36866 5236 36876
rect 5404 36932 5460 36942
rect 5460 36876 5796 36932
rect 5404 36866 5460 36876
rect 5292 36820 5348 36830
rect 4956 36318 4958 36370
rect 5010 36318 5012 36370
rect 4956 36306 5012 36318
rect 5068 36484 5124 36494
rect 5068 36370 5124 36428
rect 5068 36318 5070 36370
rect 5122 36318 5124 36370
rect 5068 36148 5124 36318
rect 5068 36082 5124 36092
rect 4620 35586 4900 35588
rect 4620 35534 4622 35586
rect 4674 35534 4900 35586
rect 4620 35532 4900 35534
rect 5292 35586 5348 36764
rect 5740 35924 5796 36876
rect 5852 36706 5908 37212
rect 6188 37266 6244 37278
rect 6188 37214 6190 37266
rect 6242 37214 6244 37266
rect 5964 37156 6020 37166
rect 5964 37062 6020 37100
rect 6188 37044 6244 37214
rect 6300 37266 6356 37436
rect 6636 37490 6692 37998
rect 7084 38052 7140 38062
rect 7084 37958 7140 37996
rect 6636 37438 6638 37490
rect 6690 37438 6692 37490
rect 6636 37426 6692 37438
rect 7532 37828 7588 38612
rect 7644 38500 7700 38782
rect 7644 38434 7700 38444
rect 7644 37828 7700 37838
rect 7532 37826 7700 37828
rect 7532 37774 7646 37826
rect 7698 37774 7700 37826
rect 7532 37772 7700 37774
rect 6300 37214 6302 37266
rect 6354 37214 6356 37266
rect 6300 37202 6356 37214
rect 6860 37378 6916 37390
rect 6860 37326 6862 37378
rect 6914 37326 6916 37378
rect 6860 37268 6916 37326
rect 6860 37202 6916 37212
rect 6972 37268 7028 37278
rect 6972 37266 7364 37268
rect 6972 37214 6974 37266
rect 7026 37214 7364 37266
rect 6972 37212 7364 37214
rect 6972 37202 7028 37212
rect 6188 36978 6244 36988
rect 5852 36654 5854 36706
rect 5906 36654 5908 36706
rect 5852 36642 5908 36654
rect 7308 36594 7364 37212
rect 7308 36542 7310 36594
rect 7362 36542 7364 36594
rect 7308 36530 7364 36542
rect 6188 36484 6244 36494
rect 5852 36372 5908 36382
rect 5852 36278 5908 36316
rect 5964 36372 6020 36382
rect 6188 36372 6244 36428
rect 6524 36482 6580 36494
rect 6524 36430 6526 36482
rect 6578 36430 6580 36482
rect 5964 36370 6244 36372
rect 5964 36318 5966 36370
rect 6018 36318 6244 36370
rect 5964 36316 6244 36318
rect 5964 36306 6020 36316
rect 5740 35922 6132 35924
rect 5740 35870 5742 35922
rect 5794 35870 6132 35922
rect 5740 35868 6132 35870
rect 5740 35858 5796 35868
rect 5292 35534 5294 35586
rect 5346 35534 5348 35586
rect 4620 35522 4676 35532
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 3724 35140 3780 35150
rect 3724 35026 3780 35084
rect 3724 34974 3726 35026
rect 3778 34974 3780 35026
rect 3724 34962 3780 34974
rect 5292 35028 5348 35534
rect 5740 35364 5796 35374
rect 5292 34972 5572 35028
rect 5180 34916 5236 34926
rect 5236 34860 5348 34916
rect 5180 34850 5236 34860
rect 4172 34804 4228 34814
rect 4172 34710 4228 34748
rect 4620 34692 4676 34702
rect 4620 34598 4676 34636
rect 5180 34692 5236 34702
rect 5180 34598 5236 34636
rect 5068 34244 5124 34254
rect 4844 34132 4900 34142
rect 4620 34020 4676 34030
rect 4284 34018 4676 34020
rect 4284 33966 4622 34018
rect 4674 33966 4676 34018
rect 4284 33964 4676 33966
rect 4284 33460 4340 33964
rect 4620 33954 4676 33964
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4508 33572 4564 33582
rect 4844 33572 4900 34076
rect 4956 34132 5012 34142
rect 5068 34132 5124 34188
rect 4956 34130 5124 34132
rect 4956 34078 4958 34130
rect 5010 34078 5124 34130
rect 4956 34076 5124 34078
rect 5180 34132 5236 34142
rect 5292 34132 5348 34860
rect 5180 34130 5348 34132
rect 5180 34078 5182 34130
rect 5234 34078 5348 34130
rect 5180 34076 5348 34078
rect 4956 34066 5012 34076
rect 5180 34066 5236 34076
rect 5516 33796 5572 34972
rect 5740 35026 5796 35308
rect 5740 34974 5742 35026
rect 5794 34974 5796 35026
rect 5740 34962 5796 34974
rect 5628 34916 5684 34926
rect 5628 34822 5684 34860
rect 5852 34692 5908 34702
rect 5628 34690 5908 34692
rect 5628 34638 5854 34690
rect 5906 34638 5908 34690
rect 5628 34636 5908 34638
rect 5628 34132 5684 34636
rect 5852 34626 5908 34636
rect 6076 34468 6132 35868
rect 6188 35698 6244 36316
rect 6300 36370 6356 36382
rect 6300 36318 6302 36370
rect 6354 36318 6356 36370
rect 6300 35812 6356 36318
rect 6412 36260 6468 36270
rect 6412 36166 6468 36204
rect 6300 35746 6356 35756
rect 6524 35924 6580 36430
rect 7196 36484 7252 36494
rect 7196 36390 7252 36428
rect 6188 35646 6190 35698
rect 6242 35646 6244 35698
rect 6188 35634 6244 35646
rect 6524 35364 6580 35868
rect 6636 36372 6692 36382
rect 6636 35698 6692 36316
rect 6860 36372 6916 36382
rect 7420 36372 7476 36382
rect 6860 36370 7140 36372
rect 6860 36318 6862 36370
rect 6914 36318 7140 36370
rect 6860 36316 7140 36318
rect 6860 36306 6916 36316
rect 7084 36036 7140 36316
rect 7420 36278 7476 36316
rect 7532 36260 7588 37772
rect 7644 37762 7700 37772
rect 7644 37492 7700 37502
rect 7644 37398 7700 37436
rect 7532 36194 7588 36204
rect 7644 36258 7700 36270
rect 7644 36206 7646 36258
rect 7698 36206 7700 36258
rect 7084 35980 7588 36036
rect 7532 35922 7588 35980
rect 7532 35870 7534 35922
rect 7586 35870 7588 35922
rect 7532 35858 7588 35870
rect 7644 35924 7700 36206
rect 7644 35830 7700 35868
rect 7084 35812 7140 35822
rect 7420 35812 7476 35822
rect 7140 35810 7476 35812
rect 7140 35758 7422 35810
rect 7474 35758 7476 35810
rect 7140 35756 7476 35758
rect 7084 35718 7140 35756
rect 7420 35746 7476 35756
rect 7756 35700 7812 40908
rect 7980 40626 8036 41132
rect 8316 41094 8372 41132
rect 9324 40962 9380 40974
rect 9324 40910 9326 40962
rect 9378 40910 9380 40962
rect 7980 40574 7982 40626
rect 8034 40574 8036 40626
rect 7980 40562 8036 40574
rect 8316 40852 8372 40862
rect 8316 39284 8372 40796
rect 8652 40404 8708 40414
rect 9100 40404 9156 40414
rect 8652 40402 9156 40404
rect 8652 40350 8654 40402
rect 8706 40350 9102 40402
rect 9154 40350 9156 40402
rect 8652 40348 9156 40350
rect 8652 40338 8708 40348
rect 8540 39730 8596 39742
rect 8540 39678 8542 39730
rect 8594 39678 8596 39730
rect 7980 39228 8372 39284
rect 8428 39396 8484 39406
rect 7980 38668 8036 39228
rect 8092 39060 8148 39070
rect 8092 38966 8148 39004
rect 8316 38948 8372 38958
rect 8316 38854 8372 38892
rect 8204 38836 8260 38846
rect 8204 38742 8260 38780
rect 8428 38668 8484 39340
rect 8540 39060 8596 39678
rect 8988 39508 9044 39518
rect 8876 39452 8988 39508
rect 8876 39394 8932 39452
rect 8988 39442 9044 39452
rect 8876 39342 8878 39394
rect 8930 39342 8932 39394
rect 8876 39330 8932 39342
rect 8540 38994 8596 39004
rect 6636 35646 6638 35698
rect 6690 35646 6692 35698
rect 6636 35634 6692 35646
rect 7532 35644 7812 35700
rect 7868 38612 8036 38668
rect 8316 38612 8484 38668
rect 8652 38948 8708 38958
rect 6524 35298 6580 35308
rect 6972 35084 7364 35140
rect 6188 34916 6244 34926
rect 6412 34916 6468 34926
rect 6188 34914 6468 34916
rect 6188 34862 6190 34914
rect 6242 34862 6414 34914
rect 6466 34862 6468 34914
rect 6188 34860 6468 34862
rect 6188 34850 6244 34860
rect 6412 34850 6468 34860
rect 6748 34916 6804 34926
rect 6748 34914 6916 34916
rect 6748 34862 6750 34914
rect 6802 34862 6916 34914
rect 6748 34860 6916 34862
rect 6748 34850 6804 34860
rect 6636 34692 6692 34702
rect 6076 34402 6132 34412
rect 6412 34690 6692 34692
rect 6412 34638 6638 34690
rect 6690 34638 6692 34690
rect 6412 34636 6692 34638
rect 6300 34132 6356 34142
rect 5628 34038 5684 34076
rect 5740 34130 6356 34132
rect 5740 34078 6302 34130
rect 6354 34078 6356 34130
rect 5740 34076 6356 34078
rect 4508 33570 4900 33572
rect 4508 33518 4510 33570
rect 4562 33518 4900 33570
rect 4508 33516 4900 33518
rect 5292 33740 5572 33796
rect 4508 33506 4564 33516
rect 4396 33460 4452 33470
rect 4284 33458 4452 33460
rect 4284 33406 4398 33458
rect 4450 33406 4452 33458
rect 4284 33404 4452 33406
rect 4396 33394 4452 33404
rect 3612 33348 3668 33358
rect 3612 33346 3892 33348
rect 3612 33294 3614 33346
rect 3666 33294 3892 33346
rect 3612 33292 3892 33294
rect 3612 33282 3668 33292
rect 3164 33234 3332 33236
rect 3164 33182 3166 33234
rect 3218 33182 3332 33234
rect 3164 33180 3332 33182
rect 3388 33180 3556 33236
rect 2940 33124 2996 33134
rect 2828 33122 2996 33124
rect 2828 33070 2942 33122
rect 2994 33070 2996 33122
rect 2828 33068 2996 33070
rect 2940 33058 2996 33068
rect 3164 32900 3220 33180
rect 3164 32834 3220 32844
rect 3388 32788 3444 33180
rect 3724 33124 3780 33134
rect 3276 32732 3444 32788
rect 3500 33122 3780 33124
rect 3500 33070 3726 33122
rect 3778 33070 3780 33122
rect 3500 33068 3780 33070
rect 3052 32676 3108 32686
rect 3052 32582 3108 32620
rect 2828 32564 2884 32574
rect 2716 32508 2828 32564
rect 2716 31556 2772 32508
rect 2828 32470 2884 32508
rect 2940 32450 2996 32462
rect 2940 32398 2942 32450
rect 2994 32398 2996 32450
rect 2940 32004 2996 32398
rect 3052 32004 3108 32014
rect 2940 32002 3108 32004
rect 2940 31950 3054 32002
rect 3106 31950 3108 32002
rect 2940 31948 3108 31950
rect 3052 31938 3108 31948
rect 3164 32004 3220 32014
rect 2828 31780 2884 31790
rect 2828 31686 2884 31724
rect 3164 31668 3220 31948
rect 2716 31500 3108 31556
rect 3052 30322 3108 31500
rect 3052 30270 3054 30322
rect 3106 30270 3108 30322
rect 3052 30258 3108 30270
rect 3164 30324 3220 31612
rect 3276 31444 3332 32732
rect 3388 32562 3444 32574
rect 3388 32510 3390 32562
rect 3442 32510 3444 32562
rect 3388 32116 3444 32510
rect 3388 32050 3444 32060
rect 3276 31378 3332 31388
rect 3388 31554 3444 31566
rect 3388 31502 3390 31554
rect 3442 31502 3444 31554
rect 3388 31332 3444 31502
rect 3388 31266 3444 31276
rect 3388 30324 3444 30334
rect 3164 30322 3444 30324
rect 3164 30270 3390 30322
rect 3442 30270 3444 30322
rect 3164 30268 3444 30270
rect 3388 30258 3444 30268
rect 2940 30212 2996 30222
rect 2940 30118 2996 30156
rect 3500 30100 3556 33068
rect 3724 33058 3780 33068
rect 3836 33012 3892 33292
rect 4060 33236 4116 33246
rect 5068 33236 5124 33246
rect 4060 33234 4340 33236
rect 4060 33182 4062 33234
rect 4114 33182 4340 33234
rect 4060 33180 4340 33182
rect 4060 33170 4116 33180
rect 3836 32946 3892 32956
rect 3948 33122 4004 33134
rect 3948 33070 3950 33122
rect 4002 33070 4004 33122
rect 3948 32788 4004 33070
rect 4172 33012 4228 33022
rect 3948 32732 4116 32788
rect 3836 32676 3892 32686
rect 3836 32582 3892 32620
rect 3612 32562 3668 32574
rect 3612 32510 3614 32562
rect 3666 32510 3668 32562
rect 3612 31780 3668 32510
rect 3948 32562 4004 32574
rect 3948 32510 3950 32562
rect 4002 32510 4004 32562
rect 3948 32452 4004 32510
rect 3948 32386 4004 32396
rect 3612 31714 3668 31724
rect 3948 32116 4004 32126
rect 3724 31668 3780 31678
rect 3724 31574 3780 31612
rect 3836 31556 3892 31566
rect 3836 31462 3892 31500
rect 3948 31554 4004 32060
rect 3948 31502 3950 31554
rect 4002 31502 4004 31554
rect 3948 30996 4004 31502
rect 4060 31220 4116 32732
rect 4060 31154 4116 31164
rect 4172 31554 4228 32956
rect 4284 31780 4340 33180
rect 5068 33234 5236 33236
rect 5068 33182 5070 33234
rect 5122 33182 5236 33234
rect 5068 33180 5236 33182
rect 5068 33170 5124 33180
rect 4732 33122 4788 33134
rect 4732 33070 4734 33122
rect 4786 33070 4788 33122
rect 4732 32340 4788 33070
rect 4956 33122 5012 33134
rect 4956 33070 4958 33122
rect 5010 33070 5012 33122
rect 4956 32788 5012 33070
rect 4956 32722 5012 32732
rect 5068 32676 5124 32686
rect 4956 32562 5012 32574
rect 4956 32510 4958 32562
rect 5010 32510 5012 32562
rect 4732 32284 4900 32340
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4844 32004 4900 32284
rect 4844 31938 4900 31948
rect 4284 31724 4900 31780
rect 4172 31502 4174 31554
rect 4226 31502 4228 31554
rect 4172 31108 4228 31502
rect 4508 31556 4564 31566
rect 4508 31332 4564 31500
rect 4732 31556 4788 31566
rect 4732 31462 4788 31500
rect 4508 31266 4564 31276
rect 4396 31108 4452 31118
rect 4172 31052 4396 31108
rect 4396 31042 4452 31052
rect 3948 30940 4228 30996
rect 3724 30324 3780 30334
rect 3500 30044 3668 30100
rect 2828 29428 2884 29438
rect 2604 29426 2884 29428
rect 2604 29374 2830 29426
rect 2882 29374 2884 29426
rect 2604 29372 2884 29374
rect 2828 29362 2884 29372
rect 3612 29426 3668 30044
rect 3612 29374 3614 29426
rect 3666 29374 3668 29426
rect 2492 28802 2548 28812
rect 3500 28644 3556 28654
rect 3612 28644 3668 29374
rect 3724 29314 3780 30268
rect 3724 29262 3726 29314
rect 3778 29262 3780 29314
rect 3724 29250 3780 29262
rect 3836 30098 3892 30110
rect 3836 30046 3838 30098
rect 3890 30046 3892 30098
rect 3500 28642 3668 28644
rect 3500 28590 3502 28642
rect 3554 28590 3668 28642
rect 3500 28588 3668 28590
rect 3500 28578 3556 28588
rect 2380 28478 2382 28530
rect 2434 28478 2436 28530
rect 2380 28466 2436 28478
rect 2604 28532 2660 28542
rect 2604 28084 2660 28476
rect 3836 28418 3892 30046
rect 4060 30100 4116 30110
rect 4060 30006 4116 30044
rect 3836 28366 3838 28418
rect 3890 28366 3892 28418
rect 3836 28354 3892 28366
rect 3948 29986 4004 29998
rect 3948 29934 3950 29986
rect 4002 29934 4004 29986
rect 2604 28018 2660 28028
rect 3836 27972 3892 27982
rect 3948 27972 4004 29934
rect 4172 29538 4228 30940
rect 4620 30882 4676 30894
rect 4620 30830 4622 30882
rect 4674 30830 4676 30882
rect 4620 30772 4676 30830
rect 4284 30716 4676 30772
rect 4284 30212 4340 30716
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4844 30436 4900 31724
rect 4956 31668 5012 32510
rect 5068 32450 5124 32620
rect 5068 32398 5070 32450
rect 5122 32398 5124 32450
rect 5068 32386 5124 32398
rect 4956 31602 5012 31612
rect 5068 31554 5124 31566
rect 5068 31502 5070 31554
rect 5122 31502 5124 31554
rect 5068 31444 5124 31502
rect 5068 31378 5124 31388
rect 5180 31220 5236 33180
rect 5292 31444 5348 33740
rect 5628 33572 5684 33582
rect 5628 32900 5684 33516
rect 5628 32450 5684 32844
rect 5740 32562 5796 34076
rect 6300 34066 6356 34076
rect 6076 33908 6132 33918
rect 6076 33570 6132 33852
rect 6076 33518 6078 33570
rect 6130 33518 6132 33570
rect 6076 33506 6132 33518
rect 6412 33572 6468 34636
rect 6636 34626 6692 34636
rect 6860 34354 6916 34860
rect 6860 34302 6862 34354
rect 6914 34302 6916 34354
rect 6860 34290 6916 34302
rect 6412 33506 6468 33516
rect 6524 34242 6580 34254
rect 6524 34190 6526 34242
rect 6578 34190 6580 34242
rect 6524 33348 6580 34190
rect 6412 33292 6580 33348
rect 6636 34130 6692 34142
rect 6636 34078 6638 34130
rect 6690 34078 6692 34130
rect 6636 33908 6692 34078
rect 6636 33348 6692 33852
rect 6636 33292 6804 33348
rect 5740 32510 5742 32562
rect 5794 32510 5796 32562
rect 5740 32498 5796 32510
rect 5852 33122 5908 33134
rect 5852 33070 5854 33122
rect 5906 33070 5908 33122
rect 5628 32398 5630 32450
rect 5682 32398 5684 32450
rect 5628 32386 5684 32398
rect 5852 32340 5908 33070
rect 5964 33122 6020 33134
rect 5964 33070 5966 33122
rect 6018 33070 6020 33122
rect 5964 32676 6020 33070
rect 5964 32610 6020 32620
rect 6300 33122 6356 33134
rect 6300 33070 6302 33122
rect 6354 33070 6356 33122
rect 6076 32394 6132 32416
rect 6076 32342 6078 32394
rect 6130 32342 6132 32394
rect 6076 32340 6132 32342
rect 5852 32284 6132 32340
rect 5964 31780 6020 31790
rect 5852 31668 5908 31678
rect 5852 31574 5908 31612
rect 5964 31554 6020 31724
rect 6076 31668 6132 32284
rect 6076 31602 6132 31612
rect 5964 31502 5966 31554
rect 6018 31502 6020 31554
rect 5964 31490 6020 31502
rect 5292 31378 5348 31388
rect 4956 31164 5236 31220
rect 6076 31220 6132 31230
rect 4956 30772 5012 31164
rect 5180 30996 5236 31006
rect 5180 30902 5236 30940
rect 6076 30994 6132 31164
rect 6076 30942 6078 30994
rect 6130 30942 6132 30994
rect 5292 30884 5348 30894
rect 5292 30882 5572 30884
rect 5292 30830 5294 30882
rect 5346 30830 5572 30882
rect 5292 30828 5572 30830
rect 5292 30818 5348 30828
rect 4956 30716 5236 30772
rect 4284 30146 4340 30156
rect 4732 30380 4900 30436
rect 4172 29486 4174 29538
rect 4226 29486 4228 29538
rect 4172 29474 4228 29486
rect 4508 29986 4564 29998
rect 4508 29934 4510 29986
rect 4562 29934 4564 29986
rect 4508 29204 4564 29934
rect 3836 27970 4004 27972
rect 3836 27918 3838 27970
rect 3890 27918 4004 27970
rect 3836 27916 4004 27918
rect 4172 29148 4564 29204
rect 4732 29204 4788 30380
rect 4956 30324 5012 30334
rect 4956 30230 5012 30268
rect 4844 30212 4900 30222
rect 4844 29538 4900 30156
rect 5068 29540 5124 29550
rect 4844 29486 4846 29538
rect 4898 29486 4900 29538
rect 4844 29474 4900 29486
rect 4956 29538 5124 29540
rect 4956 29486 5070 29538
rect 5122 29486 5124 29538
rect 4956 29484 5124 29486
rect 3836 27906 3892 27916
rect 3500 27860 3556 27870
rect 3164 26962 3220 26974
rect 3164 26910 3166 26962
rect 3218 26910 3220 26962
rect 1932 26852 2212 26908
rect 2268 26852 2436 26908
rect 2156 25620 2212 26852
rect 2156 25554 2212 25564
rect 2268 26290 2324 26302
rect 2268 26238 2270 26290
rect 2322 26238 2324 26290
rect 1820 25454 1822 25506
rect 1874 25454 1876 25506
rect 1820 25442 1876 25454
rect 2156 25172 2212 25182
rect 2156 24946 2212 25116
rect 2156 24894 2158 24946
rect 2210 24894 2212 24946
rect 2156 24882 2212 24894
rect 2268 24948 2324 26238
rect 2380 25620 2436 26852
rect 2492 26852 2548 26862
rect 2492 26850 2660 26852
rect 2492 26798 2494 26850
rect 2546 26798 2660 26850
rect 2492 26796 2660 26798
rect 2492 26786 2548 26796
rect 2492 25620 2548 25630
rect 2380 25618 2548 25620
rect 2380 25566 2494 25618
rect 2546 25566 2548 25618
rect 2380 25564 2548 25566
rect 2492 25554 2548 25564
rect 2268 24892 2436 24948
rect 2268 24722 2324 24734
rect 2268 24670 2270 24722
rect 2322 24670 2324 24722
rect 1820 23154 1876 23166
rect 1820 23102 1822 23154
rect 1874 23102 1876 23154
rect 1820 22932 1876 23102
rect 1820 22876 2100 22932
rect 1820 22484 1876 22494
rect 1708 22482 1876 22484
rect 1708 22430 1822 22482
rect 1874 22430 1876 22482
rect 1708 22428 1876 22430
rect 1708 19348 1764 19358
rect 1708 19254 1764 19292
rect 1820 18116 1876 22428
rect 2044 21700 2100 22876
rect 1932 21476 1988 21486
rect 1932 21382 1988 21420
rect 2044 20802 2100 21644
rect 2268 21476 2324 24670
rect 2380 24164 2436 24892
rect 2604 24946 2660 26796
rect 3052 26290 3108 26302
rect 3052 26238 3054 26290
rect 3106 26238 3108 26290
rect 2940 26180 2996 26190
rect 2604 24894 2606 24946
rect 2658 24894 2660 24946
rect 2380 24162 2548 24164
rect 2380 24110 2382 24162
rect 2434 24110 2548 24162
rect 2380 24108 2548 24110
rect 2380 24098 2436 24108
rect 2492 23492 2548 24108
rect 2604 23940 2660 24894
rect 2828 26178 2996 26180
rect 2828 26126 2942 26178
rect 2994 26126 2996 26178
rect 2828 26124 2996 26126
rect 2716 24724 2772 24734
rect 2716 24630 2772 24668
rect 2828 24388 2884 26124
rect 2940 26114 2996 26124
rect 2940 24836 2996 24846
rect 2940 24742 2996 24780
rect 2604 23874 2660 23884
rect 2716 24332 2884 24388
rect 2492 23426 2548 23436
rect 2380 23380 2436 23390
rect 2380 22370 2436 23324
rect 2492 23044 2548 23054
rect 2492 23042 2660 23044
rect 2492 22990 2494 23042
rect 2546 22990 2660 23042
rect 2492 22988 2660 22990
rect 2492 22978 2548 22988
rect 2380 22318 2382 22370
rect 2434 22318 2436 22370
rect 2380 22306 2436 22318
rect 2324 21420 2548 21476
rect 2268 21410 2324 21420
rect 2044 20750 2046 20802
rect 2098 20750 2100 20802
rect 2044 20738 2100 20750
rect 2492 20244 2548 21420
rect 2268 20242 2548 20244
rect 2268 20190 2494 20242
rect 2546 20190 2548 20242
rect 2268 20188 2548 20190
rect 2156 19908 2212 19918
rect 2156 19814 2212 19852
rect 1820 18050 1876 18060
rect 1932 19460 1988 19470
rect 1932 17778 1988 19404
rect 1932 17726 1934 17778
rect 1986 17726 1988 17778
rect 1932 17714 1988 17726
rect 2044 18452 2100 18462
rect 1708 17108 1764 17118
rect 1596 17106 1764 17108
rect 1596 17054 1710 17106
rect 1762 17054 1764 17106
rect 1596 17052 1764 17054
rect 1260 16940 1540 16996
rect 1148 15372 1316 15428
rect 1260 15316 1316 15372
rect 1260 15260 1428 15316
rect 1036 15138 1092 15148
rect 1372 14420 1428 15260
rect 1372 14354 1428 14364
rect 1484 13972 1540 16940
rect 1484 13906 1540 13916
rect 1708 7700 1764 17052
rect 2044 16212 2100 18396
rect 2268 17666 2324 20188
rect 2492 20178 2548 20188
rect 2268 17614 2270 17666
rect 2322 17614 2324 17666
rect 2268 17602 2324 17614
rect 2380 19012 2436 19022
rect 2268 16884 2324 16894
rect 2268 16790 2324 16828
rect 2156 16212 2212 16222
rect 2044 16210 2212 16212
rect 2044 16158 2158 16210
rect 2210 16158 2212 16210
rect 2044 16156 2212 16158
rect 2156 15538 2212 16156
rect 2380 15876 2436 18956
rect 2492 18452 2548 18462
rect 2492 18358 2548 18396
rect 2604 17108 2660 22988
rect 2716 20916 2772 24332
rect 2828 24164 2884 24174
rect 2828 22482 2884 24108
rect 3052 24052 3108 26238
rect 3164 24164 3220 26910
rect 3388 24724 3444 24734
rect 3388 24630 3444 24668
rect 3164 24098 3220 24108
rect 3052 23986 3108 23996
rect 3164 23716 3220 23726
rect 3500 23716 3556 27804
rect 4172 27860 4228 29148
rect 4732 29138 4788 29148
rect 4844 29316 4900 29326
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4508 28868 4564 28878
rect 4508 28774 4564 28812
rect 4844 28866 4900 29260
rect 4844 28814 4846 28866
rect 4898 28814 4900 28866
rect 4844 28802 4900 28814
rect 4172 27794 4228 27804
rect 4284 28644 4340 28654
rect 3220 23660 3556 23716
rect 3612 27074 3668 27086
rect 3612 27022 3614 27074
rect 3666 27022 3668 27074
rect 3164 22596 3220 23660
rect 3612 23380 3668 27022
rect 4172 26962 4228 26974
rect 4172 26910 4174 26962
rect 4226 26910 4228 26962
rect 4172 26908 4228 26910
rect 4060 26852 4228 26908
rect 4284 26908 4340 28588
rect 4508 28532 4564 28542
rect 4508 27858 4564 28476
rect 4508 27806 4510 27858
rect 4562 27806 4564 27858
rect 4508 27794 4564 27806
rect 4844 27972 4900 27982
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4844 26962 4900 27916
rect 4844 26910 4846 26962
rect 4898 26910 4900 26962
rect 4284 26852 4564 26908
rect 4844 26898 4900 26910
rect 4060 26516 4116 26852
rect 4508 26850 4564 26852
rect 4508 26798 4510 26850
rect 4562 26798 4564 26850
rect 4508 26786 4564 26798
rect 4732 26516 4788 26526
rect 4060 26514 4788 26516
rect 4060 26462 4734 26514
rect 4786 26462 4788 26514
rect 4060 26460 4788 26462
rect 3836 24836 3892 24846
rect 3836 24742 3892 24780
rect 3612 23314 3668 23324
rect 3724 24724 3780 24734
rect 3388 22596 3444 22606
rect 3164 22594 3444 22596
rect 3164 22542 3390 22594
rect 3442 22542 3444 22594
rect 3164 22540 3444 22542
rect 3388 22530 3444 22540
rect 2828 22430 2830 22482
rect 2882 22430 2884 22482
rect 2828 22418 2884 22430
rect 2716 20850 2772 20860
rect 2940 22370 2996 22382
rect 2940 22318 2942 22370
rect 2994 22318 2996 22370
rect 2716 20690 2772 20702
rect 2716 20638 2718 20690
rect 2770 20638 2772 20690
rect 2716 18788 2772 20638
rect 2716 18722 2772 18732
rect 2940 19348 2996 22318
rect 3276 21028 3332 21038
rect 3276 20242 3332 20972
rect 3276 20190 3278 20242
rect 3330 20190 3332 20242
rect 3276 20178 3332 20190
rect 3724 19908 3780 24668
rect 3948 23492 4004 23502
rect 3948 22484 4004 23436
rect 3948 22390 4004 22428
rect 4060 22260 4116 26460
rect 4732 26450 4788 26460
rect 4844 26516 4900 26526
rect 4172 26290 4228 26302
rect 4172 26238 4174 26290
rect 4226 26238 4228 26290
rect 4172 22372 4228 26238
rect 4620 26292 4676 26302
rect 4620 26198 4676 26236
rect 4732 26068 4788 26078
rect 4844 26068 4900 26460
rect 4732 26066 4900 26068
rect 4732 26014 4734 26066
rect 4786 26014 4900 26066
rect 4732 26012 4900 26014
rect 4732 26002 4788 26012
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4620 25620 4676 25630
rect 4620 25526 4676 25564
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4284 24164 4340 24174
rect 4284 23938 4340 24108
rect 4956 24050 5012 29484
rect 5068 29474 5124 29484
rect 5180 29316 5236 30716
rect 5292 29540 5348 29550
rect 5292 29446 5348 29484
rect 5180 29260 5348 29316
rect 5068 29204 5124 29214
rect 5124 29148 5236 29204
rect 5068 29138 5124 29148
rect 5068 28642 5124 28654
rect 5068 28590 5070 28642
rect 5122 28590 5124 28642
rect 5068 28532 5124 28590
rect 5068 28466 5124 28476
rect 5180 27970 5236 29148
rect 5292 28082 5348 29260
rect 5292 28030 5294 28082
rect 5346 28030 5348 28082
rect 5292 28018 5348 28030
rect 5516 28196 5572 30828
rect 6076 30324 6132 30942
rect 6076 30258 6132 30268
rect 5852 30212 5908 30222
rect 5908 30156 6020 30212
rect 5852 30146 5908 30156
rect 5852 29988 5908 29998
rect 5740 29986 5908 29988
rect 5740 29934 5854 29986
rect 5906 29934 5908 29986
rect 5740 29932 5908 29934
rect 5628 29204 5684 29214
rect 5628 29110 5684 29148
rect 5180 27918 5182 27970
rect 5234 27918 5236 27970
rect 5180 27636 5236 27918
rect 5180 27570 5236 27580
rect 5404 27634 5460 27646
rect 5404 27582 5406 27634
rect 5458 27582 5460 27634
rect 5068 27188 5124 27198
rect 5068 27074 5124 27132
rect 5068 27022 5070 27074
rect 5122 27022 5124 27074
rect 5068 27010 5124 27022
rect 5404 27076 5460 27582
rect 5404 27010 5460 27020
rect 5516 26964 5572 28140
rect 5740 26908 5796 29932
rect 5852 29922 5908 29932
rect 5852 28980 5908 28990
rect 5852 28642 5908 28924
rect 5852 28590 5854 28642
rect 5906 28590 5908 28642
rect 5852 28578 5908 28590
rect 5964 28082 6020 30156
rect 6300 29988 6356 33070
rect 6412 31668 6468 33292
rect 6636 33178 6692 33190
rect 6412 31602 6468 31612
rect 6524 33122 6580 33134
rect 6524 33070 6526 33122
rect 6578 33070 6580 33122
rect 6524 31220 6580 33070
rect 6524 31154 6580 31164
rect 6636 33126 6638 33178
rect 6690 33126 6692 33178
rect 6524 30996 6580 31006
rect 6524 30902 6580 30940
rect 6524 30772 6580 30782
rect 6188 29932 6356 29988
rect 6412 30098 6468 30110
rect 6412 30046 6414 30098
rect 6466 30046 6468 30098
rect 6076 29428 6132 29438
rect 6076 29334 6132 29372
rect 6076 28644 6132 28654
rect 6076 28550 6132 28588
rect 6188 28418 6244 29932
rect 6300 29428 6356 29438
rect 6412 29428 6468 30046
rect 6524 29650 6580 30716
rect 6636 30212 6692 33126
rect 6748 31780 6804 33292
rect 6972 32676 7028 35084
rect 7196 34916 7252 34926
rect 7084 34242 7140 34254
rect 7084 34190 7086 34242
rect 7138 34190 7140 34242
rect 7084 34132 7140 34190
rect 7196 34242 7252 34860
rect 7308 34802 7364 35084
rect 7308 34750 7310 34802
rect 7362 34750 7364 34802
rect 7308 34738 7364 34750
rect 7420 34690 7476 34702
rect 7420 34638 7422 34690
rect 7474 34638 7476 34690
rect 7420 34580 7476 34638
rect 7420 34514 7476 34524
rect 7532 34356 7588 35644
rect 7868 35476 7924 38612
rect 8316 38162 8372 38612
rect 8316 38110 8318 38162
rect 8370 38110 8372 38162
rect 8316 38098 8372 38110
rect 7644 35420 7924 35476
rect 7980 38052 8036 38062
rect 7980 35698 8036 37996
rect 8652 37938 8708 38892
rect 8652 37886 8654 37938
rect 8706 37886 8708 37938
rect 8652 37874 8708 37886
rect 8876 38722 8932 38734
rect 8876 38670 8878 38722
rect 8930 38670 8932 38722
rect 8764 37828 8820 37838
rect 8428 37380 8484 37390
rect 8428 37266 8484 37324
rect 8764 37268 8820 37772
rect 8428 37214 8430 37266
rect 8482 37214 8484 37266
rect 8428 37202 8484 37214
rect 8652 37266 8820 37268
rect 8652 37214 8766 37266
rect 8818 37214 8820 37266
rect 8652 37212 8820 37214
rect 8428 36708 8484 36718
rect 7980 35646 7982 35698
rect 8034 35646 8036 35698
rect 7644 34914 7700 35420
rect 7980 35028 8036 35646
rect 7644 34862 7646 34914
rect 7698 34862 7700 34914
rect 7644 34850 7700 34862
rect 7756 34972 8036 35028
rect 8092 36706 8484 36708
rect 8092 36654 8430 36706
rect 8482 36654 8484 36706
rect 8092 36652 8484 36654
rect 8092 36148 8148 36652
rect 8428 36642 8484 36652
rect 8204 36484 8260 36522
rect 8260 36428 8596 36484
rect 8204 36418 8260 36428
rect 7756 34356 7812 34972
rect 7868 34804 7924 34814
rect 8092 34804 8148 36092
rect 8204 36260 8260 36270
rect 8204 35308 8260 36204
rect 8540 35922 8596 36428
rect 8652 36260 8708 37212
rect 8764 37202 8820 37212
rect 8876 36820 8932 38670
rect 8988 37828 9044 37838
rect 9100 37828 9156 40348
rect 8988 37826 9156 37828
rect 8988 37774 8990 37826
rect 9042 37774 9156 37826
rect 8988 37772 9156 37774
rect 9212 39394 9268 39406
rect 9212 39342 9214 39394
rect 9266 39342 9268 39394
rect 9212 39060 9268 39342
rect 9324 39396 9380 40910
rect 9548 40514 9604 42140
rect 9548 40462 9550 40514
rect 9602 40462 9604 40514
rect 9548 39508 9604 40462
rect 9660 41972 9716 41982
rect 9660 39732 9716 41916
rect 9772 41858 9828 42364
rect 9772 41806 9774 41858
rect 9826 41806 9828 41858
rect 9772 41794 9828 41806
rect 9772 40964 9828 40974
rect 9884 40964 9940 42476
rect 10220 41970 10276 41982
rect 10220 41918 10222 41970
rect 10274 41918 10276 41970
rect 10108 41858 10164 41870
rect 10108 41806 10110 41858
rect 10162 41806 10164 41858
rect 10108 41748 10164 41806
rect 10108 41682 10164 41692
rect 10220 41188 10276 41918
rect 10220 41122 10276 41132
rect 9828 40908 9940 40964
rect 10108 40964 10164 40974
rect 10332 40964 10388 42588
rect 10668 41300 10724 41310
rect 10668 41206 10724 41244
rect 10556 40964 10612 40974
rect 10780 40964 10836 42924
rect 11340 42868 11396 43262
rect 11788 43426 11844 43438
rect 11788 43374 11790 43426
rect 11842 43374 11844 43426
rect 11788 43092 11844 43374
rect 12236 43426 12292 43438
rect 12236 43374 12238 43426
rect 12290 43374 12292 43426
rect 12236 43314 12292 43374
rect 12460 43428 12516 43596
rect 13244 43540 13300 43550
rect 13356 43540 13412 43820
rect 13916 43652 13972 43662
rect 13916 43558 13972 43596
rect 14028 43652 14084 43662
rect 14028 43650 14196 43652
rect 14028 43598 14030 43650
rect 14082 43598 14196 43650
rect 14028 43596 14196 43598
rect 14028 43586 14084 43596
rect 13244 43538 13412 43540
rect 13244 43486 13246 43538
rect 13298 43486 13412 43538
rect 13244 43484 13412 43486
rect 13580 43538 13636 43550
rect 13580 43486 13582 43538
rect 13634 43486 13636 43538
rect 13244 43474 13300 43484
rect 12460 43372 12964 43428
rect 12236 43262 12238 43314
rect 12290 43262 12292 43314
rect 12236 43250 12292 43262
rect 11788 43026 11844 43036
rect 11340 42812 11620 42868
rect 11452 42642 11508 42654
rect 11452 42590 11454 42642
rect 11506 42590 11508 42642
rect 10108 40962 10612 40964
rect 10108 40910 10110 40962
rect 10162 40910 10558 40962
rect 10610 40910 10612 40962
rect 10108 40908 10612 40910
rect 9772 40870 9828 40908
rect 10108 40898 10164 40908
rect 10556 40898 10612 40908
rect 10668 40962 10836 40964
rect 10668 40910 10782 40962
rect 10834 40910 10836 40962
rect 10668 40908 10836 40910
rect 10668 40852 10724 40908
rect 10780 40898 10836 40908
rect 11004 41356 11284 41412
rect 10668 40786 10724 40796
rect 11004 40740 11060 41356
rect 10780 40684 11060 40740
rect 11116 41186 11172 41198
rect 11116 41134 11118 41186
rect 11170 41134 11172 41186
rect 10108 40626 10164 40638
rect 10108 40574 10110 40626
rect 10162 40574 10164 40626
rect 10108 40516 10164 40574
rect 10108 40450 10164 40460
rect 10780 40514 10836 40684
rect 11116 40626 11172 41134
rect 11228 41188 11284 41356
rect 11340 41188 11396 41198
rect 11228 41186 11396 41188
rect 11228 41134 11342 41186
rect 11394 41134 11396 41186
rect 11228 41132 11396 41134
rect 11340 41122 11396 41132
rect 11116 40574 11118 40626
rect 11170 40574 11172 40626
rect 11116 40562 11172 40574
rect 11452 40628 11508 42590
rect 11564 41858 11620 42812
rect 11676 42642 11732 42654
rect 11676 42590 11678 42642
rect 11730 42590 11732 42642
rect 11676 42196 11732 42590
rect 11676 42130 11732 42140
rect 12012 42642 12068 42654
rect 12012 42590 12014 42642
rect 12066 42590 12068 42642
rect 11564 41806 11566 41858
rect 11618 41806 11620 41858
rect 11564 41412 11620 41806
rect 11564 41346 11620 41356
rect 11788 41746 11844 41758
rect 11788 41694 11790 41746
rect 11842 41694 11844 41746
rect 11676 41074 11732 41086
rect 11676 41022 11678 41074
rect 11730 41022 11732 41074
rect 11564 40962 11620 40974
rect 11564 40910 11566 40962
rect 11618 40910 11620 40962
rect 11564 40852 11620 40910
rect 11676 40964 11732 41022
rect 11788 40964 11844 41694
rect 12012 41300 12068 42590
rect 12796 42644 12852 42654
rect 12124 42532 12180 42542
rect 12124 42194 12180 42476
rect 12124 42142 12126 42194
rect 12178 42142 12180 42194
rect 12124 42130 12180 42142
rect 12348 42530 12404 42542
rect 12348 42478 12350 42530
rect 12402 42478 12404 42530
rect 12012 41234 12068 41244
rect 12348 41188 12404 42478
rect 12572 42530 12628 42542
rect 12572 42478 12574 42530
rect 12626 42478 12628 42530
rect 12348 41122 12404 41132
rect 12460 41412 12516 41422
rect 12460 41186 12516 41356
rect 12460 41134 12462 41186
rect 12514 41134 12516 41186
rect 12460 41122 12516 41134
rect 12236 40964 12292 40974
rect 11788 40908 12180 40964
rect 11676 40898 11732 40908
rect 11564 40786 11620 40796
rect 12124 40740 12180 40908
rect 12236 40870 12292 40908
rect 12572 40740 12628 42478
rect 12684 41858 12740 41870
rect 12684 41806 12686 41858
rect 12738 41806 12740 41858
rect 12684 41300 12740 41806
rect 12684 41234 12740 41244
rect 12796 41074 12852 42588
rect 12908 42642 12964 43372
rect 13580 43092 13636 43486
rect 14140 43540 14196 43596
rect 14028 43316 14084 43326
rect 13580 43026 13636 43036
rect 13692 43314 14084 43316
rect 13692 43262 14030 43314
rect 14082 43262 14084 43314
rect 13692 43260 14084 43262
rect 12908 42590 12910 42642
rect 12962 42590 12964 42642
rect 12908 42578 12964 42590
rect 13692 42754 13748 43260
rect 14028 43250 14084 43260
rect 14140 42866 14196 43484
rect 14140 42814 14142 42866
rect 14194 42814 14196 42866
rect 13692 42702 13694 42754
rect 13746 42702 13748 42754
rect 13356 42532 13412 42542
rect 13132 42530 13412 42532
rect 13132 42478 13358 42530
rect 13410 42478 13412 42530
rect 13132 42476 13412 42478
rect 13132 41970 13188 42476
rect 13356 42466 13412 42476
rect 13580 42532 13636 42542
rect 13580 42438 13636 42476
rect 13132 41918 13134 41970
rect 13186 41918 13188 41970
rect 13132 41906 13188 41918
rect 13468 41748 13524 41758
rect 13468 41654 13524 41692
rect 13468 41188 13524 41198
rect 13468 41094 13524 41132
rect 12796 41022 12798 41074
rect 12850 41022 12852 41074
rect 12796 41010 12852 41022
rect 13692 41074 13748 42702
rect 13916 42756 13972 42766
rect 13916 41858 13972 42700
rect 14140 42644 14196 42814
rect 14140 42578 14196 42588
rect 13916 41806 13918 41858
rect 13970 41806 13972 41858
rect 13916 41794 13972 41806
rect 14476 41300 14532 45052
rect 14588 45042 14644 45052
rect 14700 44996 14756 45006
rect 14700 44994 14868 44996
rect 14700 44942 14702 44994
rect 14754 44942 14868 44994
rect 14700 44940 14868 44942
rect 14700 44930 14756 44940
rect 14812 43762 14868 44940
rect 15372 44548 15428 44558
rect 15372 44454 15428 44492
rect 16044 44322 16100 45950
rect 16156 44548 16212 49200
rect 17724 46004 17780 49200
rect 19180 46116 19236 46126
rect 19292 46116 19348 49200
rect 19180 46114 19348 46116
rect 19180 46062 19182 46114
rect 19234 46062 19348 46114
rect 19180 46060 19348 46062
rect 20860 46116 20916 49200
rect 19180 46050 19236 46060
rect 20860 46050 20916 46060
rect 22092 46116 22148 46126
rect 22092 46022 22148 46060
rect 22428 46116 22484 49200
rect 23996 46788 24052 49200
rect 25564 49140 25620 49200
rect 25900 49140 25956 49308
rect 25564 49084 25956 49140
rect 22428 46050 22484 46060
rect 23548 46732 24052 46788
rect 17724 45948 17892 46004
rect 16940 45780 16996 45790
rect 16940 45686 16996 45724
rect 17500 45108 17556 45118
rect 17500 45014 17556 45052
rect 16828 44994 16884 45006
rect 16828 44942 16830 44994
rect 16882 44942 16884 44994
rect 16828 44548 16884 44942
rect 16828 44492 17780 44548
rect 16156 44482 16212 44492
rect 16044 44270 16046 44322
rect 16098 44270 16100 44322
rect 16044 44258 16100 44270
rect 16828 44322 16884 44334
rect 16828 44270 16830 44322
rect 16882 44270 16884 44322
rect 16828 44100 16884 44270
rect 17500 44212 17556 44222
rect 16828 44034 16884 44044
rect 17276 44210 17556 44212
rect 17276 44158 17502 44210
rect 17554 44158 17556 44210
rect 17276 44156 17556 44158
rect 14812 43710 14814 43762
rect 14866 43710 14868 43762
rect 14812 43698 14868 43710
rect 14700 43652 14756 43662
rect 14700 43558 14756 43596
rect 15372 43652 15428 43662
rect 15372 43558 15428 43596
rect 15260 43540 15316 43550
rect 15260 43446 15316 43484
rect 15484 43538 15540 43550
rect 15484 43486 15486 43538
rect 15538 43486 15540 43538
rect 14924 43428 14980 43438
rect 14924 43334 14980 43372
rect 15484 43316 15540 43486
rect 14588 42756 14644 42766
rect 14588 42662 14644 42700
rect 15484 42756 15540 43260
rect 15484 42690 15540 42700
rect 15708 43538 15764 43550
rect 15708 43486 15710 43538
rect 15762 43486 15764 43538
rect 15708 42980 15764 43486
rect 16156 43540 16212 43550
rect 16156 43446 16212 43484
rect 16380 43538 16436 43550
rect 16380 43486 16382 43538
rect 16434 43486 16436 43538
rect 16268 43428 16324 43438
rect 16268 43334 16324 43372
rect 16380 43316 16436 43486
rect 16828 43540 16884 43550
rect 16828 43538 16996 43540
rect 16828 43486 16830 43538
rect 16882 43486 16996 43538
rect 16828 43484 16996 43486
rect 16828 43474 16884 43484
rect 16380 43250 16436 43260
rect 16940 43316 16996 43484
rect 15708 42754 15764 42924
rect 15708 42702 15710 42754
rect 15762 42702 15764 42754
rect 15708 42690 15764 42702
rect 16156 42642 16212 42654
rect 16156 42590 16158 42642
rect 16210 42590 16212 42642
rect 16044 41860 16100 41870
rect 15932 41858 16100 41860
rect 15932 41806 16046 41858
rect 16098 41806 16100 41858
rect 15932 41804 16100 41806
rect 14588 41300 14644 41310
rect 13692 41022 13694 41074
rect 13746 41022 13748 41074
rect 13692 41010 13748 41022
rect 14140 41298 14644 41300
rect 14140 41246 14590 41298
rect 14642 41246 14644 41298
rect 14140 41244 14644 41246
rect 14028 40962 14084 40974
rect 14028 40910 14030 40962
rect 14082 40910 14084 40962
rect 12124 40684 12628 40740
rect 12684 40740 12740 40750
rect 11676 40628 11732 40638
rect 11452 40626 11732 40628
rect 11452 40574 11678 40626
rect 11730 40574 11732 40626
rect 11452 40572 11732 40574
rect 11676 40562 11732 40572
rect 10780 40462 10782 40514
rect 10834 40462 10836 40514
rect 10780 40450 10836 40462
rect 10892 40516 10948 40526
rect 9884 40404 9940 40414
rect 9772 40180 9828 40190
rect 9772 40086 9828 40124
rect 9884 39956 9940 40348
rect 9660 39638 9716 39676
rect 9772 39900 9940 39956
rect 9996 40180 10052 40190
rect 10892 40180 10948 40460
rect 11004 40514 11060 40526
rect 11004 40462 11006 40514
rect 11058 40462 11060 40514
rect 11004 40404 11060 40462
rect 12012 40516 12068 40526
rect 12012 40422 12068 40460
rect 11004 40338 11060 40348
rect 11228 40404 11284 40414
rect 11564 40404 11620 40414
rect 11228 40402 11620 40404
rect 11228 40350 11230 40402
rect 11282 40350 11566 40402
rect 11618 40350 11620 40402
rect 11228 40348 11620 40350
rect 11228 40338 11284 40348
rect 10892 40124 11172 40180
rect 9548 39442 9604 39452
rect 9324 39330 9380 39340
rect 8988 37380 9044 37772
rect 8988 37314 9044 37324
rect 9100 37604 9156 37614
rect 8988 37156 9044 37166
rect 9100 37156 9156 37548
rect 8988 37154 9156 37156
rect 8988 37102 8990 37154
rect 9042 37102 9156 37154
rect 8988 37100 9156 37102
rect 8988 37090 9044 37100
rect 8876 36754 8932 36764
rect 9212 36708 9268 39004
rect 9660 38948 9716 38958
rect 9660 38854 9716 38892
rect 9548 38834 9604 38846
rect 9548 38782 9550 38834
rect 9602 38782 9604 38834
rect 9548 38724 9604 38782
rect 9772 38668 9828 39900
rect 9996 39506 10052 40124
rect 10780 39732 10836 39742
rect 9996 39454 9998 39506
rect 10050 39454 10052 39506
rect 9996 39442 10052 39454
rect 10332 39508 10388 39518
rect 10332 39414 10388 39452
rect 9884 39396 9940 39406
rect 9884 39058 9940 39340
rect 9884 39006 9886 39058
rect 9938 39006 9940 39058
rect 9884 38994 9940 39006
rect 10220 39116 10724 39172
rect 10108 38836 10164 38846
rect 9548 38612 9716 38668
rect 9772 38612 9940 38668
rect 9660 37938 9716 38612
rect 9660 37886 9662 37938
rect 9714 37886 9716 37938
rect 9660 37874 9716 37886
rect 9324 37828 9380 37838
rect 9324 37734 9380 37772
rect 9548 37828 9604 37838
rect 9548 36932 9604 37772
rect 9100 36652 9268 36708
rect 9324 36876 9604 36932
rect 9660 37604 9716 37614
rect 8764 36594 8820 36606
rect 8764 36542 8766 36594
rect 8818 36542 8820 36594
rect 8764 36484 8820 36542
rect 8764 36418 8820 36428
rect 8652 36194 8708 36204
rect 9100 35924 9156 36652
rect 9212 36484 9268 36494
rect 9212 36390 9268 36428
rect 8540 35870 8542 35922
rect 8594 35870 8596 35922
rect 8540 35858 8596 35870
rect 8652 35868 9156 35924
rect 8540 35476 8596 35486
rect 8204 35252 8484 35308
rect 7868 34802 8148 34804
rect 7868 34750 7870 34802
rect 7922 34750 8148 34802
rect 7868 34748 8148 34750
rect 8204 34804 8260 34814
rect 7868 34738 7924 34748
rect 7196 34190 7198 34242
rect 7250 34190 7252 34242
rect 7196 34178 7252 34190
rect 7308 34300 7588 34356
rect 7644 34300 7812 34356
rect 8204 34690 8260 34748
rect 8204 34638 8206 34690
rect 8258 34638 8260 34690
rect 7084 34066 7140 34076
rect 7308 33908 7364 34300
rect 7196 33852 7364 33908
rect 6972 32610 7028 32620
rect 7084 33234 7140 33246
rect 7084 33182 7086 33234
rect 7138 33182 7140 33234
rect 6972 31780 7028 31790
rect 6748 31778 7028 31780
rect 6748 31726 6974 31778
rect 7026 31726 7028 31778
rect 6748 31724 7028 31726
rect 6972 31714 7028 31724
rect 7084 31780 7140 33182
rect 7196 32900 7252 33852
rect 7644 33796 7700 34300
rect 7868 34244 7924 34254
rect 7868 34242 8036 34244
rect 7868 34190 7870 34242
rect 7922 34190 8036 34242
rect 7868 34188 8036 34190
rect 7868 34178 7924 34188
rect 7756 34130 7812 34142
rect 7756 34078 7758 34130
rect 7810 34078 7812 34130
rect 7756 34020 7812 34078
rect 7756 33954 7812 33964
rect 7308 33740 7700 33796
rect 7308 33012 7364 33740
rect 7420 33572 7476 33582
rect 7420 33570 7924 33572
rect 7420 33518 7422 33570
rect 7474 33518 7924 33570
rect 7420 33516 7924 33518
rect 7420 33506 7476 33516
rect 7420 33346 7476 33358
rect 7420 33294 7422 33346
rect 7474 33294 7476 33346
rect 7420 33236 7476 33294
rect 7420 33170 7476 33180
rect 7308 32956 7476 33012
rect 7196 32844 7364 32900
rect 7084 31714 7140 31724
rect 7196 31668 7252 31706
rect 7196 31602 7252 31612
rect 6860 31556 6916 31566
rect 6860 31218 6916 31500
rect 6860 31166 6862 31218
rect 6914 31166 6916 31218
rect 6860 31108 6916 31166
rect 7196 31444 7252 31454
rect 7196 31218 7252 31388
rect 7196 31166 7198 31218
rect 7250 31166 7252 31218
rect 7196 31154 7252 31166
rect 6860 31042 6916 31052
rect 6636 30146 6692 30156
rect 6972 30996 7028 31006
rect 6972 30098 7028 30940
rect 7084 30212 7140 30222
rect 7084 30118 7140 30156
rect 7308 30210 7364 32844
rect 7420 31556 7476 32956
rect 7868 32788 7924 33516
rect 7980 33460 8036 34188
rect 8092 34132 8148 34142
rect 8092 34038 8148 34076
rect 8204 33684 8260 34638
rect 8316 34018 8372 34030
rect 8316 33966 8318 34018
rect 8370 33966 8372 34018
rect 8316 33908 8372 33966
rect 8316 33842 8372 33852
rect 8204 33628 8372 33684
rect 7980 33366 8036 33404
rect 7868 32732 8260 32788
rect 8204 32674 8260 32732
rect 8204 32622 8206 32674
rect 8258 32622 8260 32674
rect 8204 32610 8260 32622
rect 8316 32452 8372 33628
rect 7420 31490 7476 31500
rect 7756 32396 8372 32452
rect 7532 31332 7588 31342
rect 7308 30158 7310 30210
rect 7362 30158 7364 30210
rect 7308 30146 7364 30158
rect 7420 31276 7532 31332
rect 6972 30046 6974 30098
rect 7026 30046 7028 30098
rect 6524 29598 6526 29650
rect 6578 29598 6580 29650
rect 6524 29586 6580 29598
rect 6636 29764 6692 29774
rect 6636 29428 6692 29708
rect 6972 29538 7028 30046
rect 6972 29486 6974 29538
rect 7026 29486 7028 29538
rect 6972 29474 7028 29486
rect 6300 29426 6468 29428
rect 6300 29374 6302 29426
rect 6354 29374 6468 29426
rect 6300 29372 6468 29374
rect 6524 29372 6692 29428
rect 6748 29426 6804 29438
rect 6748 29374 6750 29426
rect 6802 29374 6804 29426
rect 6300 28756 6356 29372
rect 6300 28690 6356 28700
rect 6524 28644 6580 29372
rect 6748 29204 6804 29374
rect 7196 29204 7252 29214
rect 6524 28578 6580 28588
rect 6636 29202 7252 29204
rect 6636 29150 7198 29202
rect 7250 29150 7252 29202
rect 6636 29148 7252 29150
rect 6188 28366 6190 28418
rect 6242 28366 6244 28418
rect 6188 28354 6244 28366
rect 5964 28030 5966 28082
rect 6018 28030 6020 28082
rect 5964 28018 6020 28030
rect 6076 28196 6132 28206
rect 6076 27970 6132 28140
rect 6076 27918 6078 27970
rect 6130 27918 6132 27970
rect 6076 27906 6132 27918
rect 6524 27188 6580 27198
rect 6636 27188 6692 29148
rect 6972 28642 7028 29148
rect 7196 29138 7252 29148
rect 7420 28980 7476 31276
rect 7532 31266 7588 31276
rect 7644 30436 7700 30446
rect 7756 30436 7812 32396
rect 8428 32228 8484 35252
rect 8540 34580 8596 35420
rect 8540 34514 8596 34524
rect 8428 32162 8484 32172
rect 8540 32116 8596 32126
rect 8092 31948 8372 32004
rect 7868 31220 7924 31230
rect 7868 31108 7924 31164
rect 7868 31106 8036 31108
rect 7868 31054 7870 31106
rect 7922 31054 8036 31106
rect 7868 31052 8036 31054
rect 7868 31042 7924 31052
rect 7644 30434 7812 30436
rect 7644 30382 7646 30434
rect 7698 30382 7812 30434
rect 7644 30380 7812 30382
rect 7980 30434 8036 31052
rect 7980 30382 7982 30434
rect 8034 30382 8036 30434
rect 7644 30370 7700 30380
rect 7196 28924 7476 28980
rect 7980 29426 8036 30382
rect 7980 29374 7982 29426
rect 8034 29374 8036 29426
rect 6972 28590 6974 28642
rect 7026 28590 7028 28642
rect 6972 28578 7028 28590
rect 7084 28756 7140 28766
rect 7084 28530 7140 28700
rect 7084 28478 7086 28530
rect 7138 28478 7140 28530
rect 7084 28466 7140 28478
rect 6972 28420 7028 28430
rect 6972 28326 7028 28364
rect 6748 27972 6804 27982
rect 6748 27878 6804 27916
rect 6524 27186 6692 27188
rect 6524 27134 6526 27186
rect 6578 27134 6692 27186
rect 6524 27132 6692 27134
rect 6860 27858 6916 27870
rect 6860 27806 6862 27858
rect 6914 27806 6916 27858
rect 6860 27188 6916 27806
rect 6524 27122 6580 27132
rect 6860 27122 6916 27132
rect 5516 26898 5572 26908
rect 5628 26852 5796 26908
rect 5852 27074 5908 27086
rect 5852 27022 5854 27074
rect 5906 27022 5908 27074
rect 5628 26516 5684 26852
rect 5516 26460 5684 26516
rect 5068 25284 5124 25294
rect 5068 25190 5124 25228
rect 5516 25284 5572 26460
rect 5852 26292 5908 27022
rect 6972 27076 7028 27086
rect 5964 26964 6020 26974
rect 6972 26908 7028 27020
rect 5964 26870 6020 26908
rect 6748 26852 7028 26908
rect 5852 26226 5908 26236
rect 6076 26740 6132 26750
rect 6076 26290 6132 26684
rect 6300 26404 6356 26414
rect 6300 26310 6356 26348
rect 6076 26238 6078 26290
rect 6130 26238 6132 26290
rect 5740 26180 5796 26190
rect 5740 25506 5796 26124
rect 5740 25454 5742 25506
rect 5794 25454 5796 25506
rect 5740 25442 5796 25454
rect 5964 25396 6020 25406
rect 5964 25302 6020 25340
rect 5516 25218 5572 25228
rect 6076 25172 6132 26238
rect 6412 26290 6468 26302
rect 6412 26238 6414 26290
rect 6466 26238 6468 26290
rect 5740 25116 6132 25172
rect 6300 25506 6356 25518
rect 6300 25454 6302 25506
rect 6354 25454 6356 25506
rect 5404 25060 5460 25070
rect 5068 24948 5124 24958
rect 5068 24724 5124 24892
rect 5068 24722 5236 24724
rect 5068 24670 5070 24722
rect 5122 24670 5236 24722
rect 5068 24668 5236 24670
rect 5068 24658 5124 24668
rect 4956 23998 4958 24050
rect 5010 23998 5012 24050
rect 4956 23986 5012 23998
rect 5068 24052 5124 24062
rect 4284 23886 4286 23938
rect 4338 23886 4340 23938
rect 4284 23828 4340 23886
rect 4508 23940 4564 23950
rect 4508 23846 4564 23884
rect 4284 23762 4340 23772
rect 4844 23716 4900 23726
rect 5068 23716 5124 23996
rect 4844 23622 4900 23660
rect 4956 23714 5124 23716
rect 4956 23662 5070 23714
rect 5122 23662 5124 23714
rect 4956 23660 5124 23662
rect 4732 23380 4788 23390
rect 4732 23042 4788 23324
rect 4732 22990 4734 23042
rect 4786 22990 4788 23042
rect 4732 22978 4788 22990
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4508 22372 4564 22382
rect 4844 22372 4900 22382
rect 4956 22372 5012 23660
rect 5068 23650 5124 23660
rect 4172 22370 4676 22372
rect 4172 22318 4510 22370
rect 4562 22318 4676 22370
rect 4172 22316 4676 22318
rect 4508 22306 4564 22316
rect 3948 22204 4116 22260
rect 3836 22148 3892 22158
rect 3836 22054 3892 22092
rect 3836 19908 3892 19918
rect 3724 19852 3836 19908
rect 3836 19814 3892 19852
rect 2828 18116 2884 18126
rect 2716 17108 2772 17118
rect 2604 17106 2772 17108
rect 2604 17054 2718 17106
rect 2770 17054 2772 17106
rect 2604 17052 2772 17054
rect 2716 17042 2772 17052
rect 2604 16884 2660 16894
rect 2604 16790 2660 16828
rect 2828 16882 2884 18060
rect 2940 17892 2996 19292
rect 2940 17826 2996 17836
rect 3052 19796 3108 19806
rect 2828 16830 2830 16882
rect 2882 16830 2884 16882
rect 2828 16818 2884 16830
rect 3052 15988 3108 19740
rect 3948 19460 4004 22204
rect 4396 21700 4452 21710
rect 4284 21644 4396 21700
rect 3948 19394 4004 19404
rect 4060 21474 4116 21486
rect 4060 21422 4062 21474
rect 4114 21422 4116 21474
rect 4060 19348 4116 21422
rect 4060 19282 4116 19292
rect 4284 19348 4340 21644
rect 4396 21634 4452 21644
rect 4620 21588 4676 22316
rect 4844 22370 5012 22372
rect 4844 22318 4846 22370
rect 4898 22318 5012 22370
rect 4844 22316 5012 22318
rect 4844 22306 4900 22316
rect 4620 21522 4676 21532
rect 4732 21700 4788 21710
rect 4732 21586 4788 21644
rect 4732 21534 4734 21586
rect 4786 21534 4788 21586
rect 4732 21522 4788 21534
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4844 20914 4900 20926
rect 4844 20862 4846 20914
rect 4898 20862 4900 20914
rect 4396 20018 4452 20030
rect 4396 19966 4398 20018
rect 4450 19966 4452 20018
rect 4396 19796 4452 19966
rect 4844 19796 4900 20862
rect 4396 19740 4900 19796
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4284 19292 4564 19348
rect 3836 19122 3892 19134
rect 3836 19070 3838 19122
rect 3890 19070 3892 19122
rect 3164 18338 3220 18350
rect 3164 18286 3166 18338
rect 3218 18286 3220 18338
rect 3164 17220 3220 18286
rect 3836 18340 3892 19070
rect 4284 18452 4340 19292
rect 4508 19234 4564 19292
rect 4508 19182 4510 19234
rect 4562 19182 4564 19234
rect 4508 19170 4564 19182
rect 4284 18386 4340 18396
rect 3836 18274 3892 18284
rect 3500 18116 3556 18126
rect 4844 18116 4900 19740
rect 4956 18340 5012 22316
rect 5180 21700 5236 24668
rect 5180 21634 5236 21644
rect 5292 21588 5348 21598
rect 5292 21494 5348 21532
rect 5292 20244 5348 20254
rect 5292 19906 5348 20188
rect 5292 19854 5294 19906
rect 5346 19854 5348 19906
rect 5292 19796 5348 19854
rect 5292 19730 5348 19740
rect 5180 19348 5236 19358
rect 5404 19348 5460 25004
rect 5628 24948 5684 24958
rect 5628 24854 5684 24892
rect 5516 23828 5572 23838
rect 5628 23828 5684 23838
rect 5572 23826 5684 23828
rect 5572 23774 5630 23826
rect 5682 23774 5684 23826
rect 5572 23772 5684 23774
rect 5516 21586 5572 23772
rect 5628 23762 5684 23772
rect 5628 23380 5684 23390
rect 5628 22370 5684 23324
rect 5628 22318 5630 22370
rect 5682 22318 5684 22370
rect 5628 22306 5684 22318
rect 5516 21534 5518 21586
rect 5570 21534 5572 21586
rect 5516 21522 5572 21534
rect 5740 21364 5796 25116
rect 6188 24836 6244 24846
rect 6300 24836 6356 25454
rect 6412 24948 6468 26238
rect 6748 25732 6804 26852
rect 7196 26516 7252 28924
rect 7196 26450 7252 26460
rect 7308 28756 7364 28766
rect 7308 26404 7364 28700
rect 7980 28196 8036 29374
rect 8092 28756 8148 31948
rect 8316 31890 8372 31948
rect 8540 32002 8596 32060
rect 8540 31950 8542 32002
rect 8594 31950 8596 32002
rect 8540 31938 8596 31950
rect 8316 31838 8318 31890
rect 8370 31838 8372 31890
rect 8316 31826 8372 31838
rect 8204 31780 8260 31790
rect 8204 31106 8260 31724
rect 8652 31220 8708 35868
rect 8876 35698 8932 35710
rect 8876 35646 8878 35698
rect 8930 35646 8932 35698
rect 8876 34916 8932 35646
rect 9324 34916 9380 36876
rect 9660 36820 9716 37548
rect 9436 36764 9716 36820
rect 9772 37492 9828 37502
rect 9772 37266 9828 37436
rect 9772 37214 9774 37266
rect 9826 37214 9828 37266
rect 9436 36482 9492 36764
rect 9436 36430 9438 36482
rect 9490 36430 9492 36482
rect 9436 36418 9492 36430
rect 9548 36372 9604 36382
rect 9548 36370 9716 36372
rect 9548 36318 9550 36370
rect 9602 36318 9716 36370
rect 9548 36316 9716 36318
rect 9548 36306 9604 36316
rect 9660 35700 9716 36316
rect 9772 35924 9828 37214
rect 9884 36708 9940 38612
rect 9996 36708 10052 36718
rect 9884 36706 10052 36708
rect 9884 36654 9998 36706
rect 10050 36654 10052 36706
rect 9884 36652 10052 36654
rect 9996 36642 10052 36652
rect 10108 35924 10164 38780
rect 10220 37492 10276 39116
rect 10556 38946 10612 38958
rect 10556 38894 10558 38946
rect 10610 38894 10612 38946
rect 10332 38834 10388 38846
rect 10332 38782 10334 38834
rect 10386 38782 10388 38834
rect 10332 38050 10388 38782
rect 10556 38724 10612 38894
rect 10668 38834 10724 39116
rect 10668 38782 10670 38834
rect 10722 38782 10724 38834
rect 10668 38770 10724 38782
rect 10556 38658 10612 38668
rect 10332 37998 10334 38050
rect 10386 37998 10388 38050
rect 10332 37986 10388 37998
rect 10780 38612 10836 39676
rect 11116 39618 11172 40124
rect 11564 39844 11620 40348
rect 11788 40404 11844 40414
rect 11788 40310 11844 40348
rect 11900 40292 11956 40302
rect 11788 39844 11844 39854
rect 11564 39842 11844 39844
rect 11564 39790 11790 39842
rect 11842 39790 11844 39842
rect 11564 39788 11844 39790
rect 11788 39778 11844 39788
rect 11676 39620 11732 39630
rect 11116 39566 11118 39618
rect 11170 39566 11172 39618
rect 11116 39554 11172 39566
rect 11228 39618 11732 39620
rect 11228 39566 11678 39618
rect 11730 39566 11732 39618
rect 11228 39564 11732 39566
rect 11004 39508 11060 39518
rect 10892 39394 10948 39406
rect 10892 39342 10894 39394
rect 10946 39342 10948 39394
rect 10892 39284 10948 39342
rect 10892 39218 10948 39228
rect 11004 38948 11060 39452
rect 11228 39506 11284 39564
rect 11228 39454 11230 39506
rect 11282 39454 11284 39506
rect 11228 39442 11284 39454
rect 11116 39060 11172 39070
rect 11116 38966 11172 39004
rect 11340 39058 11396 39564
rect 11676 39554 11732 39564
rect 11788 39508 11844 39518
rect 11900 39508 11956 40236
rect 11788 39506 11956 39508
rect 11788 39454 11790 39506
rect 11842 39454 11956 39506
rect 11788 39452 11956 39454
rect 11340 39006 11342 39058
rect 11394 39006 11396 39058
rect 11340 38994 11396 39006
rect 11452 39394 11508 39406
rect 11452 39342 11454 39394
rect 11506 39342 11508 39394
rect 11004 38854 11060 38892
rect 11228 38948 11284 38958
rect 10444 37940 10500 37950
rect 10444 37846 10500 37884
rect 10668 37828 10724 37838
rect 10220 37426 10276 37436
rect 10556 37826 10724 37828
rect 10556 37774 10670 37826
rect 10722 37774 10724 37826
rect 10556 37772 10724 37774
rect 10220 37268 10276 37278
rect 10444 37268 10500 37278
rect 10220 37266 10444 37268
rect 10220 37214 10222 37266
rect 10274 37214 10444 37266
rect 10220 37212 10444 37214
rect 10220 37202 10276 37212
rect 10444 37202 10500 37212
rect 10444 37044 10500 37054
rect 10332 36820 10388 36830
rect 10332 36484 10388 36764
rect 10444 36706 10500 36988
rect 10444 36654 10446 36706
rect 10498 36654 10500 36706
rect 10444 36642 10500 36654
rect 10332 36428 10500 36484
rect 10220 35924 10276 35934
rect 10108 35922 10276 35924
rect 10108 35870 10222 35922
rect 10274 35870 10276 35922
rect 10108 35868 10276 35870
rect 9772 35830 9828 35868
rect 10220 35858 10276 35868
rect 9996 35812 10052 35822
rect 9884 35700 9940 35710
rect 9660 35698 9940 35700
rect 9660 35646 9886 35698
rect 9938 35646 9940 35698
rect 9660 35644 9940 35646
rect 9884 35634 9940 35644
rect 9884 35028 9940 35038
rect 9660 34916 9716 34926
rect 8876 34914 9716 34916
rect 8876 34862 9662 34914
rect 9714 34862 9716 34914
rect 8876 34860 9716 34862
rect 8764 34802 8820 34814
rect 8764 34750 8766 34802
rect 8818 34750 8820 34802
rect 8764 33124 8820 34750
rect 8876 34692 8932 34702
rect 9100 34692 9156 34702
rect 8876 34690 9044 34692
rect 8876 34638 8878 34690
rect 8930 34638 9044 34690
rect 8876 34636 9044 34638
rect 8876 34626 8932 34636
rect 8876 34130 8932 34142
rect 8876 34078 8878 34130
rect 8930 34078 8932 34130
rect 8876 33572 8932 34078
rect 8876 33506 8932 33516
rect 8988 33348 9044 34636
rect 9100 34598 9156 34636
rect 8988 33282 9044 33292
rect 9436 34580 9492 34590
rect 8764 32396 8820 33068
rect 8988 32562 9044 32574
rect 8988 32510 8990 32562
rect 9042 32510 9044 32562
rect 8764 32340 8932 32396
rect 8764 32004 8820 32014
rect 8764 31444 8820 31948
rect 8876 32002 8932 32340
rect 8876 31950 8878 32002
rect 8930 31950 8932 32002
rect 8876 31668 8932 31950
rect 8876 31602 8932 31612
rect 8988 31892 9044 32510
rect 9436 32004 9492 34524
rect 9660 32116 9716 34860
rect 9772 34804 9828 34814
rect 9884 34804 9940 34972
rect 9996 34916 10052 35756
rect 9996 34850 10052 34860
rect 10444 35364 10500 36428
rect 10556 36482 10612 37772
rect 10668 37762 10724 37772
rect 10668 37380 10724 37390
rect 10668 37286 10724 37324
rect 10556 36430 10558 36482
rect 10610 36430 10612 36482
rect 10556 36418 10612 36430
rect 10780 37268 10836 38556
rect 11228 38050 11284 38892
rect 11452 38836 11508 39342
rect 11788 39396 11844 39452
rect 11788 39330 11844 39340
rect 11452 38770 11508 38780
rect 11564 39060 11620 39070
rect 11564 38724 11620 39004
rect 11228 37998 11230 38050
rect 11282 37998 11284 38050
rect 11228 37986 11284 37998
rect 11340 38612 11620 38668
rect 12012 38722 12068 38734
rect 12012 38670 12014 38722
rect 12066 38670 12068 38722
rect 10892 37938 10948 37950
rect 10892 37886 10894 37938
rect 10946 37886 10948 37938
rect 10892 37492 10948 37886
rect 11004 37828 11060 37838
rect 11004 37734 11060 37772
rect 10892 37436 11172 37492
rect 11004 37268 11060 37278
rect 10780 37266 11060 37268
rect 10780 37214 11006 37266
rect 11058 37214 11060 37266
rect 10780 37212 11060 37214
rect 10668 35924 10724 35934
rect 10668 35698 10724 35868
rect 10668 35646 10670 35698
rect 10722 35646 10724 35698
rect 10668 35634 10724 35646
rect 9828 34748 9940 34804
rect 10332 34804 10388 34814
rect 9772 34738 9828 34748
rect 10332 34710 10388 34748
rect 9996 34242 10052 34254
rect 9996 34190 9998 34242
rect 10050 34190 10052 34242
rect 9772 34020 9828 34030
rect 9772 33908 9828 33964
rect 9772 33906 9940 33908
rect 9772 33854 9774 33906
rect 9826 33854 9940 33906
rect 9772 33852 9940 33854
rect 9772 33842 9828 33852
rect 9884 32452 9940 33852
rect 9996 33460 10052 34190
rect 10332 34132 10388 34142
rect 10332 34038 10388 34076
rect 10108 34020 10164 34030
rect 10108 33926 10164 33964
rect 10332 33796 10388 33806
rect 9996 33124 10052 33404
rect 10108 33740 10332 33796
rect 10108 33458 10164 33740
rect 10332 33730 10388 33740
rect 10108 33406 10110 33458
rect 10162 33406 10164 33458
rect 10108 33394 10164 33406
rect 9996 33068 10164 33124
rect 10108 32674 10164 33068
rect 10108 32622 10110 32674
rect 10162 32622 10164 32674
rect 10108 32610 10164 32622
rect 9996 32452 10052 32462
rect 9884 32450 10164 32452
rect 9884 32398 9998 32450
rect 10050 32398 10164 32450
rect 9884 32396 10164 32398
rect 9996 32386 10052 32396
rect 9772 32116 9828 32126
rect 9660 32060 9772 32116
rect 9772 32050 9828 32060
rect 9436 31938 9492 31948
rect 8764 31388 8932 31444
rect 8764 31220 8820 31230
rect 8652 31218 8820 31220
rect 8652 31166 8766 31218
rect 8818 31166 8820 31218
rect 8652 31164 8820 31166
rect 8764 31154 8820 31164
rect 8204 31054 8206 31106
rect 8258 31054 8260 31106
rect 8204 30996 8260 31054
rect 8876 30996 8932 31388
rect 8988 31108 9044 31836
rect 9772 31890 9828 31902
rect 9772 31838 9774 31890
rect 9826 31838 9828 31890
rect 9436 31780 9492 31790
rect 9436 31686 9492 31724
rect 9212 31668 9268 31678
rect 8988 31042 9044 31052
rect 9100 31666 9268 31668
rect 9100 31614 9214 31666
rect 9266 31614 9268 31666
rect 9100 31612 9268 31614
rect 8204 30930 8260 30940
rect 8652 30940 8932 30996
rect 8428 30772 8484 30782
rect 8428 30678 8484 30716
rect 8652 30210 8708 30940
rect 8652 30158 8654 30210
rect 8706 30158 8708 30210
rect 8652 30146 8708 30158
rect 8764 30100 8820 30110
rect 9100 30100 9156 31612
rect 9212 31602 9268 31612
rect 9660 31108 9716 31118
rect 9660 30994 9716 31052
rect 9660 30942 9662 30994
rect 9714 30942 9716 30994
rect 9660 30930 9716 30942
rect 9436 30772 9492 30782
rect 9212 30212 9268 30222
rect 9212 30118 9268 30156
rect 8764 30098 9156 30100
rect 8764 30046 8766 30098
rect 8818 30046 9156 30098
rect 8764 30044 9156 30046
rect 8428 29540 8484 29550
rect 8428 29446 8484 29484
rect 8540 29316 8596 29326
rect 8596 29260 8708 29316
rect 8540 29250 8596 29260
rect 8540 28868 8596 28878
rect 8092 28690 8148 28700
rect 8428 28754 8484 28766
rect 8428 28702 8430 28754
rect 8482 28702 8484 28754
rect 7980 28130 8036 28140
rect 8316 28084 8372 28094
rect 7644 27972 7700 27982
rect 7532 27860 7588 27898
rect 7532 27794 7588 27804
rect 7420 27748 7476 27758
rect 7420 27654 7476 27692
rect 7532 27636 7588 27646
rect 7532 27074 7588 27580
rect 7532 27022 7534 27074
rect 7586 27022 7588 27074
rect 7532 27010 7588 27022
rect 7308 26338 7364 26348
rect 7644 26962 7700 27916
rect 8316 27186 8372 28028
rect 8316 27134 8318 27186
rect 8370 27134 8372 27186
rect 8316 27122 8372 27134
rect 8428 27076 8484 28702
rect 8540 28642 8596 28812
rect 8540 28590 8542 28642
rect 8594 28590 8596 28642
rect 8540 28578 8596 28590
rect 8428 27010 8484 27020
rect 8540 28420 8596 28430
rect 8540 27858 8596 28364
rect 8652 27972 8708 29260
rect 8652 27878 8708 27916
rect 8540 27806 8542 27858
rect 8594 27806 8596 27858
rect 7644 26910 7646 26962
rect 7698 26910 7700 26962
rect 7084 26068 7140 26078
rect 6412 24882 6468 24892
rect 6524 25676 6804 25732
rect 6972 26012 7084 26068
rect 6972 25730 7028 26012
rect 7084 26002 7140 26012
rect 6972 25678 6974 25730
rect 7026 25678 7028 25730
rect 6524 24946 6580 25676
rect 6972 25666 7028 25678
rect 6636 25508 6692 25518
rect 6748 25508 6804 25518
rect 6636 25506 6748 25508
rect 6636 25454 6638 25506
rect 6690 25454 6748 25506
rect 6636 25452 6748 25454
rect 6636 25442 6692 25452
rect 6524 24894 6526 24946
rect 6578 24894 6580 24946
rect 6524 24882 6580 24894
rect 6244 24780 6356 24836
rect 6188 24162 6244 24780
rect 6524 24724 6580 24734
rect 6748 24724 6804 25452
rect 7420 25284 7476 25294
rect 6972 24836 7028 24846
rect 6972 24742 7028 24780
rect 6524 24722 6804 24724
rect 6524 24670 6526 24722
rect 6578 24670 6804 24722
rect 6524 24668 6804 24670
rect 6524 24658 6580 24668
rect 6188 24110 6190 24162
rect 6242 24110 6244 24162
rect 6188 24098 6244 24110
rect 6076 23940 6132 23950
rect 6076 22482 6132 23884
rect 6412 23492 6468 23502
rect 6300 23436 6412 23492
rect 6188 23156 6244 23166
rect 6188 23062 6244 23100
rect 6076 22430 6078 22482
rect 6130 22430 6132 22482
rect 6076 22418 6132 22430
rect 5852 21700 5908 21710
rect 5908 21644 6020 21700
rect 5852 21634 5908 21644
rect 5852 21364 5908 21374
rect 5796 21362 5908 21364
rect 5796 21310 5854 21362
rect 5906 21310 5908 21362
rect 5796 21308 5908 21310
rect 5740 20916 5796 21308
rect 5852 21298 5908 21308
rect 5964 21140 6020 21644
rect 5740 20850 5796 20860
rect 5852 21084 6020 21140
rect 5740 20018 5796 20030
rect 5740 19966 5742 20018
rect 5794 19966 5796 20018
rect 5180 19346 5460 19348
rect 5180 19294 5182 19346
rect 5234 19294 5460 19346
rect 5180 19292 5460 19294
rect 5628 19348 5684 19358
rect 5180 19282 5236 19292
rect 5628 19254 5684 19292
rect 5516 18452 5572 18462
rect 4956 18284 5124 18340
rect 4956 18116 5012 18126
rect 3500 17780 3556 18060
rect 4476 18060 4740 18070
rect 4844 18060 4956 18116
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4956 18050 5012 18060
rect 4476 17994 4740 18004
rect 4396 17892 4452 17902
rect 3500 17724 3780 17780
rect 3724 17666 3780 17724
rect 3724 17614 3726 17666
rect 3778 17614 3780 17666
rect 3724 17602 3780 17614
rect 3948 17668 4004 17678
rect 3948 17554 4004 17612
rect 3948 17502 3950 17554
rect 4002 17502 4004 17554
rect 3948 17490 4004 17502
rect 3276 17444 3332 17454
rect 3276 17350 3332 17388
rect 3500 17442 3556 17454
rect 3500 17390 3502 17442
rect 3554 17390 3556 17442
rect 3164 17164 3332 17220
rect 3164 16996 3220 17006
rect 3164 16902 3220 16940
rect 3164 16772 3220 16782
rect 3164 16210 3220 16716
rect 3164 16158 3166 16210
rect 3218 16158 3220 16210
rect 3164 16146 3220 16158
rect 3276 16212 3332 17164
rect 3500 16884 3556 17390
rect 3612 17442 3668 17454
rect 3612 17390 3614 17442
rect 3666 17390 3668 17442
rect 3612 16996 3668 17390
rect 3724 17220 3780 17230
rect 3724 17106 3780 17164
rect 3724 17054 3726 17106
rect 3778 17054 3780 17106
rect 4396 17108 4452 17836
rect 4844 17892 4900 17902
rect 5068 17892 5124 18284
rect 4620 17778 4676 17790
rect 4620 17726 4622 17778
rect 4674 17726 4676 17778
rect 4620 17444 4676 17726
rect 4844 17668 4900 17836
rect 4844 17602 4900 17612
rect 4956 17836 5124 17892
rect 5180 18004 5236 18014
rect 4956 17444 5012 17836
rect 5068 17668 5124 17678
rect 5180 17668 5236 17948
rect 5068 17666 5236 17668
rect 5068 17614 5070 17666
rect 5122 17614 5236 17666
rect 5068 17612 5236 17614
rect 5516 17668 5572 18396
rect 5740 18228 5796 19966
rect 5740 18162 5796 18172
rect 5852 18674 5908 21084
rect 6300 21026 6356 23436
rect 6412 23426 6468 23436
rect 6300 20974 6302 21026
rect 6354 20974 6356 21026
rect 6300 20962 6356 20974
rect 6748 21028 6804 24668
rect 7420 23266 7476 25228
rect 7420 23214 7422 23266
rect 7474 23214 7476 23266
rect 6748 20962 6804 20972
rect 6972 22484 7028 22494
rect 6972 21698 7028 22428
rect 6972 21646 6974 21698
rect 7026 21646 7028 21698
rect 6076 20802 6132 20814
rect 6076 20750 6078 20802
rect 6130 20750 6132 20802
rect 6076 20692 6132 20750
rect 6300 20804 6356 20814
rect 6748 20804 6804 20814
rect 6356 20802 6804 20804
rect 6356 20750 6750 20802
rect 6802 20750 6804 20802
rect 6356 20748 6804 20750
rect 6300 20710 6356 20748
rect 6748 20738 6804 20748
rect 6076 20626 6132 20636
rect 6524 20580 6580 20590
rect 6188 19460 6244 19470
rect 5964 19122 6020 19134
rect 5964 19070 5966 19122
rect 6018 19070 6020 19122
rect 5964 18900 6020 19070
rect 6076 19124 6132 19134
rect 6076 19030 6132 19068
rect 6188 19122 6244 19404
rect 6188 19070 6190 19122
rect 6242 19070 6244 19122
rect 6188 19012 6244 19070
rect 6188 18946 6244 18956
rect 6412 19010 6468 19022
rect 6412 18958 6414 19010
rect 6466 18958 6468 19010
rect 5964 18834 6020 18844
rect 6412 18676 6468 18958
rect 5852 18622 5854 18674
rect 5906 18622 5908 18674
rect 5852 18004 5908 18622
rect 5852 17938 5908 17948
rect 6188 18620 6412 18676
rect 6188 17668 6244 18620
rect 6412 18582 6468 18620
rect 6524 18674 6580 20524
rect 6860 20132 6916 20142
rect 6972 20132 7028 21646
rect 7420 21812 7476 23214
rect 7420 20244 7476 21756
rect 7420 20178 7476 20188
rect 6860 20130 7028 20132
rect 6860 20078 6862 20130
rect 6914 20078 7028 20130
rect 6860 20076 7028 20078
rect 6860 20066 6916 20076
rect 7644 19684 7700 26910
rect 7756 26964 7812 26974
rect 8540 26908 8596 27806
rect 8764 26908 8820 30044
rect 8876 29876 8932 29886
rect 8876 29426 8932 29820
rect 8876 29374 8878 29426
rect 8930 29374 8932 29426
rect 8876 29362 8932 29374
rect 8988 29428 9044 29438
rect 8988 28644 9044 29372
rect 9436 28866 9492 30716
rect 9548 30436 9604 30446
rect 9548 29986 9604 30380
rect 9660 30212 9716 30222
rect 9660 30118 9716 30156
rect 9548 29934 9550 29986
rect 9602 29934 9604 29986
rect 9548 29922 9604 29934
rect 9772 29876 9828 31838
rect 9884 31556 9940 31566
rect 9884 30210 9940 31500
rect 9884 30158 9886 30210
rect 9938 30158 9940 30210
rect 9884 30146 9940 30158
rect 9772 29810 9828 29820
rect 9884 29540 9940 29550
rect 9884 29446 9940 29484
rect 9548 29428 9604 29438
rect 9548 29334 9604 29372
rect 9436 28814 9438 28866
rect 9490 28814 9492 28866
rect 9436 28802 9492 28814
rect 8988 28578 9044 28588
rect 9212 28756 9268 28766
rect 9212 28642 9268 28700
rect 9212 28590 9214 28642
rect 9266 28590 9268 28642
rect 9212 28578 9268 28590
rect 10108 28754 10164 32396
rect 10220 31890 10276 31902
rect 10220 31838 10222 31890
rect 10274 31838 10276 31890
rect 10220 31220 10276 31838
rect 10332 31778 10388 31790
rect 10332 31726 10334 31778
rect 10386 31726 10388 31778
rect 10332 31332 10388 31726
rect 10332 31266 10388 31276
rect 10220 31154 10276 31164
rect 10332 30882 10388 30894
rect 10332 30830 10334 30882
rect 10386 30830 10388 30882
rect 10332 30436 10388 30830
rect 10332 30370 10388 30380
rect 10332 30210 10388 30222
rect 10332 30158 10334 30210
rect 10386 30158 10388 30210
rect 10220 30098 10276 30110
rect 10220 30046 10222 30098
rect 10274 30046 10276 30098
rect 10220 29764 10276 30046
rect 10220 29698 10276 29708
rect 10108 28702 10110 28754
rect 10162 28702 10164 28754
rect 9884 28532 9940 28542
rect 9212 28196 9268 28206
rect 7756 25506 7812 26908
rect 8428 26852 8596 26908
rect 8652 26852 8820 26908
rect 8876 27858 8932 27870
rect 8876 27806 8878 27858
rect 8930 27806 8932 27858
rect 8876 26908 8932 27806
rect 8876 26852 9044 26908
rect 8204 26290 8260 26302
rect 8204 26238 8206 26290
rect 8258 26238 8260 26290
rect 8204 26068 8260 26238
rect 8204 26002 8260 26012
rect 7756 25454 7758 25506
rect 7810 25454 7812 25506
rect 7756 23938 7812 25454
rect 8204 24724 8260 24734
rect 8204 24630 8260 24668
rect 7756 23886 7758 23938
rect 7810 23886 7812 23938
rect 7756 23874 7812 23886
rect 8092 24050 8148 24062
rect 8092 23998 8094 24050
rect 8146 23998 8148 24050
rect 7980 23154 8036 23166
rect 7980 23102 7982 23154
rect 8034 23102 8036 23154
rect 7756 22482 7812 22494
rect 7756 22430 7758 22482
rect 7810 22430 7812 22482
rect 7756 21028 7812 22430
rect 7756 20962 7812 20972
rect 7868 21586 7924 21598
rect 7868 21534 7870 21586
rect 7922 21534 7924 21586
rect 7756 20802 7812 20814
rect 7756 20750 7758 20802
rect 7810 20750 7812 20802
rect 7756 20692 7812 20750
rect 7756 20242 7812 20636
rect 7756 20190 7758 20242
rect 7810 20190 7812 20242
rect 7756 20178 7812 20190
rect 7868 20018 7924 21534
rect 7980 20468 8036 23102
rect 8092 20580 8148 23998
rect 8316 24052 8372 24062
rect 8316 23378 8372 23996
rect 8316 23326 8318 23378
rect 8370 23326 8372 23378
rect 8316 23314 8372 23326
rect 8204 23042 8260 23054
rect 8204 22990 8206 23042
rect 8258 22990 8260 23042
rect 8204 22932 8260 22990
rect 8204 22866 8260 22876
rect 8428 22820 8484 26852
rect 8652 25618 8708 26852
rect 8652 25566 8654 25618
rect 8706 25566 8708 25618
rect 8540 25508 8596 25518
rect 8540 25414 8596 25452
rect 8316 22764 8484 22820
rect 8316 21810 8372 22764
rect 8316 21758 8318 21810
rect 8370 21758 8372 21810
rect 8316 21746 8372 21758
rect 8204 21700 8260 21710
rect 8204 21586 8260 21644
rect 8204 21534 8206 21586
rect 8258 21534 8260 21586
rect 8204 21522 8260 21534
rect 8092 20514 8148 20524
rect 8540 21028 8596 21038
rect 7980 20402 8036 20412
rect 7868 19966 7870 20018
rect 7922 19966 7924 20018
rect 7644 19628 7812 19684
rect 7644 19460 7700 19470
rect 7084 19236 7140 19246
rect 6524 18622 6526 18674
rect 6578 18622 6580 18674
rect 6524 18610 6580 18622
rect 6972 19234 7140 19236
rect 6972 19182 7086 19234
rect 7138 19182 7140 19234
rect 6972 19180 7140 19182
rect 6300 18452 6356 18462
rect 6300 17778 6356 18396
rect 6300 17726 6302 17778
rect 6354 17726 6356 17778
rect 6300 17714 6356 17726
rect 6524 18450 6580 18462
rect 6524 18398 6526 18450
rect 6578 18398 6580 18450
rect 6524 18116 6580 18398
rect 5068 17602 5124 17612
rect 5404 17556 5460 17566
rect 5180 17500 5404 17556
rect 4620 17388 5124 17444
rect 4508 17108 4564 17118
rect 4396 17106 4564 17108
rect 3724 17042 3780 17054
rect 4060 17050 4116 17062
rect 4396 17054 4510 17106
rect 4562 17054 4564 17106
rect 4396 17052 4564 17054
rect 4060 16998 4062 17050
rect 4114 16998 4116 17050
rect 4508 17042 4564 17052
rect 4060 16996 4116 16998
rect 3612 16930 3668 16940
rect 3836 16940 4116 16996
rect 3276 16146 3332 16156
rect 3388 16828 3500 16884
rect 3052 15932 3332 15988
rect 2716 15876 2772 15886
rect 2380 15820 2548 15876
rect 2156 15486 2158 15538
rect 2210 15486 2212 15538
rect 2156 15316 2212 15486
rect 2492 15540 2548 15820
rect 2716 15782 2772 15820
rect 2492 15484 2772 15540
rect 2604 15316 2660 15326
rect 2156 15314 2660 15316
rect 2156 15262 2606 15314
rect 2658 15262 2660 15314
rect 2156 15260 2660 15262
rect 2380 14754 2436 14766
rect 2380 14702 2382 14754
rect 2434 14702 2436 14754
rect 2380 14642 2436 14702
rect 2380 14590 2382 14642
rect 2434 14590 2436 14642
rect 1820 14306 1876 14318
rect 1820 14254 1822 14306
rect 1874 14254 1876 14306
rect 1820 13188 1876 14254
rect 2268 13972 2324 13982
rect 2268 13878 2324 13916
rect 2044 13188 2100 13198
rect 1820 13186 2100 13188
rect 1820 13134 2046 13186
rect 2098 13134 2100 13186
rect 1820 13132 2100 13134
rect 1932 12740 1988 12750
rect 2044 12740 2100 13132
rect 2380 13074 2436 14590
rect 2492 13186 2548 15260
rect 2604 15250 2660 15260
rect 2716 14754 2772 15484
rect 3164 15202 3220 15214
rect 3164 15150 3166 15202
rect 3218 15150 3220 15202
rect 2716 14702 2718 14754
rect 2770 14702 2772 14754
rect 2716 14690 2772 14702
rect 2828 15092 2884 15102
rect 2828 14642 2884 15036
rect 2828 14590 2830 14642
rect 2882 14590 2884 14642
rect 2828 14578 2884 14590
rect 2716 14420 2772 14430
rect 2716 13970 2772 14364
rect 2716 13918 2718 13970
rect 2770 13918 2772 13970
rect 2716 13906 2772 13918
rect 3164 13748 3220 15150
rect 3276 14642 3332 15932
rect 3276 14590 3278 14642
rect 3330 14590 3332 14642
rect 3276 14578 3332 14590
rect 3164 13682 3220 13692
rect 2492 13134 2494 13186
rect 2546 13134 2548 13186
rect 2492 13122 2548 13134
rect 3052 13634 3108 13646
rect 3052 13582 3054 13634
rect 3106 13582 3108 13634
rect 3052 13186 3108 13582
rect 3052 13134 3054 13186
rect 3106 13134 3108 13186
rect 3052 13122 3108 13134
rect 3276 13188 3332 13198
rect 2380 13022 2382 13074
rect 2434 13022 2436 13074
rect 2380 13010 2436 13022
rect 2828 12740 2884 12750
rect 3276 12740 3332 13132
rect 1932 12738 2100 12740
rect 1932 12686 1934 12738
rect 1986 12686 2100 12738
rect 1932 12684 2100 12686
rect 1932 12674 1988 12684
rect 1932 12516 1988 12526
rect 1932 12402 1988 12460
rect 1932 12350 1934 12402
rect 1986 12350 1988 12402
rect 1932 12338 1988 12350
rect 2044 12068 2100 12684
rect 2716 12738 3332 12740
rect 2716 12686 2830 12738
rect 2882 12686 3278 12738
rect 3330 12686 3332 12738
rect 2716 12684 3332 12686
rect 2268 12068 2324 12078
rect 2044 12066 2324 12068
rect 2044 12014 2270 12066
rect 2322 12014 2324 12066
rect 2044 12012 2324 12014
rect 1820 11508 1876 11518
rect 2156 11508 2212 12012
rect 2268 12002 2324 12012
rect 1820 11506 2212 11508
rect 1820 11454 1822 11506
rect 1874 11454 2212 11506
rect 1820 11452 2212 11454
rect 2268 11844 2324 11854
rect 1820 11442 1876 11452
rect 2268 11394 2324 11788
rect 2268 11342 2270 11394
rect 2322 11342 2324 11394
rect 2156 10500 2212 10510
rect 2268 10500 2324 11342
rect 2492 10500 2548 10510
rect 2268 10498 2548 10500
rect 2268 10446 2494 10498
rect 2546 10446 2548 10498
rect 2268 10444 2548 10446
rect 2156 10406 2212 10444
rect 2044 9716 2100 9726
rect 2044 9622 2100 9660
rect 2380 9604 2436 9614
rect 2492 9604 2548 10444
rect 2380 9602 2548 9604
rect 2380 9550 2382 9602
rect 2434 9550 2548 9602
rect 2380 9548 2548 9550
rect 2044 9044 2100 9054
rect 2044 8950 2100 8988
rect 1932 8372 1988 8382
rect 2380 8372 2436 9548
rect 2492 8930 2548 8942
rect 2492 8878 2494 8930
rect 2546 8878 2548 8930
rect 2492 8818 2548 8878
rect 2492 8766 2494 8818
rect 2546 8766 2548 8818
rect 2492 8754 2548 8766
rect 2716 8818 2772 12684
rect 2828 12674 2884 12684
rect 3276 12674 3332 12684
rect 3388 12516 3444 16828
rect 3500 16818 3556 16828
rect 3836 16884 3892 16940
rect 4172 16884 4228 16894
rect 3836 16818 3892 16828
rect 3948 16882 4228 16884
rect 3948 16830 4174 16882
rect 4226 16830 4228 16882
rect 3948 16828 4228 16830
rect 3948 15988 4004 16828
rect 4172 16818 4228 16828
rect 4956 16884 5012 16894
rect 4956 16770 5012 16828
rect 4956 16718 4958 16770
rect 5010 16718 5012 16770
rect 4956 16706 5012 16718
rect 4060 16660 4116 16698
rect 4060 16594 4116 16604
rect 4956 16548 5012 16558
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4844 16492 4956 16548
rect 3948 15922 4004 15932
rect 4060 16324 4116 16334
rect 4060 16210 4116 16268
rect 4396 16324 4452 16334
rect 4844 16324 4900 16492
rect 4956 16482 5012 16492
rect 4396 16322 4900 16324
rect 4396 16270 4398 16322
rect 4450 16270 4900 16322
rect 4396 16268 4900 16270
rect 4396 16258 4452 16268
rect 4060 16158 4062 16210
rect 4114 16158 4116 16210
rect 3500 15874 3556 15886
rect 3500 15822 3502 15874
rect 3554 15822 3556 15874
rect 3500 15652 3556 15822
rect 3500 15538 3556 15596
rect 3500 15486 3502 15538
rect 3554 15486 3556 15538
rect 3500 15474 3556 15486
rect 3948 15540 4004 15550
rect 3948 15314 4004 15484
rect 3948 15262 3950 15314
rect 4002 15262 4004 15314
rect 3948 15250 4004 15262
rect 4060 14532 4116 16158
rect 4396 16100 4452 16110
rect 4284 15988 4340 15998
rect 4284 15894 4340 15932
rect 4396 15986 4452 16044
rect 4396 15934 4398 15986
rect 4450 15934 4452 15986
rect 4396 15922 4452 15934
rect 4844 15988 4900 15998
rect 4844 15894 4900 15932
rect 4956 15876 5012 15886
rect 4956 15782 5012 15820
rect 5068 15652 5124 17388
rect 5180 16098 5236 17500
rect 5404 17490 5460 17500
rect 5516 17108 5572 17612
rect 6076 17612 6244 17668
rect 5964 17444 6020 17454
rect 6076 17444 6132 17612
rect 6300 17556 6356 17566
rect 6300 17462 6356 17500
rect 5964 17442 6132 17444
rect 5964 17390 5966 17442
rect 6018 17390 6132 17442
rect 5964 17388 6132 17390
rect 6188 17442 6244 17454
rect 6188 17390 6190 17442
rect 6242 17390 6244 17442
rect 5516 17106 5908 17108
rect 5516 17054 5518 17106
rect 5570 17054 5908 17106
rect 5516 17052 5908 17054
rect 5516 17042 5572 17052
rect 5180 16046 5182 16098
rect 5234 16046 5236 16098
rect 5180 16034 5236 16046
rect 5740 16884 5796 16894
rect 4956 15596 5124 15652
rect 5628 15988 5684 15998
rect 4620 15540 4676 15550
rect 4172 15426 4228 15438
rect 4172 15374 4174 15426
rect 4226 15374 4228 15426
rect 4172 14756 4228 15374
rect 4620 15314 4676 15484
rect 4620 15262 4622 15314
rect 4674 15262 4676 15314
rect 4620 15250 4676 15262
rect 4844 15426 4900 15438
rect 4844 15374 4846 15426
rect 4898 15374 4900 15426
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4172 14690 4228 14700
rect 4844 14644 4900 15374
rect 4844 14578 4900 14588
rect 4060 14476 4340 14532
rect 3612 14306 3668 14318
rect 3612 14254 3614 14306
rect 3666 14254 3668 14306
rect 3500 13746 3556 13758
rect 3500 13694 3502 13746
rect 3554 13694 3556 13746
rect 3500 13076 3556 13694
rect 3500 13010 3556 13020
rect 3612 13636 3668 14254
rect 3164 12460 3444 12516
rect 3052 12180 3108 12190
rect 2828 12068 2884 12078
rect 2828 11974 2884 12012
rect 3052 11844 3108 12124
rect 3052 11778 3108 11788
rect 2940 11282 2996 11294
rect 2940 11230 2942 11282
rect 2994 11230 2996 11282
rect 2940 10836 2996 11230
rect 2940 10770 2996 10780
rect 3052 10948 3108 10958
rect 3052 10834 3108 10892
rect 3052 10782 3054 10834
rect 3106 10782 3108 10834
rect 3052 10770 3108 10782
rect 2940 10050 2996 10062
rect 2940 9998 2942 10050
rect 2994 9998 2996 10050
rect 2940 9938 2996 9998
rect 2940 9886 2942 9938
rect 2994 9886 2996 9938
rect 2940 9874 2996 9886
rect 2940 9268 2996 9278
rect 2940 9174 2996 9212
rect 2716 8766 2718 8818
rect 2770 8766 2772 8818
rect 2716 8754 2772 8766
rect 3164 8372 3220 12460
rect 3500 11508 3556 11518
rect 3500 10834 3556 11452
rect 3500 10782 3502 10834
rect 3554 10782 3556 10834
rect 3500 10770 3556 10782
rect 3612 10050 3668 13580
rect 4060 14306 4116 14318
rect 4060 14254 4062 14306
rect 4114 14254 4116 14306
rect 4060 13076 4116 14254
rect 4172 14308 4228 14318
rect 4172 13858 4228 14252
rect 4172 13806 4174 13858
rect 4226 13806 4228 13858
rect 4172 13794 4228 13806
rect 3948 13020 4060 13076
rect 3724 12740 3780 12750
rect 3948 12740 4004 13020
rect 4060 13010 4116 13020
rect 4172 12740 4228 12750
rect 3724 12738 4004 12740
rect 3724 12686 3726 12738
rect 3778 12686 4004 12738
rect 3724 12684 4004 12686
rect 3724 12674 3780 12684
rect 3836 12292 3892 12302
rect 3836 12198 3892 12236
rect 3948 12180 4004 12684
rect 3836 10612 3892 10622
rect 3948 10612 4004 12124
rect 3612 9998 3614 10050
rect 3666 9998 3668 10050
rect 3612 9986 3668 9998
rect 3724 10610 4004 10612
rect 3724 10558 3838 10610
rect 3890 10558 4004 10610
rect 3724 10556 4004 10558
rect 4060 12684 4172 12740
rect 3388 9604 3444 9642
rect 3388 9538 3444 9548
rect 3388 9380 3444 9390
rect 3388 9266 3444 9324
rect 3388 9214 3390 9266
rect 3442 9214 3444 9266
rect 3388 9202 3444 9214
rect 3724 9044 3780 10556
rect 3836 10546 3892 10556
rect 3836 9828 3892 9838
rect 3836 9734 3892 9772
rect 4060 9268 4116 12684
rect 4172 12646 4228 12684
rect 4284 10052 4340 14476
rect 4844 14420 4900 14430
rect 4620 14306 4676 14318
rect 4620 14254 4622 14306
rect 4674 14254 4676 14306
rect 4620 13524 4676 14254
rect 4620 13458 4676 13468
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4620 13186 4676 13198
rect 4620 13134 4622 13186
rect 4674 13134 4676 13186
rect 4620 13074 4676 13134
rect 4620 13022 4622 13074
rect 4674 13022 4676 13074
rect 4620 13010 4676 13022
rect 4844 12628 4900 14364
rect 4956 14418 5012 15596
rect 5292 15540 5348 15550
rect 5292 15314 5348 15484
rect 5516 15428 5572 15438
rect 5516 15334 5572 15372
rect 5292 15262 5294 15314
rect 5346 15262 5348 15314
rect 5292 15250 5348 15262
rect 5628 15148 5684 15932
rect 5740 15428 5796 16828
rect 5852 16882 5908 17052
rect 5852 16830 5854 16882
rect 5906 16830 5908 16882
rect 5852 16818 5908 16830
rect 5964 15874 6020 17388
rect 6188 16324 6244 17390
rect 6524 16660 6580 18060
rect 6972 18452 7028 19180
rect 7084 19170 7140 19180
rect 7532 19122 7588 19134
rect 7532 19070 7534 19122
rect 7586 19070 7588 19122
rect 7084 18676 7140 18686
rect 7084 18582 7140 18620
rect 6636 17668 6692 17678
rect 6972 17668 7028 18396
rect 7308 18562 7364 18574
rect 7308 18510 7310 18562
rect 7362 18510 7364 18562
rect 7196 18340 7252 18350
rect 7196 18246 7252 18284
rect 7308 17780 7364 18510
rect 6636 17666 7028 17668
rect 6636 17614 6638 17666
rect 6690 17614 7028 17666
rect 6636 17612 7028 17614
rect 7196 17724 7364 17780
rect 7420 18562 7476 18574
rect 7420 18510 7422 18562
rect 7474 18510 7476 18562
rect 6636 17602 6692 17612
rect 6636 16884 6692 16894
rect 6636 16790 6692 16828
rect 6524 16604 6692 16660
rect 6188 16268 6580 16324
rect 6076 16212 6132 16222
rect 6076 16118 6132 16156
rect 6300 15988 6356 15998
rect 6300 15894 6356 15932
rect 5964 15822 5966 15874
rect 6018 15822 6020 15874
rect 5852 15428 5908 15438
rect 5740 15426 5908 15428
rect 5740 15374 5854 15426
rect 5906 15374 5908 15426
rect 5740 15372 5908 15374
rect 5180 15092 5684 15148
rect 4956 14366 4958 14418
rect 5010 14366 5012 14418
rect 4956 14354 5012 14366
rect 5068 14532 5124 14542
rect 5068 13748 5124 14476
rect 5180 14530 5236 15092
rect 5404 14980 5460 14990
rect 5180 14478 5182 14530
rect 5234 14478 5236 14530
rect 5180 14466 5236 14478
rect 5292 14868 5348 14878
rect 5068 12740 5124 13692
rect 5292 13524 5348 14812
rect 5292 13458 5348 13468
rect 5404 14420 5460 14924
rect 5516 14756 5572 14766
rect 5516 14532 5572 14700
rect 5516 14530 5684 14532
rect 5516 14478 5518 14530
rect 5570 14478 5684 14530
rect 5516 14476 5684 14478
rect 5516 14466 5572 14476
rect 5068 12738 5348 12740
rect 5068 12686 5070 12738
rect 5122 12686 5348 12738
rect 5068 12684 5348 12686
rect 5068 12674 5124 12684
rect 4844 12562 4900 12572
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 5068 11620 5124 11630
rect 5068 11506 5124 11564
rect 5068 11454 5070 11506
rect 5122 11454 5124 11506
rect 5068 11442 5124 11454
rect 4508 11172 4564 11182
rect 4508 10722 4564 11116
rect 4508 10670 4510 10722
rect 4562 10670 4564 10722
rect 4508 10658 4564 10670
rect 5292 10276 5348 12684
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 5292 10210 5348 10220
rect 4476 10154 4740 10164
rect 4284 9996 4676 10052
rect 4620 9938 4676 9996
rect 4620 9886 4622 9938
rect 4674 9886 4676 9938
rect 4620 9874 4676 9886
rect 4284 9602 4340 9614
rect 4284 9550 4286 9602
rect 4338 9550 4340 9602
rect 4060 9202 4116 9212
rect 4172 9380 4228 9390
rect 3500 9042 3780 9044
rect 3500 8990 3726 9042
rect 3778 8990 3780 9042
rect 3500 8988 3780 8990
rect 3276 8820 3332 8830
rect 3276 8726 3332 8764
rect 3276 8372 3332 8382
rect 1932 8370 2436 8372
rect 1932 8318 1934 8370
rect 1986 8318 2436 8370
rect 1932 8316 2436 8318
rect 2492 8370 3332 8372
rect 2492 8318 3278 8370
rect 3330 8318 3332 8370
rect 2492 8316 3332 8318
rect 1932 8306 1988 8316
rect 2380 8148 2436 8158
rect 2492 8148 2548 8316
rect 2380 8146 2548 8148
rect 2380 8094 2382 8146
rect 2434 8094 2548 8146
rect 2380 8092 2548 8094
rect 2380 8082 2436 8092
rect 2828 8036 2884 8046
rect 2828 7942 2884 7980
rect 1820 7700 1876 7710
rect 1708 7698 1876 7700
rect 1708 7646 1822 7698
rect 1874 7646 1876 7698
rect 1708 7644 1876 7646
rect 1820 7634 1876 7644
rect 2716 7362 2772 7374
rect 2716 7310 2718 7362
rect 2770 7310 2772 7362
rect 2716 6916 2772 7310
rect 3164 7364 3220 7374
rect 3164 7270 3220 7308
rect 2716 6850 2772 6860
rect 2828 6914 2884 6926
rect 2828 6862 2830 6914
rect 2882 6862 2884 6914
rect 2828 6802 2884 6862
rect 2828 6750 2830 6802
rect 2882 6750 2884 6802
rect 2828 6738 2884 6750
rect 3276 6356 3332 8316
rect 3500 7474 3556 8988
rect 3724 8978 3780 8988
rect 4060 8372 4116 8382
rect 3724 8260 3780 8270
rect 3724 8166 3780 8204
rect 3500 7422 3502 7474
rect 3554 7422 3556 7474
rect 3500 6914 3556 7422
rect 3500 6862 3502 6914
rect 3554 6862 3556 6914
rect 3388 6580 3444 6590
rect 3388 6486 3444 6524
rect 3276 6300 3388 6356
rect 3332 6244 3388 6300
rect 3332 6188 3444 6244
rect 3388 2884 3444 6188
rect 3500 6132 3556 6862
rect 3836 6692 3892 6702
rect 3836 6598 3892 6636
rect 3500 6130 3892 6132
rect 3500 6078 3502 6130
rect 3554 6078 3892 6130
rect 3500 6076 3892 6078
rect 3500 6066 3556 6076
rect 3836 5906 3892 6076
rect 3836 5854 3838 5906
rect 3890 5854 3892 5906
rect 3836 5236 3892 5854
rect 3836 5170 3892 5180
rect 4060 3332 4116 8316
rect 4172 8370 4228 9324
rect 4284 9156 4340 9550
rect 5068 9602 5124 9614
rect 5068 9550 5070 9602
rect 5122 9550 5124 9602
rect 5068 9492 5124 9550
rect 5068 9426 5124 9436
rect 4284 9090 4340 9100
rect 5404 9044 5460 14364
rect 5516 13524 5572 13534
rect 5516 9492 5572 13468
rect 5628 13076 5684 14476
rect 5740 14308 5796 14318
rect 5740 14214 5796 14252
rect 5852 13188 5908 15372
rect 5964 14756 6020 15822
rect 6188 15876 6244 15886
rect 6188 15782 6244 15820
rect 6412 15316 6468 15326
rect 6412 15222 6468 15260
rect 6300 15204 6356 15214
rect 6300 14980 6356 15148
rect 6300 14914 6356 14924
rect 6524 14868 6580 16268
rect 6636 16100 6692 16604
rect 6636 16034 6692 16044
rect 6748 16098 6804 17612
rect 7196 17444 7252 17724
rect 7196 16996 7252 17388
rect 7308 17554 7364 17566
rect 7308 17502 7310 17554
rect 7362 17502 7364 17554
rect 7308 17332 7364 17502
rect 7308 17266 7364 17276
rect 7420 17220 7476 18510
rect 7532 18004 7588 19070
rect 7644 19122 7700 19404
rect 7756 19348 7812 19628
rect 7868 19572 7924 19966
rect 8092 19908 8148 19918
rect 8092 19814 8148 19852
rect 7868 19506 7924 19516
rect 7756 19292 8036 19348
rect 7644 19070 7646 19122
rect 7698 19070 7700 19122
rect 7644 19058 7700 19070
rect 7756 19124 7812 19134
rect 7756 19030 7812 19068
rect 7868 19010 7924 19022
rect 7868 18958 7870 19010
rect 7922 18958 7924 19010
rect 7644 18562 7700 18574
rect 7644 18510 7646 18562
rect 7698 18510 7700 18562
rect 7644 18452 7700 18510
rect 7644 18386 7700 18396
rect 7532 17938 7588 17948
rect 7420 17154 7476 17164
rect 7532 17554 7588 17566
rect 7532 17502 7534 17554
rect 7586 17502 7588 17554
rect 7196 16930 7252 16940
rect 6748 16046 6750 16098
rect 6802 16046 6804 16098
rect 6748 15988 6804 16046
rect 6748 15922 6804 15932
rect 7196 16212 7252 16222
rect 6860 15876 6916 15886
rect 6860 15314 6916 15820
rect 6860 15262 6862 15314
rect 6914 15262 6916 15314
rect 6860 15250 6916 15262
rect 7196 15204 7252 16156
rect 7308 16100 7364 16110
rect 7308 16006 7364 16044
rect 7196 15138 7252 15148
rect 7420 15428 7476 15438
rect 6524 14802 6580 14812
rect 5964 14690 6020 14700
rect 6076 14644 6132 14654
rect 5964 14420 6020 14430
rect 5964 14326 6020 14364
rect 6076 14308 6132 14588
rect 7084 14530 7140 14542
rect 7084 14478 7086 14530
rect 7138 14478 7140 14530
rect 6188 14420 6244 14430
rect 6412 14420 6468 14430
rect 6188 14418 6412 14420
rect 6188 14366 6190 14418
rect 6242 14366 6412 14418
rect 6188 14364 6412 14366
rect 6188 14354 6244 14364
rect 6412 14354 6468 14364
rect 6636 14420 6692 14430
rect 6636 14326 6692 14364
rect 6076 14242 6132 14252
rect 6524 14308 6580 14318
rect 6524 13972 6580 14252
rect 6748 14308 6804 14318
rect 6748 14306 7028 14308
rect 6748 14254 6750 14306
rect 6802 14254 7028 14306
rect 6748 14252 7028 14254
rect 6748 14242 6804 14252
rect 6636 13972 6692 13982
rect 6524 13970 6692 13972
rect 6524 13918 6638 13970
rect 6690 13918 6692 13970
rect 6524 13916 6692 13918
rect 6636 13906 6692 13916
rect 6860 13746 6916 13758
rect 6860 13694 6862 13746
rect 6914 13694 6916 13746
rect 6300 13634 6356 13646
rect 6300 13582 6302 13634
rect 6354 13582 6356 13634
rect 6300 13524 6356 13582
rect 6748 13634 6804 13646
rect 6748 13582 6750 13634
rect 6802 13582 6804 13634
rect 6748 13524 6804 13582
rect 6300 13458 6356 13468
rect 6636 13468 6804 13524
rect 5852 13122 5908 13132
rect 6412 13300 6468 13310
rect 5628 13020 5796 13076
rect 5628 11394 5684 13020
rect 5740 12964 5796 13020
rect 5964 12964 6020 12974
rect 5740 12962 6020 12964
rect 5740 12910 5966 12962
rect 6018 12910 6020 12962
rect 5740 12908 6020 12910
rect 5964 12898 6020 12908
rect 6412 12964 6468 13244
rect 6412 12962 6580 12964
rect 6412 12910 6414 12962
rect 6466 12910 6580 12962
rect 6412 12908 6580 12910
rect 6412 12898 6468 12908
rect 5628 11342 5630 11394
rect 5682 11342 5684 11394
rect 5628 10724 5684 11342
rect 5628 10658 5684 10668
rect 5740 12738 5796 12750
rect 5740 12686 5742 12738
rect 5794 12686 5796 12738
rect 5740 12516 5796 12686
rect 5516 9426 5572 9436
rect 5740 9380 5796 12460
rect 6188 12738 6244 12750
rect 6188 12686 6190 12738
rect 6242 12686 6244 12738
rect 6188 12292 6244 12686
rect 6188 12226 6244 12236
rect 6412 12180 6468 12190
rect 5964 12066 6020 12078
rect 5964 12014 5966 12066
rect 6018 12014 6020 12066
rect 5964 11956 6020 12014
rect 5964 11890 6020 11900
rect 6412 12066 6468 12124
rect 6412 12014 6414 12066
rect 6466 12014 6468 12066
rect 6412 11732 6468 12014
rect 5964 11676 6468 11732
rect 5852 11172 5908 11182
rect 5852 11078 5908 11116
rect 5964 9716 6020 11676
rect 6300 11396 6356 11406
rect 6300 11302 6356 11340
rect 5964 9650 6020 9660
rect 6076 11282 6132 11294
rect 6076 11230 6078 11282
rect 6130 11230 6132 11282
rect 6076 11060 6132 11230
rect 5740 9314 5796 9324
rect 5404 8978 5460 8988
rect 5516 9268 5572 9278
rect 4396 8932 4452 8942
rect 4956 8932 5012 8942
rect 4396 8930 4900 8932
rect 4396 8878 4398 8930
rect 4450 8878 4900 8930
rect 4396 8876 4900 8878
rect 4396 8866 4452 8876
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4844 8482 4900 8876
rect 4844 8430 4846 8482
rect 4898 8430 4900 8482
rect 4844 8418 4900 8430
rect 4172 8318 4174 8370
rect 4226 8318 4228 8370
rect 4172 8306 4228 8318
rect 4956 8370 5012 8876
rect 4956 8318 4958 8370
rect 5010 8318 5012 8370
rect 4956 8306 5012 8318
rect 4620 8034 4676 8046
rect 4620 7982 4622 8034
rect 4674 7982 4676 8034
rect 4620 7924 4676 7982
rect 4620 7858 4676 7868
rect 4172 7588 4228 7598
rect 4172 7494 4228 7532
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4620 6914 4676 6926
rect 4620 6862 4622 6914
rect 4674 6862 4676 6914
rect 4620 6802 4676 6862
rect 4620 6750 4622 6802
rect 4674 6750 4676 6802
rect 4620 6738 4676 6750
rect 4284 6580 4340 6590
rect 4284 6486 4340 6524
rect 5516 6580 5572 9212
rect 5740 8148 5796 8158
rect 5740 8054 5796 8092
rect 5852 8146 5908 8158
rect 5852 8094 5854 8146
rect 5906 8094 5908 8146
rect 5628 8034 5684 8046
rect 5628 7982 5630 8034
rect 5682 7982 5684 8034
rect 5628 7588 5684 7982
rect 5628 7522 5684 7532
rect 5516 6514 5572 6524
rect 5852 6690 5908 8094
rect 5852 6638 5854 6690
rect 5906 6638 5908 6690
rect 5852 6580 5908 6638
rect 5852 6514 5908 6524
rect 5964 7028 6020 7038
rect 5180 6466 5236 6478
rect 5180 6414 5182 6466
rect 5234 6414 5236 6466
rect 5180 6244 5236 6414
rect 5180 6178 5236 6188
rect 4620 5796 4676 5806
rect 4620 5702 4676 5740
rect 5628 5796 5684 5806
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 5628 5346 5684 5740
rect 5628 5294 5630 5346
rect 5682 5294 5684 5346
rect 5628 5282 5684 5294
rect 5740 5348 5796 5358
rect 4620 5236 4676 5246
rect 4620 5142 4676 5180
rect 5068 5236 5124 5246
rect 5124 5180 5348 5236
rect 5068 5142 5124 5180
rect 5292 4562 5348 5180
rect 5740 5234 5796 5292
rect 5740 5182 5742 5234
rect 5794 5182 5796 5234
rect 5740 5170 5796 5182
rect 5292 4510 5294 4562
rect 5346 4510 5348 4562
rect 5292 4498 5348 4510
rect 5852 4564 5908 4574
rect 5964 4564 6020 6972
rect 6076 6468 6132 11004
rect 6188 10500 6244 10510
rect 6188 9938 6244 10444
rect 6188 9886 6190 9938
rect 6242 9886 6244 9938
rect 6188 9874 6244 9886
rect 6412 9268 6468 9278
rect 6524 9268 6580 12908
rect 6636 12962 6692 13468
rect 6860 13300 6916 13694
rect 6972 13524 7028 14252
rect 7084 13972 7140 14478
rect 7084 13970 7364 13972
rect 7084 13918 7086 13970
rect 7138 13918 7364 13970
rect 7084 13916 7364 13918
rect 7084 13906 7140 13916
rect 6972 13458 7028 13468
rect 6860 13244 7252 13300
rect 6636 12910 6638 12962
rect 6690 12910 6692 12962
rect 6636 12898 6692 12910
rect 7084 13076 7140 13086
rect 7084 12962 7140 13020
rect 7084 12910 7086 12962
rect 7138 12910 7140 12962
rect 7084 12898 7140 12910
rect 7084 12516 7140 12526
rect 6748 12404 6804 12414
rect 6636 12348 6748 12404
rect 6636 11170 6692 12348
rect 6748 12310 6804 12348
rect 6972 12178 7028 12190
rect 6972 12126 6974 12178
rect 7026 12126 7028 12178
rect 6860 12066 6916 12078
rect 6860 12014 6862 12066
rect 6914 12014 6916 12066
rect 6860 11732 6916 12014
rect 6860 11666 6916 11676
rect 6972 11620 7028 12126
rect 6748 11396 6804 11406
rect 6748 11302 6804 11340
rect 6636 11118 6638 11170
rect 6690 11118 6692 11170
rect 6636 11106 6692 11118
rect 6860 11170 6916 11182
rect 6860 11118 6862 11170
rect 6914 11118 6916 11170
rect 6636 10500 6692 10510
rect 6860 10500 6916 11118
rect 6972 11172 7028 11564
rect 7084 11282 7140 12460
rect 7196 11956 7252 13244
rect 7308 12292 7364 13916
rect 7420 13746 7476 15372
rect 7532 15148 7588 17502
rect 7756 17556 7812 17566
rect 7756 17462 7812 17500
rect 7868 17554 7924 18958
rect 7868 17502 7870 17554
rect 7922 17502 7924 17554
rect 7644 17444 7700 17454
rect 7644 17350 7700 17388
rect 7868 17444 7924 17502
rect 7868 17378 7924 17388
rect 7868 16212 7924 16222
rect 7980 16212 8036 19292
rect 8428 19236 8484 19246
rect 8316 19180 8428 19236
rect 7868 16210 8036 16212
rect 7868 16158 7870 16210
rect 7922 16158 8036 16210
rect 7868 16156 8036 16158
rect 8092 18004 8148 18014
rect 7644 15988 7700 15998
rect 7644 15538 7700 15932
rect 7868 15764 7924 16156
rect 7868 15698 7924 15708
rect 7644 15486 7646 15538
rect 7698 15486 7700 15538
rect 7644 15474 7700 15486
rect 7868 15316 7924 15326
rect 7532 15092 7700 15148
rect 7532 14306 7588 14318
rect 7532 14254 7534 14306
rect 7586 14254 7588 14306
rect 7532 14084 7588 14254
rect 7532 14018 7588 14028
rect 7644 13748 7700 15092
rect 7868 14642 7924 15260
rect 7980 15314 8036 15326
rect 7980 15262 7982 15314
rect 8034 15262 8036 15314
rect 7980 15204 8036 15262
rect 7980 15138 8036 15148
rect 7868 14590 7870 14642
rect 7922 14590 7924 14642
rect 7868 14578 7924 14590
rect 7756 14532 7812 14542
rect 7756 14438 7812 14476
rect 7980 14308 8036 14318
rect 7868 14196 7924 14206
rect 7420 13694 7422 13746
rect 7474 13694 7476 13746
rect 7420 12404 7476 13694
rect 7532 13692 7700 13748
rect 7756 13970 7812 13982
rect 7756 13918 7758 13970
rect 7810 13918 7812 13970
rect 7532 12852 7588 13692
rect 7644 13524 7700 13534
rect 7644 12852 7700 13468
rect 7756 13074 7812 13918
rect 7756 13022 7758 13074
rect 7810 13022 7812 13074
rect 7756 13010 7812 13022
rect 7868 13746 7924 14140
rect 7980 13972 8036 14252
rect 7980 13906 8036 13916
rect 7868 13694 7870 13746
rect 7922 13694 7924 13746
rect 7644 12796 7812 12852
rect 7532 12786 7588 12796
rect 7420 12338 7476 12348
rect 7644 12628 7700 12638
rect 7644 12402 7700 12572
rect 7644 12350 7646 12402
rect 7698 12350 7700 12402
rect 7644 12338 7700 12350
rect 7308 12178 7364 12236
rect 7308 12126 7310 12178
rect 7362 12126 7364 12178
rect 7308 12114 7364 12126
rect 7756 12068 7812 12796
rect 7868 12180 7924 13694
rect 7980 13746 8036 13758
rect 7980 13694 7982 13746
rect 8034 13694 8036 13746
rect 7980 13524 8036 13694
rect 7980 13458 8036 13468
rect 7868 12114 7924 12124
rect 7980 12740 8036 12750
rect 7980 12402 8036 12684
rect 7980 12350 7982 12402
rect 8034 12350 8036 12402
rect 7644 12012 7812 12068
rect 7196 11890 7252 11900
rect 7532 11956 7588 11966
rect 7196 11732 7252 11742
rect 7252 11676 7476 11732
rect 7196 11666 7252 11676
rect 7084 11230 7086 11282
rect 7138 11230 7140 11282
rect 7084 11218 7140 11230
rect 6972 11106 7028 11116
rect 7196 10836 7252 10874
rect 7196 10770 7252 10780
rect 6972 10724 7028 10734
rect 6972 10630 7028 10668
rect 6636 10498 6916 10500
rect 6636 10446 6638 10498
rect 6690 10446 6916 10498
rect 6636 10444 6916 10446
rect 7308 10610 7364 10622
rect 7308 10558 7310 10610
rect 7362 10558 7364 10610
rect 6636 10434 6692 10444
rect 6468 9212 6580 9268
rect 6636 10276 6692 10286
rect 6636 9602 6692 10220
rect 6636 9550 6638 9602
rect 6690 9550 6692 9602
rect 6412 9202 6468 9212
rect 6524 9044 6580 9054
rect 6524 8930 6580 8988
rect 6524 8878 6526 8930
rect 6578 8878 6580 8930
rect 6524 8866 6580 8878
rect 6636 8708 6692 9550
rect 6524 8652 6692 8708
rect 6412 8370 6468 8382
rect 6412 8318 6414 8370
rect 6466 8318 6468 8370
rect 6300 8260 6356 8270
rect 6300 7588 6356 8204
rect 6412 8258 6468 8318
rect 6412 8206 6414 8258
rect 6466 8206 6468 8258
rect 6412 8194 6468 8206
rect 6524 7812 6580 8652
rect 6748 8260 6804 10444
rect 6972 10164 7028 10174
rect 6860 10108 6972 10164
rect 6860 8484 6916 10108
rect 6972 10098 7028 10108
rect 7308 10164 7364 10558
rect 7420 10610 7476 11676
rect 7532 11506 7588 11900
rect 7532 11454 7534 11506
rect 7586 11454 7588 11506
rect 7532 11442 7588 11454
rect 7644 11284 7700 12012
rect 7868 11732 7924 11742
rect 7756 11676 7868 11732
rect 7756 11618 7812 11676
rect 7756 11566 7758 11618
rect 7810 11566 7812 11618
rect 7756 11554 7812 11566
rect 7420 10558 7422 10610
rect 7474 10558 7476 10610
rect 7420 10546 7476 10558
rect 7532 11228 7700 11284
rect 7308 10098 7364 10108
rect 7308 9716 7364 9726
rect 7196 9714 7364 9716
rect 7196 9662 7310 9714
rect 7362 9662 7364 9714
rect 7196 9660 7364 9662
rect 6972 9602 7028 9614
rect 6972 9550 6974 9602
rect 7026 9550 7028 9602
rect 6972 9268 7028 9550
rect 6972 9202 7028 9212
rect 7196 9044 7252 9660
rect 7308 9650 7364 9660
rect 7532 9714 7588 11228
rect 7532 9662 7534 9714
rect 7586 9662 7588 9714
rect 7532 9650 7588 9662
rect 7644 9940 7700 9950
rect 7644 9602 7700 9884
rect 7868 9826 7924 11676
rect 7868 9774 7870 9826
rect 7922 9774 7924 9826
rect 7868 9716 7924 9774
rect 7868 9650 7924 9660
rect 7644 9550 7646 9602
rect 7698 9550 7700 9602
rect 7532 9492 7588 9502
rect 7196 8978 7252 8988
rect 7308 9436 7532 9492
rect 7308 9266 7364 9436
rect 7532 9426 7588 9436
rect 7308 9214 7310 9266
rect 7362 9214 7364 9266
rect 7308 8484 7364 9214
rect 7532 9156 7588 9166
rect 7644 9156 7700 9550
rect 7980 9492 8036 12350
rect 8092 12404 8148 17948
rect 8204 17668 8260 17678
rect 8316 17668 8372 19180
rect 8428 19142 8484 19180
rect 8540 18452 8596 20972
rect 8652 20802 8708 25566
rect 8988 26290 9044 26852
rect 8988 26238 8990 26290
rect 9042 26238 9044 26290
rect 8988 24162 9044 26238
rect 8988 24110 8990 24162
rect 9042 24110 9044 24162
rect 8988 24098 9044 24110
rect 8652 20750 8654 20802
rect 8706 20750 8708 20802
rect 8652 20738 8708 20750
rect 9100 19124 9156 19134
rect 9100 19030 9156 19068
rect 8652 18452 8708 18462
rect 8540 18450 8708 18452
rect 8540 18398 8654 18450
rect 8706 18398 8708 18450
rect 8540 18396 8708 18398
rect 8428 18228 8484 18238
rect 8428 18134 8484 18172
rect 8260 17612 8372 17668
rect 8204 17574 8260 17612
rect 8428 16884 8484 16894
rect 8316 16212 8372 16222
rect 8204 16210 8372 16212
rect 8204 16158 8318 16210
rect 8370 16158 8372 16210
rect 8204 16156 8372 16158
rect 8204 14420 8260 16156
rect 8316 16146 8372 16156
rect 8428 15538 8484 16828
rect 8652 16660 8708 18396
rect 8988 17556 9044 17566
rect 8988 17462 9044 17500
rect 9212 16884 9268 28140
rect 9884 28082 9940 28476
rect 10108 28196 10164 28702
rect 10108 28130 10164 28140
rect 10220 29538 10276 29550
rect 10220 29486 10222 29538
rect 10274 29486 10276 29538
rect 9884 28030 9886 28082
rect 9938 28030 9940 28082
rect 9884 28018 9940 28030
rect 10220 28082 10276 29486
rect 10332 29092 10388 30158
rect 10444 29988 10500 35308
rect 10556 33348 10612 33358
rect 10780 33348 10836 37212
rect 11004 37202 11060 37212
rect 10892 36594 10948 36606
rect 10892 36542 10894 36594
rect 10946 36542 10948 36594
rect 10892 35924 10948 36542
rect 10892 35858 10948 35868
rect 11004 35140 11060 35150
rect 10892 35026 10948 35038
rect 10892 34974 10894 35026
rect 10946 34974 10948 35026
rect 10892 33796 10948 34974
rect 11004 34802 11060 35084
rect 11116 35028 11172 37436
rect 11340 37268 11396 38612
rect 12012 38052 12068 38670
rect 12124 38668 12180 40684
rect 12460 40516 12516 40526
rect 12348 40460 12460 40516
rect 12348 39618 12404 40460
rect 12460 40450 12516 40460
rect 12572 40516 12628 40526
rect 12684 40516 12740 40684
rect 14028 40628 14084 40910
rect 14028 40562 14084 40572
rect 12572 40514 12740 40516
rect 12572 40462 12574 40514
rect 12626 40462 12740 40514
rect 12572 40460 12740 40462
rect 13468 40516 13524 40526
rect 12572 40180 12628 40460
rect 13468 40422 13524 40460
rect 13132 40404 13188 40414
rect 13132 40310 13188 40348
rect 13580 40292 13636 40302
rect 13580 40198 13636 40236
rect 12348 39566 12350 39618
rect 12402 39566 12404 39618
rect 12348 39554 12404 39566
rect 12460 40124 12628 40180
rect 12124 38612 12404 38668
rect 12012 37996 12292 38052
rect 11564 37828 11620 37838
rect 11564 37734 11620 37772
rect 11900 37826 11956 37838
rect 11900 37774 11902 37826
rect 11954 37774 11956 37826
rect 11340 36482 11396 37212
rect 11900 37380 11956 37774
rect 11340 36430 11342 36482
rect 11394 36430 11396 36482
rect 11340 36418 11396 36430
rect 11788 37154 11844 37166
rect 11788 37102 11790 37154
rect 11842 37102 11844 37154
rect 11788 36260 11844 37102
rect 11900 36482 11956 37324
rect 11900 36430 11902 36482
rect 11954 36430 11956 36482
rect 11900 36418 11956 36430
rect 12012 37826 12068 37838
rect 12012 37774 12014 37826
rect 12066 37774 12068 37826
rect 12012 36484 12068 37774
rect 12124 37828 12180 37838
rect 12124 37268 12180 37772
rect 12236 37380 12292 37996
rect 12348 37492 12404 38612
rect 12460 38050 12516 40124
rect 13020 39620 13076 39630
rect 13020 39526 13076 39564
rect 13804 39620 13860 39630
rect 12572 39508 12628 39518
rect 12572 39506 12740 39508
rect 12572 39454 12574 39506
rect 12626 39454 12740 39506
rect 12572 39452 12740 39454
rect 12572 39442 12628 39452
rect 12684 38948 12740 39452
rect 13468 39506 13524 39518
rect 13468 39454 13470 39506
rect 13522 39454 13524 39506
rect 12796 39394 12852 39406
rect 12796 39342 12798 39394
rect 12850 39342 12852 39394
rect 12796 39060 12852 39342
rect 12796 39004 13188 39060
rect 12684 38892 12964 38948
rect 12572 38722 12628 38734
rect 12572 38670 12574 38722
rect 12626 38670 12628 38722
rect 12572 38668 12628 38670
rect 12572 38612 12852 38668
rect 12460 37998 12462 38050
rect 12514 37998 12516 38050
rect 12460 37986 12516 37998
rect 12348 37436 12628 37492
rect 12236 37324 12404 37380
rect 12124 37202 12180 37212
rect 12348 37156 12404 37324
rect 12012 36418 12068 36428
rect 12236 37100 12404 37156
rect 12460 37268 12516 37278
rect 12124 36260 12180 36270
rect 11788 36258 12180 36260
rect 11788 36206 12126 36258
rect 12178 36206 12180 36258
rect 11788 36204 12180 36206
rect 12124 36194 12180 36204
rect 11788 35810 11844 35822
rect 11788 35758 11790 35810
rect 11842 35758 11844 35810
rect 11228 35698 11284 35710
rect 11228 35646 11230 35698
rect 11282 35646 11284 35698
rect 11228 35476 11284 35646
rect 11788 35588 11844 35758
rect 11788 35522 11844 35532
rect 11900 35700 11956 35710
rect 12124 35700 12180 35710
rect 11900 35586 11956 35644
rect 11900 35534 11902 35586
rect 11954 35534 11956 35586
rect 11900 35522 11956 35534
rect 12012 35698 12180 35700
rect 12012 35646 12126 35698
rect 12178 35646 12180 35698
rect 12012 35644 12180 35646
rect 11564 35476 11620 35486
rect 11228 35474 11620 35476
rect 11228 35422 11566 35474
rect 11618 35422 11620 35474
rect 11228 35420 11620 35422
rect 11116 34962 11172 34972
rect 11004 34750 11006 34802
rect 11058 34750 11060 34802
rect 11004 34738 11060 34750
rect 11228 34802 11284 34814
rect 11228 34750 11230 34802
rect 11282 34750 11284 34802
rect 11116 34692 11172 34702
rect 11116 34130 11172 34636
rect 11116 34078 11118 34130
rect 11170 34078 11172 34130
rect 11004 34020 11060 34030
rect 11004 33926 11060 33964
rect 10892 33730 10948 33740
rect 10892 33348 10948 33358
rect 10780 33346 10948 33348
rect 10780 33294 10894 33346
rect 10946 33294 10948 33346
rect 10780 33292 10948 33294
rect 10556 30212 10612 33292
rect 10892 32452 10948 33292
rect 10892 32386 10948 32396
rect 11004 32676 11060 32686
rect 10892 32116 10948 32126
rect 10556 30146 10612 30156
rect 10780 30210 10836 30222
rect 10780 30158 10782 30210
rect 10834 30158 10836 30210
rect 10668 30098 10724 30110
rect 10668 30046 10670 30098
rect 10722 30046 10724 30098
rect 10444 29932 10612 29988
rect 10556 29652 10612 29932
rect 10556 29586 10612 29596
rect 10332 29026 10388 29036
rect 10444 29540 10500 29550
rect 10220 28030 10222 28082
rect 10274 28030 10276 28082
rect 10220 28018 10276 28030
rect 9660 27970 9716 27982
rect 9660 27918 9662 27970
rect 9714 27918 9716 27970
rect 9548 27858 9604 27870
rect 9548 27806 9550 27858
rect 9602 27806 9604 27858
rect 9436 25394 9492 25406
rect 9436 25342 9438 25394
rect 9490 25342 9492 25394
rect 9436 25172 9492 25342
rect 9548 25396 9604 27806
rect 9660 27860 9716 27918
rect 9660 27524 9716 27804
rect 10108 27972 10164 27982
rect 10108 27858 10164 27916
rect 10108 27806 10110 27858
rect 10162 27806 10164 27858
rect 10108 27794 10164 27806
rect 9660 27458 9716 27468
rect 10332 27076 10388 27086
rect 9548 25330 9604 25340
rect 10220 26402 10276 26414
rect 10220 26350 10222 26402
rect 10274 26350 10276 26402
rect 10220 25396 10276 26350
rect 10220 25330 10276 25340
rect 9436 25116 9716 25172
rect 9548 24948 9604 24958
rect 9436 24722 9492 24734
rect 9436 24670 9438 24722
rect 9490 24670 9492 24722
rect 9436 21588 9492 24670
rect 9548 23266 9604 24892
rect 9660 23940 9716 25116
rect 9772 24948 9828 24958
rect 9772 24946 10052 24948
rect 9772 24894 9774 24946
rect 9826 24894 10052 24946
rect 9772 24892 10052 24894
rect 9772 24882 9828 24892
rect 9660 23846 9716 23884
rect 9884 24722 9940 24734
rect 9884 24670 9886 24722
rect 9938 24670 9940 24722
rect 9548 23214 9550 23266
rect 9602 23214 9604 23266
rect 9548 23202 9604 23214
rect 9660 23268 9716 23278
rect 9660 21812 9716 23212
rect 9772 21812 9828 21822
rect 9660 21810 9828 21812
rect 9660 21758 9774 21810
rect 9826 21758 9828 21810
rect 9660 21756 9828 21758
rect 9772 21746 9828 21756
rect 9660 21588 9716 21598
rect 9436 21586 9716 21588
rect 9436 21534 9662 21586
rect 9714 21534 9716 21586
rect 9436 21532 9716 21534
rect 9548 18004 9604 21532
rect 9660 21522 9716 21532
rect 9884 21588 9940 24670
rect 9996 22482 10052 24892
rect 10108 24722 10164 24734
rect 10108 24670 10110 24722
rect 10162 24670 10164 24722
rect 10108 23268 10164 24670
rect 10108 23202 10164 23212
rect 10220 23380 10276 23390
rect 9996 22430 9998 22482
rect 10050 22430 10052 22482
rect 9996 22418 10052 22430
rect 10108 22930 10164 22942
rect 10108 22878 10110 22930
rect 10162 22878 10164 22930
rect 9884 21586 10052 21588
rect 9884 21534 9886 21586
rect 9938 21534 10052 21586
rect 9884 21532 10052 21534
rect 9884 21522 9940 21532
rect 9772 20916 9828 20926
rect 9772 20802 9828 20860
rect 9772 20750 9774 20802
rect 9826 20750 9828 20802
rect 9772 20738 9828 20750
rect 9884 20468 9940 20478
rect 9884 20242 9940 20412
rect 9884 20190 9886 20242
rect 9938 20190 9940 20242
rect 9884 20178 9940 20190
rect 9996 20244 10052 21532
rect 9884 20020 9940 20058
rect 9884 19954 9940 19964
rect 9996 19796 10052 20188
rect 9884 19740 10052 19796
rect 9660 18450 9716 18462
rect 9660 18398 9662 18450
rect 9714 18398 9716 18450
rect 9660 18228 9716 18398
rect 9660 18162 9716 18172
rect 9548 17948 9716 18004
rect 9548 16884 9604 16894
rect 9212 16882 9604 16884
rect 9212 16830 9550 16882
rect 9602 16830 9604 16882
rect 9212 16828 9604 16830
rect 9548 16818 9604 16828
rect 8764 16772 8820 16782
rect 8764 16770 9268 16772
rect 8764 16718 8766 16770
rect 8818 16718 9268 16770
rect 8764 16716 9268 16718
rect 8764 16706 8820 16716
rect 8652 16594 8708 16604
rect 8428 15486 8430 15538
rect 8482 15486 8484 15538
rect 8428 15474 8484 15486
rect 8316 15428 8372 15438
rect 8316 15334 8372 15372
rect 8652 15314 8708 15326
rect 8652 15262 8654 15314
rect 8706 15262 8708 15314
rect 8204 14354 8260 14364
rect 8316 14756 8372 14766
rect 8316 14418 8372 14700
rect 8316 14366 8318 14418
rect 8370 14366 8372 14418
rect 8316 14354 8372 14366
rect 8540 14530 8596 14542
rect 8540 14478 8542 14530
rect 8594 14478 8596 14530
rect 8540 14084 8596 14478
rect 8316 14028 8596 14084
rect 8092 12338 8148 12348
rect 8204 13076 8260 13086
rect 8092 11396 8148 11406
rect 8092 11302 8148 11340
rect 8092 10836 8148 10846
rect 8204 10836 8260 13020
rect 8316 12740 8372 14028
rect 8652 13972 8708 15262
rect 8764 15316 8820 15326
rect 8764 15222 8820 15260
rect 8988 15204 9044 15214
rect 8652 13906 8708 13916
rect 8764 15092 9044 15148
rect 8428 13748 8484 13758
rect 8428 13654 8484 13692
rect 8540 13746 8596 13758
rect 8540 13694 8542 13746
rect 8594 13694 8596 13746
rect 8540 13524 8596 13694
rect 8540 13458 8596 13468
rect 8652 13746 8708 13758
rect 8652 13694 8654 13746
rect 8706 13694 8708 13746
rect 8652 13188 8708 13694
rect 8652 13122 8708 13132
rect 8316 12674 8372 12684
rect 8764 12516 8820 15092
rect 9100 14530 9156 14542
rect 9100 14478 9102 14530
rect 9154 14478 9156 14530
rect 9100 14420 9156 14478
rect 9212 14532 9268 16716
rect 9436 14644 9492 14654
rect 9436 14550 9492 14588
rect 9212 14438 9268 14476
rect 9660 14530 9716 17948
rect 9884 15652 9940 19740
rect 10108 19684 10164 22878
rect 10220 21924 10276 23324
rect 10220 21586 10276 21868
rect 10220 21534 10222 21586
rect 10274 21534 10276 21586
rect 10220 21522 10276 21534
rect 10332 21026 10388 27020
rect 10444 27074 10500 29484
rect 10556 29428 10612 29438
rect 10668 29428 10724 30046
rect 10556 29426 10724 29428
rect 10556 29374 10558 29426
rect 10610 29374 10724 29426
rect 10556 29372 10724 29374
rect 10556 28756 10612 29372
rect 10556 28690 10612 28700
rect 10668 29204 10724 29214
rect 10668 28530 10724 29148
rect 10668 28478 10670 28530
rect 10722 28478 10724 28530
rect 10668 28420 10724 28478
rect 10668 28354 10724 28364
rect 10780 27972 10836 30158
rect 10780 27906 10836 27916
rect 10892 27636 10948 32060
rect 11004 30100 11060 32620
rect 11116 32564 11172 34078
rect 11228 32788 11284 34750
rect 11564 33348 11620 35420
rect 11900 35140 11956 35150
rect 11676 34914 11732 34926
rect 11676 34862 11678 34914
rect 11730 34862 11732 34914
rect 11676 34692 11732 34862
rect 11900 34802 11956 35084
rect 11900 34750 11902 34802
rect 11954 34750 11956 34802
rect 11900 34738 11956 34750
rect 12012 34804 12068 35644
rect 12124 35634 12180 35644
rect 12236 34916 12292 37100
rect 12460 36932 12516 37212
rect 12348 36876 12516 36932
rect 12348 36482 12404 36876
rect 12348 36430 12350 36482
rect 12402 36430 12404 36482
rect 12348 36418 12404 36430
rect 12460 36484 12516 36494
rect 12460 36390 12516 36428
rect 12572 35924 12628 37436
rect 12796 37380 12852 38612
rect 12908 38052 12964 38892
rect 13020 38836 13076 38846
rect 13020 38742 13076 38780
rect 13132 38722 13188 39004
rect 13132 38670 13134 38722
rect 13186 38670 13188 38722
rect 13132 38658 13188 38670
rect 12908 37604 12964 37996
rect 13020 37828 13076 37838
rect 13020 37826 13188 37828
rect 13020 37774 13022 37826
rect 13074 37774 13188 37826
rect 13020 37772 13188 37774
rect 13020 37762 13076 37772
rect 12908 37538 12964 37548
rect 13020 37380 13076 37390
rect 12796 37324 13020 37380
rect 12460 35868 12628 35924
rect 12684 35924 12740 35934
rect 12460 35476 12516 35868
rect 12684 35830 12740 35868
rect 12572 35700 12628 35710
rect 12572 35606 12628 35644
rect 12796 35698 12852 35710
rect 12796 35646 12798 35698
rect 12850 35646 12852 35698
rect 12796 35476 12852 35646
rect 12460 35420 12740 35476
rect 12012 34738 12068 34748
rect 12124 34860 12292 34916
rect 12572 34916 12628 34926
rect 11676 34626 11732 34636
rect 11676 34244 11732 34254
rect 11676 34150 11732 34188
rect 11340 33292 11620 33348
rect 11676 33348 11732 33358
rect 11340 32900 11396 33292
rect 11676 33254 11732 33292
rect 12012 33348 12068 33358
rect 12012 33254 12068 33292
rect 11452 33124 11508 33134
rect 11452 33030 11508 33068
rect 11564 33122 11620 33134
rect 11564 33070 11566 33122
rect 11618 33070 11620 33122
rect 11340 32844 11508 32900
rect 11228 32722 11284 32732
rect 11340 32564 11396 32574
rect 11116 32562 11396 32564
rect 11116 32510 11342 32562
rect 11394 32510 11396 32562
rect 11116 32508 11396 32510
rect 11340 32498 11396 32508
rect 11340 31892 11396 31902
rect 11340 31554 11396 31836
rect 11340 31502 11342 31554
rect 11394 31502 11396 31554
rect 11340 31332 11396 31502
rect 11340 31266 11396 31276
rect 11452 30772 11508 32844
rect 11564 31556 11620 33070
rect 11900 32788 11956 32798
rect 11900 32694 11956 32732
rect 11788 32004 11844 32014
rect 11788 31910 11844 31948
rect 11564 31490 11620 31500
rect 11676 31666 11732 31678
rect 11676 31614 11678 31666
rect 11730 31614 11732 31666
rect 11564 30772 11620 30782
rect 11452 30716 11564 30772
rect 11564 30706 11620 30716
rect 11676 30212 11732 31614
rect 11900 31668 11956 31678
rect 11900 31666 12068 31668
rect 11900 31614 11902 31666
rect 11954 31614 12068 31666
rect 11900 31612 12068 31614
rect 11900 31602 11956 31612
rect 11004 30034 11060 30044
rect 11116 30156 11732 30212
rect 11004 29092 11060 29102
rect 11004 27860 11060 29036
rect 11116 28532 11172 30156
rect 11900 30098 11956 30110
rect 11900 30046 11902 30098
rect 11954 30046 11956 30098
rect 11228 29986 11284 29998
rect 11228 29934 11230 29986
rect 11282 29934 11284 29986
rect 11228 28868 11284 29934
rect 11900 29876 11956 30046
rect 11900 29810 11956 29820
rect 11228 28802 11284 28812
rect 11340 29764 11396 29774
rect 11116 28466 11172 28476
rect 11340 28196 11396 29708
rect 11788 29652 11844 29662
rect 11788 29558 11844 29596
rect 12012 29316 12068 31612
rect 12124 31108 12180 34860
rect 12572 34802 12628 34860
rect 12572 34750 12574 34802
rect 12626 34750 12628 34802
rect 12572 34738 12628 34750
rect 12236 34690 12292 34702
rect 12236 34638 12238 34690
rect 12290 34638 12292 34690
rect 12236 33684 12292 34638
rect 12348 34356 12404 34366
rect 12348 34262 12404 34300
rect 12684 34244 12740 35420
rect 12796 35410 12852 35420
rect 12684 34188 12964 34244
rect 12236 33618 12292 33628
rect 12684 34018 12740 34030
rect 12684 33966 12686 34018
rect 12738 33966 12740 34018
rect 12572 33236 12628 33246
rect 12236 33234 12628 33236
rect 12236 33182 12574 33234
rect 12626 33182 12628 33234
rect 12236 33180 12628 33182
rect 12236 32004 12292 33180
rect 12572 33170 12628 33180
rect 12684 32564 12740 33966
rect 12908 33570 12964 34188
rect 12908 33518 12910 33570
rect 12962 33518 12964 33570
rect 12908 33506 12964 33518
rect 12684 32498 12740 32508
rect 12908 33346 12964 33358
rect 12908 33294 12910 33346
rect 12962 33294 12964 33346
rect 12572 32452 12628 32462
rect 12572 32358 12628 32396
rect 12236 32002 12740 32004
rect 12236 31950 12238 32002
rect 12290 31950 12740 32002
rect 12236 31948 12740 31950
rect 12236 31938 12292 31948
rect 12460 31780 12516 31790
rect 12460 31686 12516 31724
rect 12124 31042 12180 31052
rect 12460 30882 12516 30894
rect 12460 30830 12462 30882
rect 12514 30830 12516 30882
rect 12236 30660 12292 30670
rect 11900 29260 12068 29316
rect 12124 30210 12180 30222
rect 12124 30158 12126 30210
rect 12178 30158 12180 30210
rect 11676 28868 11732 28878
rect 11676 28642 11732 28812
rect 11676 28590 11678 28642
rect 11730 28590 11732 28642
rect 11676 28578 11732 28590
rect 11228 28084 11284 28094
rect 11228 27990 11284 28028
rect 11340 27970 11396 28140
rect 11340 27918 11342 27970
rect 11394 27918 11396 27970
rect 11340 27906 11396 27918
rect 11788 27972 11844 27982
rect 11004 27858 11284 27860
rect 11004 27806 11006 27858
rect 11058 27806 11284 27858
rect 11004 27804 11284 27806
rect 11004 27794 11060 27804
rect 11228 27748 11284 27804
rect 11228 27692 11732 27748
rect 10892 27580 11060 27636
rect 10444 27022 10446 27074
rect 10498 27022 10500 27074
rect 10444 27010 10500 27022
rect 10892 27074 10948 27086
rect 10892 27022 10894 27074
rect 10946 27022 10948 27074
rect 10556 26402 10612 26414
rect 10556 26350 10558 26402
rect 10610 26350 10612 26402
rect 10556 25956 10612 26350
rect 10556 25890 10612 25900
rect 10668 26068 10724 26078
rect 10556 24276 10612 24286
rect 10556 23938 10612 24220
rect 10556 23886 10558 23938
rect 10610 23886 10612 23938
rect 10556 23874 10612 23886
rect 10668 22932 10724 26012
rect 10780 26066 10836 26078
rect 10780 26014 10782 26066
rect 10834 26014 10836 26066
rect 10780 25732 10836 26014
rect 10780 25666 10836 25676
rect 10892 24388 10948 27022
rect 11004 26908 11060 27580
rect 11340 27524 11396 27534
rect 11004 26852 11284 26908
rect 11116 26516 11172 26526
rect 11228 26516 11284 26852
rect 11116 26514 11284 26516
rect 11116 26462 11118 26514
rect 11170 26462 11284 26514
rect 11116 26460 11284 26462
rect 11116 26450 11172 26460
rect 11340 26404 11396 27468
rect 11228 26348 11396 26404
rect 11228 26292 11284 26348
rect 10780 24332 10948 24388
rect 11004 26236 11284 26292
rect 11564 26292 11620 26302
rect 10780 23492 10836 24332
rect 10892 24164 10948 24174
rect 10892 23826 10948 24108
rect 10892 23774 10894 23826
rect 10946 23774 10948 23826
rect 10892 23762 10948 23774
rect 10780 23426 10836 23436
rect 10668 22876 10836 22932
rect 10668 22370 10724 22382
rect 10668 22318 10670 22370
rect 10722 22318 10724 22370
rect 10332 20974 10334 21026
rect 10386 20974 10388 21026
rect 10332 20962 10388 20974
rect 10444 21924 10500 21934
rect 10220 20914 10276 20926
rect 10220 20862 10222 20914
rect 10274 20862 10276 20914
rect 10220 20580 10276 20862
rect 10220 20514 10276 20524
rect 10444 20020 10500 21868
rect 10668 21588 10724 22318
rect 10780 21812 10836 22876
rect 10780 21718 10836 21756
rect 10892 22708 10948 22718
rect 9996 19628 10164 19684
rect 10220 19964 10500 20020
rect 10556 20580 10612 20590
rect 10556 20018 10612 20524
rect 10556 19966 10558 20018
rect 10610 19966 10612 20018
rect 9996 16882 10052 19628
rect 10220 18452 10276 19964
rect 10556 19796 10612 19966
rect 10220 18386 10276 18396
rect 10444 19740 10612 19796
rect 10444 18228 10500 19740
rect 10668 19236 10724 21532
rect 10668 19170 10724 19180
rect 10780 21252 10836 21262
rect 10780 19012 10836 21196
rect 10220 18172 10500 18228
rect 10556 18956 10836 19012
rect 10892 20018 10948 22652
rect 10892 19966 10894 20018
rect 10946 19966 10948 20018
rect 9996 16830 9998 16882
rect 10050 16830 10052 16882
rect 9996 16818 10052 16830
rect 10108 17556 10164 17566
rect 10108 17332 10164 17500
rect 9884 15314 9940 15596
rect 9884 15262 9886 15314
rect 9938 15262 9940 15314
rect 9884 15250 9940 15262
rect 9660 14478 9662 14530
rect 9714 14478 9716 14530
rect 9100 14354 9156 14364
rect 9100 13972 9156 13982
rect 8092 10834 8260 10836
rect 8092 10782 8094 10834
rect 8146 10782 8260 10834
rect 8092 10780 8260 10782
rect 8428 12460 8820 12516
rect 8876 13858 8932 13870
rect 8876 13806 8878 13858
rect 8930 13806 8932 13858
rect 8092 10770 8148 10780
rect 8092 9940 8148 9950
rect 8148 9884 8260 9940
rect 8092 9874 8148 9884
rect 8204 9826 8260 9884
rect 8204 9774 8206 9826
rect 8258 9774 8260 9826
rect 8204 9762 8260 9774
rect 7532 9154 7700 9156
rect 7532 9102 7534 9154
rect 7586 9102 7700 9154
rect 7532 9100 7700 9102
rect 7756 9436 8036 9492
rect 8316 9602 8372 9614
rect 8316 9550 8318 9602
rect 8370 9550 8372 9602
rect 8316 9492 8372 9550
rect 7532 9090 7588 9100
rect 7756 9044 7812 9436
rect 7644 8988 7812 9044
rect 7980 9044 8036 9054
rect 8204 9044 8260 9054
rect 7420 8930 7476 8942
rect 7420 8878 7422 8930
rect 7474 8878 7476 8930
rect 7420 8820 7476 8878
rect 7420 8754 7476 8764
rect 7420 8484 7476 8494
rect 7308 8482 7476 8484
rect 7308 8430 7422 8482
rect 7474 8430 7476 8482
rect 7308 8428 7476 8430
rect 6860 8418 6916 8428
rect 7420 8418 7476 8428
rect 6636 8204 6804 8260
rect 6860 8260 6916 8270
rect 7308 8260 7364 8270
rect 6860 8258 7364 8260
rect 6860 8206 6862 8258
rect 6914 8206 7310 8258
rect 7362 8206 7364 8258
rect 6860 8204 7364 8206
rect 6636 7812 6692 8204
rect 6860 8194 6916 8204
rect 7308 8194 7364 8204
rect 6748 8036 6804 8046
rect 6972 8036 7028 8046
rect 6748 8034 6916 8036
rect 6748 7982 6750 8034
rect 6802 7982 6916 8034
rect 6748 7980 6916 7982
rect 6748 7970 6804 7980
rect 6636 7756 6804 7812
rect 6524 7746 6580 7756
rect 6636 7588 6692 7598
rect 6300 7586 6692 7588
rect 6300 7534 6638 7586
rect 6690 7534 6692 7586
rect 6300 7532 6692 7534
rect 6300 7362 6356 7532
rect 6636 7522 6692 7532
rect 6300 7310 6302 7362
rect 6354 7310 6356 7362
rect 6300 7298 6356 7310
rect 6748 7252 6804 7756
rect 6860 7700 6916 7980
rect 6860 7634 6916 7644
rect 6972 7698 7028 7980
rect 6972 7646 6974 7698
rect 7026 7646 7028 7698
rect 6972 7634 7028 7646
rect 7532 8036 7588 8046
rect 7532 7700 7588 7980
rect 7644 7924 7700 8988
rect 7868 8932 7924 8942
rect 7868 8838 7924 8876
rect 7980 8708 8036 8988
rect 7980 8642 8036 8652
rect 8092 9042 8260 9044
rect 8092 8990 8206 9042
rect 8258 8990 8260 9042
rect 8092 8988 8260 8990
rect 8092 8484 8148 8988
rect 8204 8978 8260 8988
rect 7980 8428 8148 8484
rect 7980 8258 8036 8428
rect 7980 8206 7982 8258
rect 8034 8206 8036 8258
rect 7756 8036 7812 8046
rect 7868 8036 7924 8046
rect 7756 8034 7868 8036
rect 7756 7982 7758 8034
rect 7810 7982 7868 8034
rect 7756 7980 7868 7982
rect 7756 7970 7812 7980
rect 7644 7858 7700 7868
rect 7532 7644 7812 7700
rect 6972 7476 7028 7486
rect 6972 7382 7028 7420
rect 7308 7474 7364 7486
rect 7308 7422 7310 7474
rect 7362 7422 7364 7474
rect 6748 7196 6916 7252
rect 6748 6804 6804 6814
rect 6748 6690 6804 6748
rect 6748 6638 6750 6690
rect 6802 6638 6804 6690
rect 6076 6402 6132 6412
rect 6188 6466 6244 6478
rect 6188 6414 6190 6466
rect 6242 6414 6244 6466
rect 6188 6132 6244 6414
rect 6188 5572 6244 6076
rect 6300 6466 6356 6478
rect 6300 6414 6302 6466
rect 6354 6414 6356 6466
rect 6300 5796 6356 6414
rect 6412 6468 6468 6478
rect 6468 6412 6692 6468
rect 6412 6374 6468 6412
rect 6300 5730 6356 5740
rect 6188 5516 6468 5572
rect 5852 4562 6020 4564
rect 5852 4510 5854 4562
rect 5906 4510 6020 4562
rect 5852 4508 6020 4510
rect 5852 4498 5908 4508
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 5964 3388 6020 4508
rect 6188 5236 6244 5246
rect 6188 4340 6244 5180
rect 6412 5234 6468 5516
rect 6636 5346 6692 6412
rect 6748 5794 6804 6638
rect 6860 6692 6916 7196
rect 6972 6692 7028 6702
rect 6860 6690 7028 6692
rect 6860 6638 6974 6690
rect 7026 6638 7028 6690
rect 6860 6636 7028 6638
rect 7308 6692 7364 7422
rect 7532 7476 7588 7486
rect 7420 6692 7476 6702
rect 7308 6636 7420 6692
rect 6972 6626 7028 6636
rect 7420 6598 7476 6636
rect 7084 6468 7140 6478
rect 7084 6374 7140 6412
rect 7420 6468 7476 6478
rect 7084 6132 7140 6142
rect 7084 6038 7140 6076
rect 7420 5906 7476 6412
rect 7420 5854 7422 5906
rect 7474 5854 7476 5906
rect 7420 5842 7476 5854
rect 6748 5742 6750 5794
rect 6802 5742 6804 5794
rect 6748 5730 6804 5742
rect 7308 5796 7364 5806
rect 6636 5294 6638 5346
rect 6690 5294 6692 5346
rect 6636 5282 6692 5294
rect 7308 5346 7364 5740
rect 7308 5294 7310 5346
rect 7362 5294 7364 5346
rect 7308 5282 7364 5294
rect 7420 5348 7476 5358
rect 7532 5348 7588 7420
rect 7756 7474 7812 7644
rect 7756 7422 7758 7474
rect 7810 7422 7812 7474
rect 7756 7410 7812 7422
rect 7868 7252 7924 7980
rect 7756 7196 7924 7252
rect 7756 6020 7812 7196
rect 7980 7028 8036 8206
rect 8204 8260 8260 8270
rect 8204 8166 8260 8204
rect 8092 8148 8148 8158
rect 8092 8054 8148 8092
rect 8092 7700 8148 7710
rect 8316 7700 8372 9436
rect 8428 9604 8484 12460
rect 8652 12292 8708 12302
rect 8876 12292 8932 13806
rect 8708 12236 8932 12292
rect 9100 13524 9156 13916
rect 9660 13970 9716 14478
rect 9884 15092 9940 15102
rect 10108 15092 10164 17276
rect 10220 15148 10276 18172
rect 10556 17108 10612 18956
rect 10780 18564 10836 18574
rect 10556 17106 10724 17108
rect 10556 17054 10558 17106
rect 10610 17054 10724 17106
rect 10556 17052 10724 17054
rect 10556 17042 10612 17052
rect 10444 16882 10500 16894
rect 10444 16830 10446 16882
rect 10498 16830 10500 16882
rect 10332 16660 10388 16670
rect 10332 16100 10388 16604
rect 10444 16212 10500 16830
rect 10444 16156 10612 16212
rect 10332 15314 10388 16044
rect 10444 15988 10500 15998
rect 10444 15894 10500 15932
rect 10332 15262 10334 15314
rect 10386 15262 10388 15314
rect 10332 15250 10388 15262
rect 10220 15092 10388 15148
rect 9884 14530 9940 15036
rect 9996 15036 10164 15092
rect 9996 14756 10052 15036
rect 10220 14980 10276 14990
rect 9996 14690 10052 14700
rect 10108 14924 10220 14980
rect 9884 14478 9886 14530
rect 9938 14478 9940 14530
rect 9884 14466 9940 14478
rect 9660 13918 9662 13970
rect 9714 13918 9716 13970
rect 9660 13906 9716 13918
rect 9772 14420 9828 14430
rect 9100 12964 9156 13468
rect 8652 12198 8708 12236
rect 8988 12178 9044 12190
rect 8988 12126 8990 12178
rect 9042 12126 9044 12178
rect 8988 12068 9044 12126
rect 9100 12180 9156 12908
rect 9660 12964 9716 12974
rect 9548 12516 9604 12526
rect 9548 12402 9604 12460
rect 9548 12350 9550 12402
rect 9602 12350 9604 12402
rect 9548 12338 9604 12350
rect 9100 12114 9156 12124
rect 8988 12002 9044 12012
rect 9660 11844 9716 12908
rect 9660 11778 9716 11788
rect 9772 11620 9828 14364
rect 9996 13522 10052 13534
rect 9996 13470 9998 13522
rect 10050 13470 10052 13522
rect 9884 13188 9940 13198
rect 9884 13074 9940 13132
rect 9884 13022 9886 13074
rect 9938 13022 9940 13074
rect 9884 13010 9940 13022
rect 9996 12964 10052 13470
rect 9996 12898 10052 12908
rect 10108 12628 10164 14924
rect 10220 14914 10276 14924
rect 10220 13860 10276 13870
rect 10220 13746 10276 13804
rect 10220 13694 10222 13746
rect 10274 13694 10276 13746
rect 10220 13682 10276 13694
rect 10332 13412 10388 15092
rect 10444 14756 10500 14766
rect 10444 14642 10500 14700
rect 10444 14590 10446 14642
rect 10498 14590 10500 14642
rect 10444 14578 10500 14590
rect 10556 13972 10612 16156
rect 10668 14980 10724 17052
rect 10780 17106 10836 18508
rect 10892 18338 10948 19966
rect 10892 18286 10894 18338
rect 10946 18286 10948 18338
rect 10892 18274 10948 18286
rect 11004 18340 11060 26236
rect 11564 26198 11620 26236
rect 11340 26180 11396 26190
rect 11228 26124 11340 26180
rect 11116 25506 11172 25518
rect 11116 25454 11118 25506
rect 11170 25454 11172 25506
rect 11116 22594 11172 25454
rect 11116 22542 11118 22594
rect 11170 22542 11172 22594
rect 11116 22372 11172 22542
rect 11116 22306 11172 22316
rect 11116 21700 11172 21710
rect 11116 21476 11172 21644
rect 11116 21410 11172 21420
rect 11228 21252 11284 26124
rect 11340 26114 11396 26124
rect 11340 24612 11396 24622
rect 11340 24610 11508 24612
rect 11340 24558 11342 24610
rect 11394 24558 11508 24610
rect 11340 24556 11508 24558
rect 11340 24546 11396 24556
rect 11452 23268 11508 24556
rect 11564 24164 11620 24174
rect 11676 24164 11732 27692
rect 11788 27074 11844 27916
rect 11788 27022 11790 27074
rect 11842 27022 11844 27074
rect 11788 24948 11844 27022
rect 11788 24882 11844 24892
rect 11900 24724 11956 29260
rect 12012 27858 12068 27870
rect 12012 27806 12014 27858
rect 12066 27806 12068 27858
rect 12012 26962 12068 27806
rect 12012 26910 12014 26962
rect 12066 26910 12068 26962
rect 12012 26898 12068 26910
rect 12124 26516 12180 30158
rect 12236 27076 12292 30604
rect 12348 30322 12404 30334
rect 12348 30270 12350 30322
rect 12402 30270 12404 30322
rect 12348 29764 12404 30270
rect 12460 30212 12516 30830
rect 12460 30146 12516 30156
rect 12348 29698 12404 29708
rect 12684 29652 12740 31948
rect 12908 30436 12964 33294
rect 12908 30370 12964 30380
rect 12908 30212 12964 30222
rect 13020 30212 13076 37324
rect 13132 36820 13188 37772
rect 13132 36754 13188 36764
rect 13468 36596 13524 39454
rect 13580 39394 13636 39406
rect 13580 39342 13582 39394
rect 13634 39342 13636 39394
rect 13580 38948 13636 39342
rect 13580 38882 13636 38892
rect 13804 38668 13860 39564
rect 14140 39618 14196 41244
rect 14588 41234 14644 41244
rect 15932 41298 15988 41804
rect 16044 41794 16100 41804
rect 16044 41412 16100 41422
rect 16156 41412 16212 42590
rect 16940 42532 16996 43260
rect 16940 42438 16996 42476
rect 16828 41972 16884 41982
rect 16828 41878 16884 41916
rect 16044 41410 16212 41412
rect 16044 41358 16046 41410
rect 16098 41358 16212 41410
rect 16044 41356 16212 41358
rect 16044 41346 16100 41356
rect 15932 41246 15934 41298
rect 15986 41246 15988 41298
rect 15932 41234 15988 41246
rect 15484 40964 15540 40974
rect 15820 40964 15876 40974
rect 15484 40962 15876 40964
rect 15484 40910 15486 40962
rect 15538 40910 15822 40962
rect 15874 40910 15876 40962
rect 15484 40908 15876 40910
rect 15484 40898 15540 40908
rect 15260 40404 15316 40414
rect 15708 40404 15764 40414
rect 15260 40402 15764 40404
rect 15260 40350 15262 40402
rect 15314 40350 15710 40402
rect 15762 40350 15764 40402
rect 15260 40348 15764 40350
rect 15260 40338 15316 40348
rect 14476 40292 14532 40302
rect 14476 40198 14532 40236
rect 14140 39566 14142 39618
rect 14194 39566 14196 39618
rect 14140 39554 14196 39566
rect 14812 39508 14868 39518
rect 15260 39508 15316 39518
rect 14812 39506 15204 39508
rect 14812 39454 14814 39506
rect 14866 39454 15204 39506
rect 14812 39452 15204 39454
rect 14812 39442 14868 39452
rect 14924 39284 14980 39294
rect 13916 39172 13972 39182
rect 13916 38946 13972 39116
rect 14924 39058 14980 39228
rect 14924 39006 14926 39058
rect 14978 39006 14980 39058
rect 13916 38894 13918 38946
rect 13970 38894 13972 38946
rect 13916 38882 13972 38894
rect 14364 38946 14420 38958
rect 14364 38894 14366 38946
rect 14418 38894 14420 38946
rect 14028 38836 14084 38846
rect 13804 38612 13972 38668
rect 13580 38052 13636 38062
rect 13580 37958 13636 37996
rect 13916 38050 13972 38612
rect 13916 37998 13918 38050
rect 13970 37998 13972 38050
rect 13916 37986 13972 37998
rect 13916 37156 13972 37166
rect 14028 37156 14084 38780
rect 14252 38834 14308 38846
rect 14252 38782 14254 38834
rect 14306 38782 14308 38834
rect 13916 37154 14084 37156
rect 13916 37102 13918 37154
rect 13970 37102 14084 37154
rect 13916 37100 14084 37102
rect 14140 37268 14196 37278
rect 13916 37090 13972 37100
rect 13132 36540 13524 36596
rect 13132 35924 13188 36540
rect 13916 36484 13972 36494
rect 14140 36484 14196 37212
rect 14252 37156 14308 38782
rect 14364 37492 14420 38894
rect 14588 38834 14644 38846
rect 14588 38782 14590 38834
rect 14642 38782 14644 38834
rect 14588 38052 14644 38782
rect 14588 37986 14644 37996
rect 14364 37436 14756 37492
rect 14700 37380 14756 37436
rect 14700 37378 14868 37380
rect 14700 37326 14702 37378
rect 14754 37326 14868 37378
rect 14700 37324 14868 37326
rect 14700 37314 14756 37324
rect 14364 37156 14420 37166
rect 14252 37154 14420 37156
rect 14252 37102 14366 37154
rect 14418 37102 14420 37154
rect 14252 37100 14420 37102
rect 14364 36708 14420 37100
rect 14364 36642 14420 36652
rect 14700 36708 14756 36718
rect 13916 36482 14196 36484
rect 13916 36430 13918 36482
rect 13970 36430 14142 36482
rect 14194 36430 14196 36482
rect 13916 36428 14196 36430
rect 13916 36418 13972 36428
rect 14140 36418 14196 36428
rect 13580 36370 13636 36382
rect 13580 36318 13582 36370
rect 13634 36318 13636 36370
rect 13132 35698 13188 35868
rect 13132 35646 13134 35698
rect 13186 35646 13188 35698
rect 13132 35634 13188 35646
rect 13244 36148 13300 36158
rect 13244 35140 13300 36092
rect 13468 35588 13524 35598
rect 13244 35074 13300 35084
rect 13356 35474 13412 35486
rect 13356 35422 13358 35474
rect 13410 35422 13412 35474
rect 13356 35138 13412 35422
rect 13356 35086 13358 35138
rect 13410 35086 13412 35138
rect 13356 35074 13412 35086
rect 13244 34130 13300 34142
rect 13244 34078 13246 34130
rect 13298 34078 13300 34130
rect 13244 31892 13300 34078
rect 13244 31826 13300 31836
rect 12908 30210 13076 30212
rect 12908 30158 12910 30210
rect 12962 30158 13076 30210
rect 12908 30156 13076 30158
rect 13132 31668 13188 31678
rect 12908 29876 12964 30156
rect 12348 29428 12404 29438
rect 12348 29334 12404 29372
rect 12684 29426 12740 29596
rect 12684 29374 12686 29426
rect 12738 29374 12740 29426
rect 12572 27860 12628 27870
rect 12684 27860 12740 29374
rect 12572 27858 12740 27860
rect 12572 27806 12574 27858
rect 12626 27806 12740 27858
rect 12572 27804 12740 27806
rect 12796 29820 12964 29876
rect 12572 27794 12628 27804
rect 12796 27636 12852 29820
rect 12908 29652 12964 29662
rect 12908 28866 12964 29596
rect 12908 28814 12910 28866
rect 12962 28814 12964 28866
rect 12908 28802 12964 28814
rect 12908 28196 12964 28206
rect 12908 27860 12964 28140
rect 12908 27858 13076 27860
rect 12908 27806 12910 27858
rect 12962 27806 13076 27858
rect 12908 27804 13076 27806
rect 12908 27794 12964 27804
rect 12796 27580 12964 27636
rect 12684 27188 12740 27198
rect 12348 27076 12404 27086
rect 12292 27074 12404 27076
rect 12292 27022 12350 27074
rect 12402 27022 12404 27074
rect 12292 27020 12404 27022
rect 12236 26982 12292 27020
rect 12348 27010 12404 27020
rect 12684 27074 12740 27132
rect 12684 27022 12686 27074
rect 12738 27022 12740 27074
rect 12684 27010 12740 27022
rect 12796 26964 12852 27002
rect 12796 26898 12852 26908
rect 12908 26908 12964 27580
rect 13020 27412 13076 27804
rect 13132 27746 13188 31612
rect 13468 31668 13524 35532
rect 13580 35364 13636 36318
rect 13692 36260 13748 36270
rect 14252 36260 14308 36270
rect 13692 36258 13860 36260
rect 13692 36206 13694 36258
rect 13746 36206 13860 36258
rect 13692 36204 13860 36206
rect 13692 36194 13748 36204
rect 13692 35924 13748 35934
rect 13692 35830 13748 35868
rect 13580 35298 13636 35308
rect 13804 35252 13860 36204
rect 14140 36258 14308 36260
rect 14140 36206 14254 36258
rect 14306 36206 14308 36258
rect 14140 36204 14308 36206
rect 14028 35812 14084 35822
rect 14028 35718 14084 35756
rect 13804 35186 13860 35196
rect 14028 35476 14084 35486
rect 13804 34914 13860 34926
rect 13804 34862 13806 34914
rect 13858 34862 13860 34914
rect 13804 34804 13860 34862
rect 13804 34738 13860 34748
rect 13916 34916 13972 34926
rect 13580 34130 13636 34142
rect 13580 34078 13582 34130
rect 13634 34078 13636 34130
rect 13580 33908 13636 34078
rect 13916 34130 13972 34860
rect 13916 34078 13918 34130
rect 13970 34078 13972 34130
rect 13916 34066 13972 34078
rect 14028 34914 14084 35420
rect 14140 35140 14196 36204
rect 14252 36194 14308 36204
rect 14476 36260 14532 36270
rect 14476 36258 14644 36260
rect 14476 36206 14478 36258
rect 14530 36206 14644 36258
rect 14476 36204 14644 36206
rect 14476 36194 14532 36204
rect 14476 36036 14532 36046
rect 14140 35074 14196 35084
rect 14252 35700 14308 35710
rect 14252 35026 14308 35644
rect 14364 35698 14420 35710
rect 14364 35646 14366 35698
rect 14418 35646 14420 35698
rect 14364 35588 14420 35646
rect 14364 35522 14420 35532
rect 14252 34974 14254 35026
rect 14306 34974 14308 35026
rect 14252 34962 14308 34974
rect 14364 35252 14420 35262
rect 14028 34862 14030 34914
rect 14082 34862 14084 34914
rect 13580 33842 13636 33852
rect 14028 33908 14084 34862
rect 14364 34356 14420 35196
rect 14364 34290 14420 34300
rect 14364 34132 14420 34142
rect 14364 34038 14420 34076
rect 14028 33842 14084 33852
rect 14252 33684 14308 33694
rect 14028 33572 14084 33582
rect 13468 31602 13524 31612
rect 13580 33460 13636 33470
rect 13580 33236 13636 33404
rect 13244 31108 13300 31118
rect 13244 30882 13300 31052
rect 13244 30830 13246 30882
rect 13298 30830 13300 30882
rect 13244 30818 13300 30830
rect 13468 30436 13524 30446
rect 13244 29876 13300 29886
rect 13300 29820 13412 29876
rect 13244 29810 13300 29820
rect 13356 29316 13412 29820
rect 13132 27694 13134 27746
rect 13186 27694 13188 27746
rect 13132 27682 13188 27694
rect 13244 29260 13412 29316
rect 13020 27346 13076 27356
rect 13020 27076 13076 27114
rect 13020 27010 13076 27020
rect 12908 26852 13076 26908
rect 12012 26460 12180 26516
rect 12012 26180 12068 26460
rect 12012 26114 12068 26124
rect 12124 26290 12180 26302
rect 12124 26238 12126 26290
rect 12178 26238 12180 26290
rect 11900 24668 12068 24724
rect 11564 24162 11732 24164
rect 11564 24110 11566 24162
rect 11618 24110 11732 24162
rect 11564 24108 11732 24110
rect 11564 24098 11620 24108
rect 12012 24052 12068 24668
rect 12124 24500 12180 26238
rect 12348 26292 12404 26302
rect 12236 25394 12292 25406
rect 12236 25342 12238 25394
rect 12290 25342 12292 25394
rect 12236 24724 12292 25342
rect 12236 24658 12292 24668
rect 12124 24444 12292 24500
rect 12012 23958 12068 23996
rect 11676 23938 11732 23950
rect 11900 23940 11956 23950
rect 11676 23886 11678 23938
rect 11730 23886 11732 23938
rect 11676 23492 11732 23886
rect 11564 23268 11620 23278
rect 11452 23212 11564 23268
rect 11564 21588 11620 23212
rect 11676 23044 11732 23436
rect 11676 22978 11732 22988
rect 11788 23884 11900 23940
rect 11676 22370 11732 22382
rect 11676 22318 11678 22370
rect 11730 22318 11732 22370
rect 11676 21812 11732 22318
rect 11676 21746 11732 21756
rect 11676 21588 11732 21598
rect 11564 21586 11732 21588
rect 11564 21534 11678 21586
rect 11730 21534 11732 21586
rect 11564 21532 11732 21534
rect 11116 21196 11284 21252
rect 11116 20130 11172 21196
rect 11676 20692 11732 21532
rect 11676 20626 11732 20636
rect 11116 20078 11118 20130
rect 11170 20078 11172 20130
rect 11116 20066 11172 20078
rect 11564 20132 11620 20142
rect 11788 20132 11844 23884
rect 11900 23874 11956 23884
rect 12124 23828 12180 23838
rect 12012 23772 12124 23828
rect 12012 23268 12068 23772
rect 12124 23762 12180 23772
rect 12124 23492 12180 23502
rect 12236 23492 12292 24444
rect 12180 23436 12292 23492
rect 12124 23426 12180 23436
rect 12348 23378 12404 26236
rect 12460 26180 12516 26190
rect 12460 26086 12516 26124
rect 13020 25956 13076 26852
rect 12348 23326 12350 23378
rect 12402 23326 12404 23378
rect 12348 23314 12404 23326
rect 12460 25900 13076 25956
rect 12460 23938 12516 25900
rect 12796 25732 12852 25742
rect 12796 25638 12852 25676
rect 12572 25620 12628 25630
rect 12572 24836 12628 25564
rect 12908 25508 12964 25518
rect 12908 25506 13188 25508
rect 12908 25454 12910 25506
rect 12962 25454 13188 25506
rect 12908 25452 13188 25454
rect 12908 25442 12964 25452
rect 13020 24948 13076 24958
rect 12572 24834 12852 24836
rect 12572 24782 12574 24834
rect 12626 24782 12852 24834
rect 12572 24780 12852 24782
rect 12572 24770 12628 24780
rect 12460 23886 12462 23938
rect 12514 23886 12516 23938
rect 11900 23212 12068 23268
rect 12236 23268 12292 23278
rect 11900 20690 11956 23212
rect 12236 23154 12292 23212
rect 12236 23102 12238 23154
rect 12290 23102 12292 23154
rect 12236 23090 12292 23102
rect 12012 23042 12068 23054
rect 12012 22990 12014 23042
rect 12066 22990 12068 23042
rect 12012 22932 12068 22990
rect 12068 22876 12292 22932
rect 12012 22866 12068 22876
rect 11900 20638 11902 20690
rect 11954 20638 11956 20690
rect 11900 20468 11956 20638
rect 11900 20402 11956 20412
rect 12012 21588 12068 21598
rect 11900 20132 11956 20142
rect 11788 20130 11956 20132
rect 11788 20078 11902 20130
rect 11954 20078 11956 20130
rect 11788 20076 11956 20078
rect 11564 20038 11620 20076
rect 11900 20066 11956 20076
rect 11228 20020 11284 20030
rect 12012 20020 12068 21532
rect 12236 21588 12292 22876
rect 12348 22148 12404 22158
rect 12348 22054 12404 22092
rect 12236 20692 12292 21532
rect 12348 20692 12404 20702
rect 12236 20690 12404 20692
rect 12236 20638 12350 20690
rect 12402 20638 12404 20690
rect 12236 20636 12404 20638
rect 12348 20626 12404 20636
rect 12460 20468 12516 23886
rect 12796 23266 12852 24780
rect 13020 23716 13076 24892
rect 13020 23650 13076 23660
rect 13132 24722 13188 25452
rect 13132 24670 13134 24722
rect 13186 24670 13188 24722
rect 12796 23214 12798 23266
rect 12850 23214 12852 23266
rect 12796 22708 12852 23214
rect 12796 22642 12852 22652
rect 12908 22596 12964 22606
rect 12908 22482 12964 22540
rect 12908 22430 12910 22482
rect 12962 22430 12964 22482
rect 12908 22418 12964 22430
rect 12908 22036 12964 22046
rect 12796 21474 12852 21486
rect 12796 21422 12798 21474
rect 12850 21422 12852 21474
rect 12572 20804 12628 20814
rect 12572 20692 12628 20748
rect 12572 20636 12740 20692
rect 12236 20412 12516 20468
rect 12124 20020 12180 20030
rect 12012 20018 12180 20020
rect 12012 19966 12126 20018
rect 12178 19966 12180 20018
rect 12012 19964 12180 19966
rect 11228 19346 11284 19964
rect 12124 19954 12180 19964
rect 11228 19294 11230 19346
rect 11282 19294 11284 19346
rect 11228 19282 11284 19294
rect 11004 17780 11060 18284
rect 11228 19124 11284 19134
rect 11116 17780 11172 17790
rect 11004 17778 11172 17780
rect 11004 17726 11118 17778
rect 11170 17726 11172 17778
rect 11004 17724 11172 17726
rect 11116 17714 11172 17724
rect 10780 17054 10782 17106
rect 10834 17054 10836 17106
rect 10780 17042 10836 17054
rect 11228 16884 11284 19068
rect 11452 19124 11508 19134
rect 11452 18564 11508 19068
rect 11452 18498 11508 18508
rect 11676 19122 11732 19134
rect 11676 19070 11678 19122
rect 11730 19070 11732 19122
rect 11004 16772 11060 16782
rect 10668 14914 10724 14924
rect 10892 16770 11060 16772
rect 10892 16718 11006 16770
rect 11058 16718 11060 16770
rect 10892 16716 11060 16718
rect 10892 14756 10948 16716
rect 11004 16706 11060 16716
rect 11228 16100 11284 16828
rect 11116 16098 11284 16100
rect 11116 16046 11230 16098
rect 11282 16046 11284 16098
rect 11116 16044 11284 16046
rect 11116 15148 11172 16044
rect 11228 16034 11284 16044
rect 11340 18340 11396 18350
rect 10892 14690 10948 14700
rect 11004 15092 11172 15148
rect 11228 15202 11284 15214
rect 11228 15150 11230 15202
rect 11282 15150 11284 15202
rect 10780 14306 10836 14318
rect 10780 14254 10782 14306
rect 10834 14254 10836 14306
rect 10780 13972 10836 14254
rect 9996 12572 10164 12628
rect 10220 13356 10388 13412
rect 10444 13916 10836 13972
rect 9884 12178 9940 12190
rect 9884 12126 9886 12178
rect 9938 12126 9940 12178
rect 9884 12068 9940 12126
rect 9996 12068 10052 12572
rect 10108 12404 10164 12414
rect 10220 12404 10276 13356
rect 10332 12964 10388 12974
rect 10332 12870 10388 12908
rect 10332 12404 10388 12414
rect 10220 12402 10388 12404
rect 10220 12350 10334 12402
rect 10386 12350 10388 12402
rect 10220 12348 10388 12350
rect 10108 12290 10164 12348
rect 10332 12338 10388 12348
rect 10108 12238 10110 12290
rect 10162 12238 10164 12290
rect 10108 12226 10164 12238
rect 10444 12292 10500 13916
rect 10668 13748 10724 13758
rect 10556 13188 10612 13198
rect 10556 12962 10612 13132
rect 10668 13076 10724 13692
rect 10668 13010 10724 13020
rect 10892 13636 10948 13646
rect 10556 12910 10558 12962
rect 10610 12910 10612 12962
rect 10556 12898 10612 12910
rect 10780 12962 10836 12974
rect 10780 12910 10782 12962
rect 10834 12910 10836 12962
rect 10668 12852 10724 12862
rect 10556 12740 10612 12750
rect 10556 12646 10612 12684
rect 10668 12402 10724 12796
rect 10668 12350 10670 12402
rect 10722 12350 10724 12402
rect 10668 12338 10724 12350
rect 10556 12292 10612 12302
rect 10444 12236 10556 12292
rect 10220 12180 10276 12190
rect 10276 12124 10388 12180
rect 10220 12114 10276 12124
rect 9996 12012 10164 12068
rect 9884 12002 9940 12012
rect 8540 11564 9604 11620
rect 9772 11564 10052 11620
rect 8540 11282 8596 11564
rect 8988 11396 9044 11406
rect 9436 11396 9492 11406
rect 9044 11394 9492 11396
rect 9044 11342 9438 11394
rect 9490 11342 9492 11394
rect 9044 11340 9492 11342
rect 8988 11302 9044 11340
rect 9436 11330 9492 11340
rect 9548 11396 9604 11564
rect 9660 11396 9716 11406
rect 9884 11396 9940 11406
rect 9548 11394 9716 11396
rect 9548 11342 9662 11394
rect 9714 11342 9716 11394
rect 9548 11340 9716 11342
rect 8540 11230 8542 11282
rect 8594 11230 8596 11282
rect 8540 9826 8596 11230
rect 8652 11284 8708 11294
rect 8652 10834 8708 11228
rect 8652 10782 8654 10834
rect 8706 10782 8708 10834
rect 8652 10770 8708 10782
rect 8764 11170 8820 11182
rect 8764 11118 8766 11170
rect 8818 11118 8820 11170
rect 8764 10052 8820 11118
rect 8876 11172 8932 11182
rect 8876 11078 8932 11116
rect 9100 10500 9156 10510
rect 9100 10406 9156 10444
rect 8540 9774 8542 9826
rect 8594 9774 8596 9826
rect 8540 9762 8596 9774
rect 8652 9996 8764 10052
rect 8428 9380 8484 9548
rect 8428 9324 8596 9380
rect 8428 9154 8484 9166
rect 8428 9102 8430 9154
rect 8482 9102 8484 9154
rect 8428 8036 8484 9102
rect 8428 7970 8484 7980
rect 8092 7698 8372 7700
rect 8092 7646 8094 7698
rect 8146 7646 8372 7698
rect 8092 7644 8372 7646
rect 8540 7700 8596 9324
rect 8652 8370 8708 9996
rect 8764 9986 8820 9996
rect 9324 9828 9380 9838
rect 9548 9828 9604 11340
rect 9660 11330 9716 11340
rect 9772 11394 9940 11396
rect 9772 11342 9886 11394
rect 9938 11342 9940 11394
rect 9772 11340 9940 11342
rect 9772 10498 9828 11340
rect 9884 11330 9940 11340
rect 9772 10446 9774 10498
rect 9826 10446 9828 10498
rect 9772 10052 9828 10446
rect 9772 9986 9828 9996
rect 9324 9826 9604 9828
rect 9324 9774 9326 9826
rect 9378 9774 9604 9826
rect 9324 9772 9604 9774
rect 9324 9762 9380 9772
rect 9660 9716 9716 9726
rect 9996 9716 10052 11564
rect 10108 10164 10164 12012
rect 10332 11956 10388 12124
rect 10444 12178 10500 12236
rect 10444 12126 10446 12178
rect 10498 12126 10500 12178
rect 10444 12114 10500 12126
rect 10556 11956 10612 12236
rect 10780 12180 10836 12910
rect 10892 12402 10948 13580
rect 10892 12350 10894 12402
rect 10946 12350 10948 12402
rect 10892 12338 10948 12350
rect 11004 12404 11060 15092
rect 11228 14644 11284 15150
rect 11228 14578 11284 14588
rect 11116 14532 11172 14542
rect 11116 14438 11172 14476
rect 11340 13860 11396 18284
rect 11676 17780 11732 19070
rect 11788 19010 11844 19022
rect 11788 18958 11790 19010
rect 11842 18958 11844 19010
rect 11788 18452 11844 18958
rect 11788 18386 11844 18396
rect 12124 19010 12180 19022
rect 12124 18958 12126 19010
rect 12178 18958 12180 19010
rect 11676 17714 11732 17724
rect 11788 17668 11844 17678
rect 11788 17556 11844 17612
rect 11788 17554 12068 17556
rect 11788 17502 11790 17554
rect 11842 17502 12068 17554
rect 11788 17500 12068 17502
rect 11788 17490 11844 17500
rect 11452 17442 11508 17454
rect 11452 17390 11454 17442
rect 11506 17390 11508 17442
rect 11452 17108 11508 17390
rect 11452 17042 11508 17052
rect 11900 16100 11956 16110
rect 11900 16006 11956 16044
rect 11452 15316 11508 15326
rect 11452 15314 11620 15316
rect 11452 15262 11454 15314
rect 11506 15262 11620 15314
rect 11452 15260 11620 15262
rect 11452 15250 11508 15260
rect 11564 15148 11620 15260
rect 11228 13804 11396 13860
rect 11452 15092 11620 15148
rect 11788 15204 11844 15242
rect 11788 15138 11844 15148
rect 12012 15148 12068 17500
rect 12124 17444 12180 18958
rect 12236 17892 12292 20412
rect 12460 19124 12516 19134
rect 12460 19030 12516 19068
rect 12572 19122 12628 19134
rect 12572 19070 12574 19122
rect 12626 19070 12628 19122
rect 12348 19010 12404 19022
rect 12348 18958 12350 19010
rect 12402 18958 12404 19010
rect 12348 18900 12404 18958
rect 12348 18834 12404 18844
rect 12572 18676 12628 19070
rect 12236 17826 12292 17836
rect 12348 18620 12628 18676
rect 12348 17780 12404 18620
rect 12572 18450 12628 18462
rect 12572 18398 12574 18450
rect 12626 18398 12628 18450
rect 12572 18228 12628 18398
rect 12572 18162 12628 18172
rect 12348 17724 12628 17780
rect 12460 17554 12516 17566
rect 12460 17502 12462 17554
rect 12514 17502 12516 17554
rect 12180 17388 12292 17444
rect 12124 17350 12180 17388
rect 12236 15538 12292 17388
rect 12348 17442 12404 17454
rect 12348 17390 12350 17442
rect 12402 17390 12404 17442
rect 12348 15876 12404 17390
rect 12460 16324 12516 17502
rect 12572 17556 12628 17724
rect 12572 17462 12628 17500
rect 12460 16258 12516 16268
rect 12684 16322 12740 20636
rect 12796 19124 12852 21422
rect 12908 20804 12964 21980
rect 13020 21252 13076 21262
rect 13020 20914 13076 21196
rect 13020 20862 13022 20914
rect 13074 20862 13076 20914
rect 13020 20850 13076 20862
rect 12908 20710 12964 20748
rect 13132 20580 13188 24670
rect 13244 21700 13300 29260
rect 13356 27412 13412 27422
rect 13356 26404 13412 27356
rect 13468 26908 13524 30380
rect 13580 30322 13636 33180
rect 14028 33458 14084 33516
rect 14028 33406 14030 33458
rect 14082 33406 14084 33458
rect 13692 33124 13748 33134
rect 13692 33030 13748 33068
rect 14028 32900 14084 33406
rect 14252 33346 14308 33628
rect 14252 33294 14254 33346
rect 14306 33294 14308 33346
rect 14252 33282 14308 33294
rect 14476 33124 14532 35980
rect 14588 34468 14644 36204
rect 14700 34916 14756 36652
rect 14812 36484 14868 37324
rect 14812 36418 14868 36428
rect 14812 35140 14868 35150
rect 14812 35046 14868 35084
rect 14700 34850 14756 34860
rect 14588 34412 14868 34468
rect 14812 34130 14868 34412
rect 14812 34078 14814 34130
rect 14866 34078 14868 34130
rect 14812 34066 14868 34078
rect 14924 33460 14980 39006
rect 15036 38948 15092 38958
rect 15036 38162 15092 38892
rect 15148 38724 15204 39452
rect 15260 38948 15316 39452
rect 15596 39396 15652 39406
rect 15260 38882 15316 38892
rect 15372 38948 15428 38958
rect 15484 38948 15540 38958
rect 15372 38946 15484 38948
rect 15372 38894 15374 38946
rect 15426 38894 15484 38946
rect 15372 38892 15484 38894
rect 15372 38882 15428 38892
rect 15260 38724 15316 38734
rect 15148 38722 15316 38724
rect 15148 38670 15262 38722
rect 15314 38670 15316 38722
rect 15148 38668 15316 38670
rect 15260 38658 15316 38668
rect 15036 38110 15038 38162
rect 15090 38110 15092 38162
rect 15036 38098 15092 38110
rect 15372 38052 15428 38062
rect 15372 37958 15428 37996
rect 15036 37044 15092 37054
rect 15036 36706 15092 36988
rect 15036 36654 15038 36706
rect 15090 36654 15092 36706
rect 15036 36642 15092 36654
rect 15372 36594 15428 36606
rect 15372 36542 15374 36594
rect 15426 36542 15428 36594
rect 15036 36484 15092 36494
rect 15372 36484 15428 36542
rect 15092 36428 15428 36484
rect 15036 36390 15092 36428
rect 15148 36148 15204 36158
rect 15148 35922 15204 36092
rect 15484 36148 15540 38892
rect 15596 38946 15652 39340
rect 15596 38894 15598 38946
rect 15650 38894 15652 38946
rect 15596 38882 15652 38894
rect 15596 38162 15652 38174
rect 15596 38110 15598 38162
rect 15650 38110 15652 38162
rect 15596 37940 15652 38110
rect 15596 37874 15652 37884
rect 15708 37828 15764 40348
rect 15820 40180 15876 40908
rect 16828 40740 16884 40750
rect 17276 40740 17332 44156
rect 17500 44146 17556 44156
rect 17612 44100 17668 44110
rect 17500 43540 17556 43550
rect 17612 43540 17668 44044
rect 17500 43538 17668 43540
rect 17500 43486 17502 43538
rect 17554 43486 17668 43538
rect 17500 43484 17668 43486
rect 17500 43474 17556 43484
rect 17388 42642 17444 42654
rect 17388 42590 17390 42642
rect 17442 42590 17444 42642
rect 17388 41860 17444 42590
rect 17500 42532 17556 42542
rect 17500 42438 17556 42476
rect 17388 41794 17444 41804
rect 17500 41972 17556 41982
rect 17612 41972 17668 43484
rect 17724 42756 17780 44492
rect 17836 42980 17892 45948
rect 19740 45892 19796 45902
rect 21084 45892 21140 45902
rect 19628 45890 19796 45892
rect 19628 45838 19742 45890
rect 19794 45838 19796 45890
rect 19628 45836 19796 45838
rect 17948 45106 18004 45118
rect 17948 45054 17950 45106
rect 18002 45054 18004 45106
rect 17948 44100 18004 45054
rect 18620 44996 18676 45006
rect 18620 44902 18676 44940
rect 19628 44434 19684 45836
rect 19740 45826 19796 45836
rect 20748 45890 21140 45892
rect 20748 45838 21086 45890
rect 21138 45838 21140 45890
rect 20748 45836 21140 45838
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 20748 44994 20804 45836
rect 21084 45826 21140 45836
rect 20748 44942 20750 44994
rect 20802 44942 20804 44994
rect 20748 44930 20804 44942
rect 21084 45106 21140 45118
rect 21084 45054 21086 45106
rect 21138 45054 21140 45106
rect 19628 44382 19630 44434
rect 19682 44382 19684 44434
rect 19628 44370 19684 44382
rect 17948 44034 18004 44044
rect 20076 44100 20132 44138
rect 20076 44034 20132 44044
rect 20524 44100 20580 44110
rect 20524 44006 20580 44044
rect 21084 44100 21140 45054
rect 21308 44996 21364 45006
rect 21308 44546 21364 44940
rect 21868 44996 21924 45006
rect 21868 44902 21924 44940
rect 21308 44494 21310 44546
rect 21362 44494 21364 44546
rect 21308 44482 21364 44494
rect 21084 44034 21140 44044
rect 21420 44210 21476 44222
rect 21420 44158 21422 44210
rect 21474 44158 21476 44210
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 20972 43652 21028 43662
rect 20972 43650 21364 43652
rect 20972 43598 20974 43650
rect 21026 43598 21364 43650
rect 20972 43596 21364 43598
rect 20972 43586 21028 43596
rect 18172 43428 18228 43438
rect 18172 43334 18228 43372
rect 20300 43426 20356 43438
rect 20300 43374 20302 43426
rect 20354 43374 20356 43426
rect 17948 42980 18004 42990
rect 17836 42924 17948 42980
rect 17948 42914 18004 42924
rect 18956 42980 19012 42990
rect 18956 42886 19012 42924
rect 17948 42756 18004 42766
rect 17724 42754 18004 42756
rect 17724 42702 17950 42754
rect 18002 42702 18004 42754
rect 17724 42700 18004 42702
rect 17948 42690 18004 42700
rect 20300 42756 20356 43374
rect 20860 43428 20916 43438
rect 20860 43334 20916 43372
rect 17724 42532 17780 42542
rect 19180 42532 19236 42542
rect 17724 42530 18004 42532
rect 17724 42478 17726 42530
rect 17778 42478 18004 42530
rect 17724 42476 18004 42478
rect 17724 42466 17780 42476
rect 17556 41916 17668 41972
rect 17948 41970 18004 42476
rect 17948 41918 17950 41970
rect 18002 41918 18004 41970
rect 17500 41858 17556 41916
rect 17948 41906 18004 41918
rect 18396 41972 18452 41982
rect 18396 41878 18452 41916
rect 18620 41972 18676 41982
rect 18620 41970 19012 41972
rect 18620 41918 18622 41970
rect 18674 41918 19012 41970
rect 18620 41916 19012 41918
rect 18620 41906 18676 41916
rect 18172 41860 18228 41870
rect 17500 41806 17502 41858
rect 17554 41806 17556 41858
rect 17500 40964 17556 41806
rect 17500 40898 17556 40908
rect 18060 41858 18228 41860
rect 18060 41806 18174 41858
rect 18226 41806 18228 41858
rect 18060 41804 18228 41806
rect 17276 40684 17780 40740
rect 16716 40514 16772 40526
rect 16716 40462 16718 40514
rect 16770 40462 16772 40514
rect 16604 40402 16660 40414
rect 16604 40350 16606 40402
rect 16658 40350 16660 40402
rect 15820 40114 15876 40124
rect 16268 40290 16324 40302
rect 16268 40238 16270 40290
rect 16322 40238 16324 40290
rect 15932 39060 15988 39070
rect 15932 38966 15988 39004
rect 16044 38836 16100 38846
rect 16044 38742 16100 38780
rect 16268 38388 16324 40238
rect 16604 40068 16660 40350
rect 16604 40002 16660 40012
rect 16716 39732 16772 40462
rect 16828 39956 16884 40684
rect 16940 40628 16996 40638
rect 16940 40626 17668 40628
rect 16940 40574 16942 40626
rect 16994 40574 17668 40626
rect 16940 40572 17668 40574
rect 16940 40562 16996 40572
rect 17612 40514 17668 40572
rect 17724 40626 17780 40684
rect 17724 40574 17726 40626
rect 17778 40574 17780 40626
rect 17724 40562 17780 40574
rect 17612 40462 17614 40514
rect 17666 40462 17668 40514
rect 17612 40450 17668 40462
rect 17500 40402 17556 40414
rect 17500 40350 17502 40402
rect 17554 40350 17556 40402
rect 16828 39900 17332 39956
rect 16940 39732 16996 39742
rect 16716 39730 16996 39732
rect 16716 39678 16942 39730
rect 16994 39678 16996 39730
rect 16716 39676 16996 39678
rect 16380 38948 16436 38958
rect 16380 38834 16436 38892
rect 16380 38782 16382 38834
rect 16434 38782 16436 38834
rect 16380 38770 16436 38782
rect 16940 38836 16996 39676
rect 16940 38770 16996 38780
rect 17276 39732 17332 39900
rect 17276 38834 17332 39676
rect 17388 39396 17444 39406
rect 17388 39302 17444 39340
rect 17500 39060 17556 40350
rect 18060 40402 18116 41804
rect 18172 41794 18228 41804
rect 18956 41412 19012 41916
rect 19068 41860 19124 41870
rect 19068 41766 19124 41804
rect 19068 41412 19124 41422
rect 18956 41410 19124 41412
rect 18956 41358 19070 41410
rect 19122 41358 19124 41410
rect 18956 41356 19124 41358
rect 19068 41346 19124 41356
rect 19180 41074 19236 42476
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19628 42084 19684 42094
rect 20300 42084 20356 42700
rect 19628 42082 20356 42084
rect 19628 42030 19630 42082
rect 19682 42030 20356 42082
rect 19628 42028 20356 42030
rect 21196 43314 21252 43326
rect 21196 43262 21198 43314
rect 21250 43262 21252 43314
rect 21196 42082 21252 43262
rect 21308 42980 21364 43596
rect 21420 43540 21476 44158
rect 23324 44212 23380 44222
rect 23548 44212 23604 46732
rect 25228 46116 25284 46126
rect 25228 46022 25284 46060
rect 24444 45332 24500 45342
rect 23996 45330 24500 45332
rect 23996 45278 24446 45330
rect 24498 45278 24500 45330
rect 23996 45276 24500 45278
rect 23996 44994 24052 45276
rect 24444 45266 24500 45276
rect 26684 45330 26740 49308
rect 27104 49200 27216 50000
rect 28672 49200 28784 50000
rect 30240 49200 30352 50000
rect 31808 49200 31920 50000
rect 33376 49200 33488 50000
rect 34944 49200 35056 50000
rect 36512 49200 36624 50000
rect 38080 49200 38192 50000
rect 39648 49200 39760 50000
rect 41216 49200 41328 50000
rect 42784 49200 42896 50000
rect 44352 49200 44464 50000
rect 45920 49200 46032 50000
rect 27132 47460 27188 49200
rect 27132 47404 27524 47460
rect 27132 45890 27188 45902
rect 27132 45838 27134 45890
rect 27186 45838 27188 45890
rect 27132 45444 27188 45838
rect 27468 45778 27524 47404
rect 27468 45726 27470 45778
rect 27522 45726 27524 45778
rect 27468 45714 27524 45726
rect 28700 45778 28756 49200
rect 30268 46002 30324 49200
rect 30268 45950 30270 46002
rect 30322 45950 30324 46002
rect 30268 45938 30324 45950
rect 28700 45726 28702 45778
rect 28754 45726 28756 45778
rect 28700 45714 28756 45726
rect 31164 45890 31220 45902
rect 31164 45838 31166 45890
rect 31218 45838 31220 45890
rect 27132 45378 27188 45388
rect 26684 45278 26686 45330
rect 26738 45278 26740 45330
rect 26684 45266 26740 45278
rect 30940 45332 30996 45342
rect 30940 45238 30996 45276
rect 25452 45220 25508 45230
rect 25340 45218 25508 45220
rect 25340 45166 25454 45218
rect 25506 45166 25508 45218
rect 25340 45164 25508 45166
rect 24332 45108 24388 45118
rect 24332 45106 24612 45108
rect 24332 45054 24334 45106
rect 24386 45054 24612 45106
rect 24332 45052 24612 45054
rect 24332 45042 24388 45052
rect 23996 44942 23998 44994
rect 24050 44942 24052 44994
rect 23996 44324 24052 44942
rect 24220 44324 24276 44334
rect 23996 44322 24388 44324
rect 23996 44270 24222 44322
rect 24274 44270 24388 44322
rect 23996 44268 24388 44270
rect 24220 44258 24276 44268
rect 23324 44210 23604 44212
rect 23324 44158 23326 44210
rect 23378 44158 23604 44210
rect 23324 44156 23604 44158
rect 23324 44146 23380 44156
rect 21868 44100 21924 44110
rect 21868 44006 21924 44044
rect 22316 44100 22372 44110
rect 22316 44006 22372 44044
rect 22988 44100 23044 44110
rect 22988 44006 23044 44044
rect 21420 43474 21476 43484
rect 22540 43708 22820 43764
rect 21980 43428 22036 43438
rect 22428 43428 22484 43438
rect 21980 43426 22148 43428
rect 21980 43374 21982 43426
rect 22034 43374 22148 43426
rect 21980 43372 22148 43374
rect 21980 43362 22036 43372
rect 21308 42924 21700 42980
rect 21420 42756 21476 42766
rect 21420 42662 21476 42700
rect 21308 42532 21364 42542
rect 21308 42438 21364 42476
rect 21196 42030 21198 42082
rect 21250 42030 21252 42082
rect 19628 42018 19684 42028
rect 21196 42018 21252 42030
rect 21532 42082 21588 42094
rect 21532 42030 21534 42082
rect 21586 42030 21588 42082
rect 20524 41972 20580 41982
rect 20524 41878 20580 41916
rect 21420 41972 21476 41982
rect 19404 41860 19460 41870
rect 19404 41410 19460 41804
rect 19404 41358 19406 41410
rect 19458 41358 19460 41410
rect 19404 41346 19460 41358
rect 21420 41298 21476 41916
rect 21532 41860 21588 42030
rect 21532 41794 21588 41804
rect 21420 41246 21422 41298
rect 21474 41246 21476 41298
rect 21420 41234 21476 41246
rect 19180 41022 19182 41074
rect 19234 41022 19236 41074
rect 19180 41010 19236 41022
rect 18284 40962 18340 40974
rect 18284 40910 18286 40962
rect 18338 40910 18340 40962
rect 18284 40740 18340 40910
rect 18284 40674 18340 40684
rect 18396 40964 18452 40974
rect 18396 40404 18452 40908
rect 20524 40964 20580 40974
rect 20524 40870 20580 40908
rect 21308 40962 21364 40974
rect 21308 40910 21310 40962
rect 21362 40910 21364 40962
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 21308 40628 21364 40910
rect 18060 40350 18062 40402
rect 18114 40350 18116 40402
rect 17948 39620 18004 39630
rect 18060 39620 18116 40350
rect 18284 40402 18452 40404
rect 18284 40350 18398 40402
rect 18450 40350 18452 40402
rect 18284 40348 18452 40350
rect 17948 39618 18116 39620
rect 17948 39566 17950 39618
rect 18002 39566 18116 39618
rect 17948 39564 18116 39566
rect 18172 40068 18228 40078
rect 17948 39554 18004 39564
rect 17836 39060 17892 39070
rect 17500 39058 17892 39060
rect 17500 39006 17838 39058
rect 17890 39006 17892 39058
rect 17500 39004 17892 39006
rect 17836 38994 17892 39004
rect 17948 39060 18004 39070
rect 18172 39060 18228 40012
rect 17948 39058 18228 39060
rect 17948 39006 17950 39058
rect 18002 39006 18228 39058
rect 17948 39004 18228 39006
rect 17948 38994 18004 39004
rect 17276 38782 17278 38834
rect 17330 38782 17332 38834
rect 17276 38668 17332 38782
rect 17724 38836 17780 38846
rect 17724 38742 17780 38780
rect 16268 38322 16324 38332
rect 16380 38610 16436 38622
rect 16716 38612 16772 38622
rect 16380 38558 16382 38610
rect 16434 38558 16436 38610
rect 16268 38162 16324 38174
rect 16268 38110 16270 38162
rect 16322 38110 16324 38162
rect 15708 37762 15764 37772
rect 16156 38050 16212 38062
rect 16156 37998 16158 38050
rect 16210 37998 16212 38050
rect 15484 36082 15540 36092
rect 15932 37268 15988 37278
rect 16156 37268 16212 37998
rect 15932 37266 16212 37268
rect 15932 37214 15934 37266
rect 15986 37214 16212 37266
rect 15932 37212 16212 37214
rect 15148 35870 15150 35922
rect 15202 35870 15204 35922
rect 15148 35858 15204 35870
rect 15708 35812 15764 35822
rect 15708 35810 15876 35812
rect 15708 35758 15710 35810
rect 15762 35758 15876 35810
rect 15708 35756 15876 35758
rect 15708 35746 15764 35756
rect 15260 35586 15316 35598
rect 15260 35534 15262 35586
rect 15314 35534 15316 35586
rect 15036 35364 15092 35374
rect 15036 35028 15092 35308
rect 15148 35028 15204 35038
rect 15036 35026 15204 35028
rect 15036 34974 15150 35026
rect 15202 34974 15204 35026
rect 15036 34972 15204 34974
rect 15148 34962 15204 34972
rect 15260 34580 15316 35534
rect 15372 35476 15428 35486
rect 15372 35474 15652 35476
rect 15372 35422 15374 35474
rect 15426 35422 15652 35474
rect 15372 35420 15652 35422
rect 15372 35410 15428 35420
rect 15260 34514 15316 34524
rect 15372 35028 15428 35038
rect 15372 34802 15428 34972
rect 15372 34750 15374 34802
rect 15426 34750 15428 34802
rect 15036 34468 15092 34478
rect 15036 33684 15092 34412
rect 15148 34244 15204 34254
rect 15148 34130 15204 34188
rect 15148 34078 15150 34130
rect 15202 34078 15204 34130
rect 15148 34066 15204 34078
rect 15036 33618 15092 33628
rect 14028 32834 14084 32844
rect 14140 33068 14532 33124
rect 14812 33404 14980 33460
rect 15372 33460 15428 34750
rect 15596 34244 15652 35420
rect 15820 34860 15876 35756
rect 15932 35026 15988 37212
rect 16268 37156 16324 38110
rect 16268 37090 16324 37100
rect 16380 37044 16436 38558
rect 16492 38610 16772 38612
rect 16492 38558 16718 38610
rect 16770 38558 16772 38610
rect 16492 38556 16772 38558
rect 16492 37378 16548 38556
rect 16716 38546 16772 38556
rect 17164 38612 17332 38668
rect 16492 37326 16494 37378
rect 16546 37326 16548 37378
rect 16492 37314 16548 37326
rect 16604 38388 16660 38398
rect 16380 36978 16436 36988
rect 16492 35810 16548 35822
rect 16492 35758 16494 35810
rect 16546 35758 16548 35810
rect 15932 34974 15934 35026
rect 15986 34974 15988 35026
rect 15932 34962 15988 34974
rect 16044 35698 16100 35710
rect 16044 35646 16046 35698
rect 16098 35646 16100 35698
rect 15708 34802 15764 34814
rect 15820 34804 15988 34860
rect 15708 34750 15710 34802
rect 15762 34750 15764 34802
rect 15708 34468 15764 34750
rect 15708 34412 15876 34468
rect 15708 34244 15764 34254
rect 15596 34242 15764 34244
rect 15596 34190 15710 34242
rect 15762 34190 15764 34242
rect 15596 34188 15764 34190
rect 15708 34178 15764 34188
rect 15820 34244 15876 34412
rect 15820 34178 15876 34188
rect 15484 33460 15540 33470
rect 15372 33458 15540 33460
rect 15372 33406 15486 33458
rect 15538 33406 15540 33458
rect 15372 33404 15540 33406
rect 13804 31890 13860 31902
rect 13804 31838 13806 31890
rect 13858 31838 13860 31890
rect 13692 31778 13748 31790
rect 13692 31726 13694 31778
rect 13746 31726 13748 31778
rect 13692 31668 13748 31726
rect 13692 31602 13748 31612
rect 13692 30772 13748 30782
rect 13804 30772 13860 31838
rect 13748 30716 13860 30772
rect 13692 30706 13748 30716
rect 13580 30270 13582 30322
rect 13634 30270 13636 30322
rect 13580 30258 13636 30270
rect 14140 29988 14196 33068
rect 14476 32562 14532 32574
rect 14476 32510 14478 32562
rect 14530 32510 14532 32562
rect 14476 32340 14532 32510
rect 14476 32274 14532 32284
rect 14476 31892 14532 31902
rect 14140 29894 14196 29932
rect 14252 31780 14308 31790
rect 13916 29764 13972 29774
rect 13580 29540 13636 29550
rect 13636 29484 13748 29540
rect 13580 29446 13636 29484
rect 13580 28756 13636 28766
rect 13580 28662 13636 28700
rect 13692 27860 13748 29484
rect 13916 28642 13972 29708
rect 14252 29428 14308 31724
rect 14476 31108 14532 31836
rect 14588 31780 14644 31790
rect 14588 31686 14644 31724
rect 14476 30210 14532 31052
rect 14476 30158 14478 30210
rect 14530 30158 14532 30210
rect 14476 30146 14532 30158
rect 14812 29876 14868 33404
rect 15484 33394 15540 33404
rect 15932 33348 15988 34804
rect 16044 34468 16100 35646
rect 16044 34402 16100 34412
rect 16156 35364 16212 35374
rect 15708 33292 15988 33348
rect 16044 34132 16100 34142
rect 14924 33236 14980 33246
rect 14924 33142 14980 33180
rect 15372 32788 15428 32798
rect 15036 32732 15372 32788
rect 14924 32340 14980 32350
rect 14924 30996 14980 32284
rect 14924 30930 14980 30940
rect 14924 30100 14980 30110
rect 15036 30100 15092 32732
rect 15372 32694 15428 32732
rect 15260 32564 15316 32574
rect 15260 32470 15316 32508
rect 15596 32562 15652 32574
rect 15596 32510 15598 32562
rect 15650 32510 15652 32562
rect 15596 32340 15652 32510
rect 15596 32274 15652 32284
rect 15596 31668 15652 31678
rect 15260 31554 15316 31566
rect 15260 31502 15262 31554
rect 15314 31502 15316 31554
rect 15260 30436 15316 31502
rect 15372 30996 15428 31006
rect 15372 30902 15428 30940
rect 15260 30370 15316 30380
rect 14924 30098 15092 30100
rect 14924 30046 14926 30098
rect 14978 30046 15092 30098
rect 14924 30044 15092 30046
rect 15148 30324 15204 30334
rect 14924 30034 14980 30044
rect 14812 29810 14868 29820
rect 14364 29428 14420 29438
rect 13916 28590 13918 28642
rect 13970 28590 13972 28642
rect 13916 28578 13972 28590
rect 14028 29426 14420 29428
rect 14028 29374 14366 29426
rect 14418 29374 14420 29426
rect 14028 29372 14420 29374
rect 14028 28420 14084 29372
rect 14364 29362 14420 29372
rect 13804 28364 14084 28420
rect 14364 28642 14420 28654
rect 14364 28590 14366 28642
rect 14418 28590 14420 28642
rect 13804 28082 13860 28364
rect 13804 28030 13806 28082
rect 13858 28030 13860 28082
rect 13804 28018 13860 28030
rect 14252 27972 14308 27982
rect 14252 27878 14308 27916
rect 14140 27860 14196 27870
rect 13692 27804 13860 27860
rect 13580 27524 13636 27534
rect 13580 27186 13636 27468
rect 13580 27134 13582 27186
rect 13634 27134 13636 27186
rect 13580 27122 13636 27134
rect 13692 27074 13748 27086
rect 13692 27022 13694 27074
rect 13746 27022 13748 27074
rect 13468 26852 13636 26908
rect 13356 26338 13412 26348
rect 13580 24500 13636 26852
rect 13692 25620 13748 27022
rect 13692 25554 13748 25564
rect 13692 25396 13748 25406
rect 13692 25302 13748 25340
rect 13804 24836 13860 27804
rect 13916 25844 13972 25854
rect 13916 25730 13972 25788
rect 13916 25678 13918 25730
rect 13970 25678 13972 25730
rect 13916 25666 13972 25678
rect 13804 24770 13860 24780
rect 13468 23940 13524 23950
rect 13468 23846 13524 23884
rect 13580 23826 13636 24444
rect 14028 24724 14084 24734
rect 13580 23774 13582 23826
rect 13634 23774 13636 23826
rect 13580 23762 13636 23774
rect 13804 24276 13860 24286
rect 13468 23716 13524 23726
rect 13468 22370 13524 23660
rect 13468 22318 13470 22370
rect 13522 22318 13524 22370
rect 13468 22306 13524 22318
rect 13692 22372 13748 22382
rect 13244 21028 13300 21644
rect 13244 20962 13300 20972
rect 13132 20514 13188 20524
rect 13468 20690 13524 20702
rect 13468 20638 13470 20690
rect 13522 20638 13524 20690
rect 13468 20020 13524 20638
rect 13468 19954 13524 19964
rect 13020 19906 13076 19918
rect 13020 19854 13022 19906
rect 13074 19854 13076 19906
rect 12908 19348 12964 19358
rect 13020 19348 13076 19854
rect 12908 19346 13076 19348
rect 12908 19294 12910 19346
rect 12962 19294 13076 19346
rect 12908 19292 13076 19294
rect 12908 19282 12964 19292
rect 13692 19234 13748 22316
rect 13692 19182 13694 19234
rect 13746 19182 13748 19234
rect 13692 19170 13748 19182
rect 12796 19068 12964 19124
rect 12796 18450 12852 18462
rect 12796 18398 12798 18450
rect 12850 18398 12852 18450
rect 12796 18340 12852 18398
rect 12796 18274 12852 18284
rect 12908 17778 12964 19068
rect 13356 18340 13412 18350
rect 13244 18226 13300 18238
rect 13244 18174 13246 18226
rect 13298 18174 13300 18226
rect 13244 17892 13300 18174
rect 13244 17826 13300 17836
rect 12908 17726 12910 17778
rect 12962 17726 12964 17778
rect 12908 17714 12964 17726
rect 13132 16772 13188 16782
rect 13132 16678 13188 16716
rect 12684 16270 12686 16322
rect 12738 16270 12740 16322
rect 12684 16258 12740 16270
rect 12404 15820 12852 15876
rect 12348 15782 12404 15820
rect 12236 15486 12238 15538
rect 12290 15486 12292 15538
rect 12236 15474 12292 15486
rect 12348 15652 12404 15662
rect 12012 15092 12180 15148
rect 11116 13636 11172 13646
rect 11228 13636 11284 13804
rect 11172 13580 11284 13636
rect 11340 13636 11396 13646
rect 11116 13570 11172 13580
rect 11340 13542 11396 13580
rect 11228 13300 11284 13310
rect 11228 12738 11284 13244
rect 11452 13076 11508 15092
rect 11564 14868 11620 14878
rect 11564 14642 11620 14812
rect 11564 14590 11566 14642
rect 11618 14590 11620 14642
rect 11564 14578 11620 14590
rect 11900 14756 11956 14766
rect 11452 12982 11508 13020
rect 11900 14530 11956 14700
rect 11900 14478 11902 14530
rect 11954 14478 11956 14530
rect 11788 12962 11844 12974
rect 11788 12910 11790 12962
rect 11842 12910 11844 12962
rect 11228 12686 11230 12738
rect 11282 12686 11284 12738
rect 11004 12348 11172 12404
rect 10892 12180 10948 12190
rect 10780 12124 10892 12180
rect 10892 12114 10948 12124
rect 11004 12178 11060 12190
rect 11004 12126 11006 12178
rect 11058 12126 11060 12178
rect 11004 11956 11060 12126
rect 10332 11900 10500 11956
rect 10556 11900 11060 11956
rect 10220 11844 10276 11854
rect 10276 11788 10388 11844
rect 10220 11778 10276 11788
rect 10108 10108 10276 10164
rect 10220 10050 10276 10108
rect 10220 9998 10222 10050
rect 10274 9998 10276 10050
rect 10220 9986 10276 9998
rect 10108 9940 10164 9950
rect 10108 9846 10164 9884
rect 10332 9828 10388 11788
rect 10444 9828 10500 11900
rect 10556 11732 10612 11742
rect 10556 11284 10612 11676
rect 11116 11620 11172 12348
rect 11228 11956 11284 12686
rect 11228 11890 11284 11900
rect 11452 12738 11508 12750
rect 11452 12686 11454 12738
rect 11506 12686 11508 12738
rect 11452 11844 11508 12686
rect 11788 12740 11844 12910
rect 11676 12404 11732 12414
rect 11676 12310 11732 12348
rect 10780 11564 11172 11620
rect 11228 11732 11508 11788
rect 11564 12178 11620 12190
rect 11564 12126 11566 12178
rect 11618 12126 11620 12178
rect 10668 11396 10724 11406
rect 10668 11302 10724 11340
rect 10556 11218 10612 11228
rect 10780 10724 10836 11564
rect 11228 11508 11284 11732
rect 11116 11452 11284 11508
rect 11116 11396 11172 11452
rect 11116 11302 11172 11340
rect 11340 11396 11396 11406
rect 11228 11284 11284 11294
rect 11228 11190 11284 11228
rect 11340 11170 11396 11340
rect 11564 11172 11620 12126
rect 11788 11956 11844 12684
rect 11900 12628 11956 14478
rect 12124 14308 12180 15092
rect 12124 14242 12180 14252
rect 12236 14756 12292 14766
rect 12236 14530 12292 14700
rect 12236 14478 12238 14530
rect 12290 14478 12292 14530
rect 12236 14084 12292 14478
rect 12236 14018 12292 14028
rect 12124 13636 12180 13646
rect 12124 13074 12180 13580
rect 12124 13022 12126 13074
rect 12178 13022 12180 13074
rect 12124 13010 12180 13022
rect 12236 13076 12292 13086
rect 12348 13076 12404 15596
rect 12684 15652 12740 15662
rect 12572 15314 12628 15326
rect 12572 15262 12574 15314
rect 12626 15262 12628 15314
rect 12572 14980 12628 15262
rect 12572 14532 12628 14924
rect 12572 14466 12628 14476
rect 12684 14868 12740 15596
rect 12684 14530 12740 14812
rect 12796 14644 12852 15820
rect 13244 15540 13300 15550
rect 13020 15202 13076 15214
rect 13020 15150 13022 15202
rect 13074 15150 13076 15202
rect 13020 15148 13076 15150
rect 13244 15148 13300 15484
rect 13020 15092 13300 15148
rect 12796 14588 13188 14644
rect 12684 14478 12686 14530
rect 12738 14478 12740 14530
rect 12684 14466 12740 14478
rect 12796 14420 12852 14430
rect 12796 14326 12852 14364
rect 12908 14308 12964 14318
rect 12908 14214 12964 14252
rect 12348 13020 12516 13076
rect 12236 12962 12292 13020
rect 12236 12910 12238 12962
rect 12290 12910 12292 12962
rect 12236 12898 12292 12910
rect 11900 12562 11956 12572
rect 12012 12850 12068 12862
rect 12012 12798 12014 12850
rect 12066 12798 12068 12850
rect 12012 12404 12068 12798
rect 12236 12740 12292 12750
rect 12124 12404 12180 12414
rect 12012 12402 12180 12404
rect 12012 12350 12126 12402
rect 12178 12350 12180 12402
rect 12012 12348 12180 12350
rect 12124 12338 12180 12348
rect 11788 11890 11844 11900
rect 11900 12178 11956 12190
rect 11900 12126 11902 12178
rect 11954 12126 11956 12178
rect 11900 11396 11956 12126
rect 12236 11732 12292 12684
rect 12348 12180 12404 12190
rect 12348 12086 12404 12124
rect 12460 12068 12516 13020
rect 12572 12852 12628 12862
rect 12572 12758 12628 12796
rect 13020 12402 13076 12414
rect 13020 12350 13022 12402
rect 13074 12350 13076 12402
rect 12572 12292 12628 12302
rect 13020 12292 13076 12350
rect 12572 12290 13076 12292
rect 12572 12238 12574 12290
rect 12626 12238 13076 12290
rect 12572 12236 13076 12238
rect 12572 12226 12628 12236
rect 13132 12180 13188 14588
rect 12908 12124 13188 12180
rect 12460 12012 12628 12068
rect 12236 11666 12292 11676
rect 12124 11620 12180 11630
rect 12124 11396 12180 11564
rect 12460 11508 12516 11518
rect 12236 11396 12292 11406
rect 12124 11394 12292 11396
rect 12124 11342 12238 11394
rect 12290 11342 12292 11394
rect 12124 11340 12292 11342
rect 11900 11330 11956 11340
rect 12236 11330 12292 11340
rect 11340 11118 11342 11170
rect 11394 11118 11396 11170
rect 10780 10668 11060 10724
rect 11004 9938 11060 10668
rect 11340 10612 11396 11118
rect 11452 11116 11620 11172
rect 11788 11282 11844 11294
rect 11788 11230 11790 11282
rect 11842 11230 11844 11282
rect 11788 11172 11844 11230
rect 12012 11284 12068 11294
rect 12012 11190 12068 11228
rect 11452 10948 11508 11116
rect 11788 11106 11844 11116
rect 12124 11170 12180 11182
rect 12460 11172 12516 11452
rect 12124 11118 12126 11170
rect 12178 11118 12180 11170
rect 11508 10892 11732 10948
rect 11452 10882 11508 10892
rect 11340 10546 11396 10556
rect 11004 9886 11006 9938
rect 11058 9886 11060 9938
rect 10444 9772 10612 9828
rect 10332 9762 10388 9772
rect 9996 9660 10164 9716
rect 8988 9604 9044 9614
rect 8876 9602 9044 9604
rect 8876 9550 8990 9602
rect 9042 9550 9044 9602
rect 8876 9548 9044 9550
rect 8876 9042 8932 9548
rect 8988 9538 9044 9548
rect 9212 9602 9268 9614
rect 9212 9550 9214 9602
rect 9266 9550 9268 9602
rect 8876 8990 8878 9042
rect 8930 8990 8932 9042
rect 8876 8978 8932 8990
rect 8764 8820 8820 8830
rect 8764 8726 8820 8764
rect 8876 8708 8932 8718
rect 8876 8482 8932 8652
rect 9212 8596 9268 9550
rect 8876 8430 8878 8482
rect 8930 8430 8932 8482
rect 8876 8418 8932 8430
rect 8988 8540 9268 8596
rect 9324 9492 9380 9502
rect 8652 8318 8654 8370
rect 8706 8318 8708 8370
rect 8652 8306 8708 8318
rect 8652 7700 8708 7710
rect 8540 7698 8932 7700
rect 8540 7646 8654 7698
rect 8706 7646 8932 7698
rect 8540 7644 8932 7646
rect 8092 7634 8148 7644
rect 8652 7634 8708 7644
rect 7980 6962 8036 6972
rect 7644 5908 7700 5918
rect 7644 5814 7700 5852
rect 7420 5346 7588 5348
rect 7420 5294 7422 5346
rect 7474 5294 7588 5346
rect 7420 5292 7588 5294
rect 7644 5460 7700 5470
rect 6412 5182 6414 5234
rect 6466 5182 6468 5234
rect 6412 5170 6468 5182
rect 6972 5124 7028 5134
rect 7420 5124 7476 5292
rect 6972 5122 7476 5124
rect 6972 5070 6974 5122
rect 7026 5070 7476 5122
rect 6972 5068 7476 5070
rect 6972 5058 7028 5068
rect 6188 4338 6468 4340
rect 6188 4286 6190 4338
rect 6242 4286 6468 4338
rect 6188 4284 6468 4286
rect 6188 4274 6244 4284
rect 6412 3668 6468 4284
rect 6860 4228 6916 4238
rect 6860 4226 7588 4228
rect 6860 4174 6862 4226
rect 6914 4174 7588 4226
rect 6860 4172 7588 4174
rect 6860 4162 6916 4172
rect 7532 3778 7588 4172
rect 7532 3726 7534 3778
rect 7586 3726 7588 3778
rect 7532 3714 7588 3726
rect 6860 3668 6916 3678
rect 7308 3668 7364 3678
rect 6412 3666 7364 3668
rect 6412 3614 6414 3666
rect 6466 3614 6862 3666
rect 6914 3614 7310 3666
rect 7362 3614 7364 3666
rect 6412 3612 7364 3614
rect 6412 3602 6468 3612
rect 6860 3602 6916 3612
rect 7308 3602 7364 3612
rect 7644 3666 7700 5404
rect 7756 5010 7812 5964
rect 7868 6804 7924 6814
rect 8428 6804 8484 6814
rect 7868 5684 7924 6748
rect 7980 6802 8484 6804
rect 7980 6750 8430 6802
rect 8482 6750 8484 6802
rect 7980 6748 8484 6750
rect 7980 5906 8036 6748
rect 8428 6738 8484 6748
rect 8092 6468 8148 6478
rect 8316 6468 8372 6478
rect 8092 6466 8260 6468
rect 8092 6414 8094 6466
rect 8146 6414 8260 6466
rect 8092 6412 8260 6414
rect 8092 6402 8148 6412
rect 7980 5854 7982 5906
rect 8034 5854 8036 5906
rect 7980 5842 8036 5854
rect 8092 6132 8148 6142
rect 8092 5906 8148 6076
rect 8092 5854 8094 5906
rect 8146 5854 8148 5906
rect 8092 5842 8148 5854
rect 8204 5796 8260 6412
rect 8316 6374 8372 6412
rect 8540 6466 8596 6478
rect 8540 6414 8542 6466
rect 8594 6414 8596 6466
rect 8540 6356 8596 6414
rect 8428 6020 8484 6030
rect 8428 5926 8484 5964
rect 8540 5908 8596 6300
rect 8540 5842 8596 5852
rect 8652 5906 8708 5918
rect 8652 5854 8654 5906
rect 8706 5854 8708 5906
rect 8652 5796 8708 5854
rect 8204 5740 8372 5796
rect 7868 5628 8260 5684
rect 8092 5348 8148 5358
rect 7980 5124 8036 5134
rect 7980 5030 8036 5068
rect 8092 5122 8148 5292
rect 8092 5070 8094 5122
rect 8146 5070 8148 5122
rect 8092 5058 8148 5070
rect 8204 5122 8260 5628
rect 8204 5070 8206 5122
rect 8258 5070 8260 5122
rect 8204 5058 8260 5070
rect 7756 4958 7758 5010
rect 7810 4958 7812 5010
rect 7756 4946 7812 4958
rect 8316 4900 8372 5740
rect 8652 5124 8708 5740
rect 8764 5906 8820 5918
rect 8764 5854 8766 5906
rect 8818 5854 8820 5906
rect 8764 5460 8820 5854
rect 8764 5394 8820 5404
rect 8652 5058 8708 5068
rect 8764 5122 8820 5134
rect 8764 5070 8766 5122
rect 8818 5070 8820 5122
rect 8764 5012 8820 5070
rect 8764 4946 8820 4956
rect 8316 4834 8372 4844
rect 7644 3614 7646 3666
rect 7698 3614 7700 3666
rect 7644 3602 7700 3614
rect 8428 4788 8484 4798
rect 8428 3666 8484 4732
rect 8876 4004 8932 7644
rect 8988 7364 9044 8540
rect 9324 8484 9380 9436
rect 9660 9266 9716 9660
rect 9660 9214 9662 9266
rect 9714 9214 9716 9266
rect 9660 9202 9716 9214
rect 9212 8428 9380 8484
rect 9996 9042 10052 9054
rect 9996 8990 9998 9042
rect 10050 8990 10052 9042
rect 9100 8260 9156 8270
rect 9100 8166 9156 8204
rect 9100 7700 9156 7710
rect 9212 7700 9268 8428
rect 9100 7698 9268 7700
rect 9100 7646 9102 7698
rect 9154 7646 9268 7698
rect 9100 7644 9268 7646
rect 9324 8258 9380 8270
rect 9324 8206 9326 8258
rect 9378 8206 9380 8258
rect 9100 7634 9156 7644
rect 8988 6916 9044 7308
rect 9212 7476 9268 7486
rect 9100 6916 9156 6926
rect 8988 6860 9100 6916
rect 9100 6850 9156 6860
rect 8988 6690 9044 6702
rect 8988 6638 8990 6690
rect 9042 6638 9044 6690
rect 8988 6580 9044 6638
rect 9212 6692 9268 7420
rect 9324 6804 9380 8206
rect 9772 8034 9828 8046
rect 9772 7982 9774 8034
rect 9826 7982 9828 8034
rect 9324 6738 9380 6748
rect 9436 7924 9492 7934
rect 9212 6598 9268 6636
rect 8988 6132 9044 6524
rect 9324 6468 9380 6478
rect 9324 6374 9380 6412
rect 8988 6066 9044 6076
rect 8988 5908 9044 5918
rect 8988 4226 9044 5852
rect 8988 4174 8990 4226
rect 9042 4174 9044 4226
rect 8988 4162 9044 4174
rect 8876 3948 9268 4004
rect 8428 3614 8430 3666
rect 8482 3614 8484 3666
rect 8428 3602 8484 3614
rect 8876 3668 8932 3678
rect 8876 3574 8932 3612
rect 5964 3332 6804 3388
rect 4060 3266 4116 3276
rect 3388 2818 3444 2828
rect 6748 2324 6804 3332
rect 9212 2996 9268 3948
rect 9324 2996 9380 3006
rect 9212 2940 9324 2996
rect 9324 2930 9380 2940
rect 9436 2772 9492 7868
rect 9772 7588 9828 7982
rect 9772 7522 9828 7532
rect 9996 7698 10052 8990
rect 10108 8260 10164 9660
rect 10332 9604 10388 9614
rect 10444 9604 10500 9614
rect 10388 9602 10500 9604
rect 10388 9550 10446 9602
rect 10498 9550 10500 9602
rect 10388 9548 10500 9550
rect 10220 8596 10276 8606
rect 10332 8596 10388 9548
rect 10444 9538 10500 9548
rect 10444 9268 10500 9278
rect 10556 9268 10612 9772
rect 11004 9492 11060 9886
rect 11564 10050 11620 10062
rect 11564 9998 11566 10050
rect 11618 9998 11620 10050
rect 11564 9828 11620 9998
rect 11676 10052 11732 10892
rect 12124 10836 12180 11118
rect 11900 10780 12180 10836
rect 12236 11116 12516 11172
rect 11900 10722 11956 10780
rect 11900 10670 11902 10722
rect 11954 10670 11956 10722
rect 11900 10658 11956 10670
rect 11676 9996 12068 10052
rect 12012 9940 12068 9996
rect 12012 9846 12068 9884
rect 11676 9828 11732 9838
rect 11564 9826 11732 9828
rect 11564 9774 11678 9826
rect 11730 9774 11732 9826
rect 11564 9772 11732 9774
rect 11676 9762 11732 9772
rect 11004 9426 11060 9436
rect 10444 9266 10612 9268
rect 10444 9214 10446 9266
rect 10498 9214 10612 9266
rect 10444 9212 10612 9214
rect 10444 9202 10500 9212
rect 11228 9044 11284 9054
rect 10276 8540 10388 8596
rect 10780 8930 10836 8942
rect 10780 8878 10782 8930
rect 10834 8878 10836 8930
rect 10220 8530 10276 8540
rect 10780 8372 10836 8878
rect 10780 8306 10836 8316
rect 10108 8194 10164 8204
rect 10668 8258 10724 8270
rect 10668 8206 10670 8258
rect 10722 8206 10724 8258
rect 10444 8148 10500 8158
rect 10444 8054 10500 8092
rect 10220 8036 10276 8046
rect 10220 7942 10276 7980
rect 9996 7646 9998 7698
rect 10050 7646 10052 7698
rect 9996 7476 10052 7646
rect 10332 7700 10388 7710
rect 10332 7606 10388 7644
rect 9996 7410 10052 7420
rect 9772 7362 9828 7374
rect 10668 7364 10724 8206
rect 11116 8036 11172 8046
rect 11004 8034 11172 8036
rect 11004 7982 11118 8034
rect 11170 7982 11172 8034
rect 11004 7980 11172 7982
rect 10892 7700 10948 7710
rect 10892 7606 10948 7644
rect 10780 7588 10836 7598
rect 10780 7494 10836 7532
rect 9772 7310 9774 7362
rect 9826 7310 9828 7362
rect 9772 6804 9828 7310
rect 9772 6738 9828 6748
rect 10332 7308 10668 7364
rect 9548 6692 9604 6702
rect 9548 6598 9604 6636
rect 9660 6690 9716 6702
rect 9660 6638 9662 6690
rect 9714 6638 9716 6690
rect 9660 6580 9716 6638
rect 9660 5908 9716 6524
rect 10108 6466 10164 6478
rect 10108 6414 10110 6466
rect 10162 6414 10164 6466
rect 10108 6356 10164 6414
rect 10108 6290 10164 6300
rect 9772 6132 9828 6142
rect 10332 6132 10388 7308
rect 10668 7270 10724 7308
rect 11004 6804 11060 7980
rect 11116 7970 11172 7980
rect 11228 7140 11284 8988
rect 12236 8484 12292 11116
rect 12124 8428 12292 8484
rect 12460 10948 12516 10958
rect 11676 8372 11732 8382
rect 11452 8036 11508 8046
rect 11452 8034 11620 8036
rect 11452 7982 11454 8034
rect 11506 7982 11620 8034
rect 11452 7980 11620 7982
rect 11452 7970 11508 7980
rect 11228 7074 11284 7084
rect 11452 6916 11508 6926
rect 10892 6748 11060 6804
rect 11116 6914 11508 6916
rect 11116 6862 11454 6914
rect 11506 6862 11508 6914
rect 11116 6860 11508 6862
rect 9772 6038 9828 6076
rect 9884 6076 10388 6132
rect 10444 6690 10500 6702
rect 10444 6638 10446 6690
rect 10498 6638 10500 6690
rect 9884 5908 9940 6076
rect 9660 5842 9716 5852
rect 9772 5852 9940 5908
rect 9996 5906 10052 5918
rect 9996 5854 9998 5906
rect 10050 5854 10052 5906
rect 9548 5124 9604 5134
rect 9548 5030 9604 5068
rect 9772 4788 9828 5852
rect 9996 5684 10052 5854
rect 10220 5908 10276 5918
rect 10444 5908 10500 6638
rect 10668 6692 10724 6702
rect 10668 6690 10836 6692
rect 10668 6638 10670 6690
rect 10722 6638 10836 6690
rect 10668 6636 10836 6638
rect 10668 6626 10724 6636
rect 10276 5852 10500 5908
rect 10668 6356 10724 6366
rect 10668 5906 10724 6300
rect 10668 5854 10670 5906
rect 10722 5854 10724 5906
rect 10220 5814 10276 5852
rect 10668 5842 10724 5854
rect 10108 5794 10164 5806
rect 10108 5742 10110 5794
rect 10162 5742 10164 5794
rect 10108 5684 10164 5742
rect 10556 5684 10612 5694
rect 10108 5682 10612 5684
rect 10108 5630 10558 5682
rect 10610 5630 10612 5682
rect 10108 5628 10612 5630
rect 9996 5618 10052 5628
rect 10556 5618 10612 5628
rect 10668 5684 10724 5694
rect 10780 5684 10836 6636
rect 10892 6132 10948 6748
rect 11004 6580 11060 6590
rect 11004 6486 11060 6524
rect 10892 6066 10948 6076
rect 11004 6018 11060 6030
rect 11004 5966 11006 6018
rect 11058 5966 11060 6018
rect 10724 5628 10836 5684
rect 10892 5908 10948 5918
rect 10668 5618 10724 5628
rect 10892 5572 10948 5852
rect 10892 5506 10948 5516
rect 11004 5236 11060 5966
rect 11004 5170 11060 5180
rect 11116 5348 11172 6860
rect 11452 6850 11508 6860
rect 11228 6692 11284 6702
rect 11228 6690 11508 6692
rect 11228 6638 11230 6690
rect 11282 6638 11508 6690
rect 11228 6636 11508 6638
rect 11228 6626 11284 6636
rect 11228 6468 11284 6478
rect 11228 5906 11284 6412
rect 11452 6020 11508 6636
rect 11452 5926 11508 5964
rect 11228 5854 11230 5906
rect 11282 5854 11284 5906
rect 11228 5796 11284 5854
rect 11228 5730 11284 5740
rect 11340 5906 11396 5918
rect 11340 5854 11342 5906
rect 11394 5854 11396 5906
rect 10220 5124 10276 5134
rect 9772 4722 9828 4732
rect 9884 5012 9940 5022
rect 9884 4564 9940 4956
rect 9884 4470 9940 4508
rect 10220 4562 10276 5068
rect 11116 4900 11172 5292
rect 10668 4844 11172 4900
rect 10220 4510 10222 4562
rect 10274 4510 10276 4562
rect 10220 4498 10276 4510
rect 10444 4788 10500 4798
rect 10332 4226 10388 4238
rect 10332 4174 10334 4226
rect 10386 4174 10388 4226
rect 9996 3780 10052 3790
rect 9996 3666 10052 3724
rect 10332 3778 10388 4174
rect 10332 3726 10334 3778
rect 10386 3726 10388 3778
rect 10332 3714 10388 3726
rect 9996 3614 9998 3666
rect 10050 3614 10052 3666
rect 9996 3602 10052 3614
rect 10444 3666 10500 4732
rect 10668 4226 10724 4844
rect 10668 4174 10670 4226
rect 10722 4174 10724 4226
rect 10668 4162 10724 4174
rect 10780 4676 10836 4686
rect 10444 3614 10446 3666
rect 10498 3614 10500 3666
rect 10444 3602 10500 3614
rect 10780 3668 10836 4620
rect 11340 3892 11396 5854
rect 11228 3836 11396 3892
rect 11452 5796 11508 5806
rect 11228 3778 11284 3836
rect 11228 3726 11230 3778
rect 11282 3726 11284 3778
rect 11228 3714 11284 3726
rect 9548 3444 9604 3482
rect 9548 3378 9604 3388
rect 9548 2772 9604 2782
rect 9436 2716 9548 2772
rect 9548 2706 9604 2716
rect 6748 2258 6804 2268
rect 10780 1428 10836 3612
rect 11340 3668 11396 3678
rect 11452 3668 11508 5740
rect 11564 4676 11620 7980
rect 11676 6914 11732 8316
rect 12012 8372 12068 8382
rect 12012 8258 12068 8316
rect 12012 8206 12014 8258
rect 12066 8206 12068 8258
rect 12012 8194 12068 8206
rect 12124 6916 12180 8428
rect 12348 8258 12404 8270
rect 12348 8206 12350 8258
rect 12402 8206 12404 8258
rect 12348 7700 12404 8206
rect 11676 6862 11678 6914
rect 11730 6862 11732 6914
rect 11676 6850 11732 6862
rect 12012 6860 12180 6916
rect 12236 7474 12292 7486
rect 12236 7422 12238 7474
rect 12290 7422 12292 7474
rect 11676 6020 11732 6030
rect 11676 5236 11732 5964
rect 12012 5348 12068 6860
rect 12124 6692 12180 6702
rect 12236 6692 12292 7422
rect 12124 6690 12292 6692
rect 12124 6638 12126 6690
rect 12178 6638 12292 6690
rect 12124 6636 12292 6638
rect 12124 6626 12180 6636
rect 12348 6020 12404 7644
rect 12460 6244 12516 10892
rect 12572 9938 12628 12012
rect 12684 11284 12740 11294
rect 12684 11282 12852 11284
rect 12684 11230 12686 11282
rect 12738 11230 12852 11282
rect 12684 11228 12852 11230
rect 12684 11218 12740 11228
rect 12684 10724 12740 10734
rect 12684 10610 12740 10668
rect 12684 10558 12686 10610
rect 12738 10558 12740 10610
rect 12684 10546 12740 10558
rect 12796 10050 12852 11228
rect 12908 10500 12964 12124
rect 13020 11956 13076 11966
rect 13020 11862 13076 11900
rect 13132 11954 13188 11966
rect 13132 11902 13134 11954
rect 13186 11902 13188 11954
rect 13132 11844 13188 11902
rect 13132 11778 13188 11788
rect 12908 10434 12964 10444
rect 13020 11732 13076 11742
rect 12796 9998 12798 10050
rect 12850 9998 12852 10050
rect 12796 9986 12852 9998
rect 12908 10052 12964 10062
rect 12572 9886 12574 9938
rect 12626 9886 12628 9938
rect 12572 9874 12628 9886
rect 12908 9938 12964 9996
rect 12908 9886 12910 9938
rect 12962 9886 12964 9938
rect 12908 9874 12964 9886
rect 12908 8932 12964 8942
rect 12908 8838 12964 8876
rect 12684 8708 12740 8718
rect 12684 7924 12740 8652
rect 12796 8596 12852 8606
rect 12796 8370 12852 8540
rect 12796 8318 12798 8370
rect 12850 8318 12852 8370
rect 12796 8306 12852 8318
rect 12796 8148 12852 8158
rect 12796 8054 12852 8092
rect 12684 7868 12852 7924
rect 12572 6580 12628 6590
rect 12572 6486 12628 6524
rect 12460 6188 12628 6244
rect 12236 5964 12404 6020
rect 12236 5460 12292 5964
rect 12572 5908 12628 6188
rect 12348 5852 12628 5908
rect 12348 5794 12404 5852
rect 12348 5742 12350 5794
rect 12402 5742 12404 5794
rect 12348 5730 12404 5742
rect 12572 5684 12628 5694
rect 12628 5628 12740 5684
rect 12572 5590 12628 5628
rect 12236 5394 12292 5404
rect 12460 5572 12516 5582
rect 12012 5292 12180 5348
rect 11676 5234 12068 5236
rect 11676 5182 11678 5234
rect 11730 5182 12068 5234
rect 11676 5180 12068 5182
rect 11676 5170 11732 5180
rect 12012 5122 12068 5180
rect 12012 5070 12014 5122
rect 12066 5070 12068 5122
rect 12012 5058 12068 5070
rect 12124 4900 12180 5292
rect 12348 5236 12404 5246
rect 12348 5122 12404 5180
rect 12460 5234 12516 5516
rect 12460 5182 12462 5234
rect 12514 5182 12516 5234
rect 12460 5170 12516 5182
rect 12572 5460 12628 5470
rect 12348 5070 12350 5122
rect 12402 5070 12404 5122
rect 12348 5058 12404 5070
rect 12572 5122 12628 5404
rect 12572 5070 12574 5122
rect 12626 5070 12628 5122
rect 12572 5058 12628 5070
rect 12684 5124 12740 5628
rect 12684 5058 12740 5068
rect 12796 4900 12852 7868
rect 12908 7812 12964 7822
rect 12908 6580 12964 7756
rect 13020 6802 13076 11676
rect 13244 10722 13300 15092
rect 13356 12404 13412 18284
rect 13468 17442 13524 17454
rect 13468 17390 13470 17442
rect 13522 17390 13524 17442
rect 13468 17220 13524 17390
rect 13468 17154 13524 17164
rect 13804 17442 13860 24220
rect 14028 23156 14084 24668
rect 14140 24612 14196 27804
rect 14252 26404 14308 26414
rect 14252 26310 14308 26348
rect 14252 25620 14308 25630
rect 14252 25526 14308 25564
rect 14364 25284 14420 28590
rect 15148 27860 15204 30268
rect 15596 29986 15652 31612
rect 15708 30098 15764 33292
rect 16044 33236 16100 34076
rect 15820 33180 16100 33236
rect 16156 34018 16212 35308
rect 16268 35140 16324 35150
rect 16268 34914 16324 35084
rect 16268 34862 16270 34914
rect 16322 34862 16324 34914
rect 16268 34850 16324 34862
rect 16156 33966 16158 34018
rect 16210 33966 16212 34018
rect 15820 31778 15876 33180
rect 15820 31726 15822 31778
rect 15874 31726 15876 31778
rect 15820 31714 15876 31726
rect 15932 32900 15988 32910
rect 15820 30996 15876 31006
rect 15820 30902 15876 30940
rect 15932 30212 15988 32844
rect 16156 32788 16212 33966
rect 16156 32722 16212 32732
rect 16268 33908 16324 33918
rect 16044 32452 16100 32462
rect 16044 32450 16212 32452
rect 16044 32398 16046 32450
rect 16098 32398 16212 32450
rect 16044 32396 16212 32398
rect 16044 32386 16100 32396
rect 16156 31890 16212 32396
rect 16156 31838 16158 31890
rect 16210 31838 16212 31890
rect 16156 31780 16212 31838
rect 16156 31714 16212 31724
rect 16268 31666 16324 33852
rect 16380 32564 16436 32574
rect 16380 32470 16436 32508
rect 16492 32340 16548 35758
rect 16604 35812 16660 38332
rect 16828 35812 16884 35822
rect 16604 35810 16884 35812
rect 16604 35758 16830 35810
rect 16882 35758 16884 35810
rect 16604 35756 16884 35758
rect 16604 35252 16660 35756
rect 16828 35746 16884 35756
rect 16604 35186 16660 35196
rect 16716 35476 16772 35486
rect 16604 34916 16660 34954
rect 16604 34850 16660 34860
rect 16716 34356 16772 35420
rect 16268 31614 16270 31666
rect 16322 31614 16324 31666
rect 16268 31602 16324 31614
rect 16380 32284 16548 32340
rect 16604 34300 16772 34356
rect 16156 31108 16212 31118
rect 16156 31014 16212 31052
rect 16268 30772 16324 30782
rect 15932 30118 15988 30156
rect 16156 30716 16268 30772
rect 15708 30046 15710 30098
rect 15762 30046 15764 30098
rect 15708 30034 15764 30046
rect 15596 29934 15598 29986
rect 15650 29934 15652 29986
rect 15596 29922 15652 29934
rect 15820 29876 15876 29886
rect 15372 29426 15428 29438
rect 15372 29374 15374 29426
rect 15426 29374 15428 29426
rect 15148 27766 15204 27804
rect 15260 28532 15316 28542
rect 15148 26962 15204 26974
rect 15148 26910 15150 26962
rect 15202 26910 15204 26962
rect 14364 25218 14420 25228
rect 14588 26740 14644 26750
rect 14140 24518 14196 24556
rect 14588 24388 14644 26684
rect 15148 26404 15204 26910
rect 15148 26290 15204 26348
rect 15148 26238 15150 26290
rect 15202 26238 15204 26290
rect 15148 26226 15204 26238
rect 14700 25732 14756 25742
rect 14700 25506 14756 25676
rect 14700 25454 14702 25506
rect 14754 25454 14756 25506
rect 14700 25442 14756 25454
rect 15036 25284 15092 25294
rect 14812 24836 14868 24846
rect 14140 24052 14196 24062
rect 14140 23958 14196 23996
rect 14252 23492 14308 23502
rect 14140 23156 14196 23166
rect 14028 23154 14196 23156
rect 14028 23102 14142 23154
rect 14194 23102 14196 23154
rect 14028 23100 14196 23102
rect 14140 22036 14196 23100
rect 14140 21970 14196 21980
rect 14252 22258 14308 23436
rect 14476 23044 14532 23054
rect 14476 22950 14532 22988
rect 14252 22206 14254 22258
rect 14306 22206 14308 22258
rect 14028 20580 14084 20590
rect 14028 20486 14084 20524
rect 14252 20132 14308 22206
rect 14252 20066 14308 20076
rect 14588 18676 14644 24332
rect 14700 24724 14756 24734
rect 14700 23938 14756 24668
rect 14700 23886 14702 23938
rect 14754 23886 14756 23938
rect 14700 23874 14756 23886
rect 14812 20468 14868 24780
rect 14924 24612 14980 24622
rect 14924 22036 14980 24556
rect 15036 23938 15092 25228
rect 15036 23886 15038 23938
rect 15090 23886 15092 23938
rect 15036 23874 15092 23886
rect 15148 22596 15204 22606
rect 15148 22502 15204 22540
rect 15260 22482 15316 28476
rect 15372 27748 15428 29374
rect 15484 28980 15540 28990
rect 15540 28924 15652 28980
rect 15484 28914 15540 28924
rect 15484 27748 15540 27758
rect 15372 27692 15484 27748
rect 15484 27654 15540 27692
rect 15596 26962 15652 28924
rect 15820 27074 15876 29820
rect 15820 27022 15822 27074
rect 15874 27022 15876 27074
rect 15820 27010 15876 27022
rect 15932 28868 15988 28878
rect 15596 26910 15598 26962
rect 15650 26910 15652 26962
rect 15596 26740 15652 26910
rect 15596 26674 15652 26684
rect 15708 26964 15764 26974
rect 15932 26908 15988 28812
rect 16156 26908 16212 30716
rect 16268 30706 16324 30716
rect 16268 30212 16324 30222
rect 16268 28754 16324 30156
rect 16380 29426 16436 32284
rect 16604 31948 16660 34300
rect 16716 34130 16772 34142
rect 16716 34078 16718 34130
rect 16770 34078 16772 34130
rect 16716 32900 16772 34078
rect 17164 33348 17220 38612
rect 18284 38164 18340 40348
rect 18396 40338 18452 40348
rect 20636 40572 21364 40628
rect 21532 40962 21588 40974
rect 21532 40910 21534 40962
rect 21586 40910 21588 40962
rect 19068 40292 19124 40302
rect 19068 40198 19124 40236
rect 20188 40180 20244 40190
rect 19404 40068 19460 40078
rect 19404 39730 19460 40012
rect 19404 39678 19406 39730
rect 19458 39678 19460 39730
rect 19404 39666 19460 39678
rect 19964 39732 20020 39742
rect 19964 39638 20020 39676
rect 18844 39506 18900 39518
rect 18844 39454 18846 39506
rect 18898 39454 18900 39506
rect 18844 38836 18900 39454
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19852 38948 19908 38958
rect 18844 38770 18900 38780
rect 18956 38946 19908 38948
rect 18956 38894 19854 38946
rect 19906 38894 19908 38946
rect 18956 38892 19908 38894
rect 17500 38108 18340 38164
rect 17500 38050 17556 38108
rect 17500 37998 17502 38050
rect 17554 37998 17556 38050
rect 17500 37986 17556 37998
rect 18172 37940 18228 37950
rect 18172 37846 18228 37884
rect 17948 37716 18004 37726
rect 17500 37268 17556 37278
rect 17500 37174 17556 37212
rect 17388 37044 17444 37054
rect 17276 37042 17444 37044
rect 17276 36990 17390 37042
rect 17442 36990 17444 37042
rect 17276 36988 17444 36990
rect 17276 34916 17332 36988
rect 17388 36978 17444 36988
rect 17500 37044 17556 37054
rect 17500 36594 17556 36988
rect 17500 36542 17502 36594
rect 17554 36542 17556 36594
rect 17500 36530 17556 36542
rect 17388 35700 17444 35710
rect 17388 35606 17444 35644
rect 17836 35028 17892 35038
rect 17276 34850 17332 34860
rect 17724 35026 17892 35028
rect 17724 34974 17838 35026
rect 17890 34974 17892 35026
rect 17724 34972 17892 34974
rect 17388 34692 17444 34702
rect 17164 33282 17220 33292
rect 17276 34690 17444 34692
rect 17276 34638 17390 34690
rect 17442 34638 17444 34690
rect 17276 34636 17444 34638
rect 16716 32834 16772 32844
rect 16716 32676 16772 32686
rect 16716 32564 16772 32620
rect 16828 32564 16884 32574
rect 16716 32562 16884 32564
rect 16716 32510 16830 32562
rect 16882 32510 16884 32562
rect 16716 32508 16884 32510
rect 16828 32498 16884 32508
rect 16604 31892 16772 31948
rect 16604 31780 16660 31790
rect 16604 31686 16660 31724
rect 16604 30994 16660 31006
rect 16604 30942 16606 30994
rect 16658 30942 16660 30994
rect 16604 30322 16660 30942
rect 16604 30270 16606 30322
rect 16658 30270 16660 30322
rect 16380 29374 16382 29426
rect 16434 29374 16436 29426
rect 16380 29362 16436 29374
rect 16492 30212 16548 30222
rect 16268 28702 16270 28754
rect 16322 28702 16324 28754
rect 16268 28690 16324 28702
rect 16492 28308 16548 30156
rect 16604 29650 16660 30270
rect 16604 29598 16606 29650
rect 16658 29598 16660 29650
rect 16604 29586 16660 29598
rect 16716 29428 16772 31892
rect 16940 31668 16996 31678
rect 17276 31668 17332 34636
rect 17388 34626 17444 34636
rect 17612 34580 17668 34590
rect 17388 34130 17444 34142
rect 17388 34078 17390 34130
rect 17442 34078 17444 34130
rect 17388 31780 17444 34078
rect 17500 34018 17556 34030
rect 17500 33966 17502 34018
rect 17554 33966 17556 34018
rect 17500 32564 17556 33966
rect 17612 33458 17668 34524
rect 17724 34244 17780 34972
rect 17836 34962 17892 34972
rect 17724 34150 17780 34188
rect 17836 34132 17892 34142
rect 17836 34038 17892 34076
rect 17612 33406 17614 33458
rect 17666 33406 17668 33458
rect 17612 33394 17668 33406
rect 17500 32498 17556 32508
rect 17388 31714 17444 31724
rect 17500 31778 17556 31790
rect 17500 31726 17502 31778
rect 17554 31726 17556 31778
rect 16940 31666 17332 31668
rect 16940 31614 16942 31666
rect 16994 31614 17332 31666
rect 16940 31612 17332 31614
rect 16940 31108 16996 31612
rect 16492 28242 16548 28252
rect 16604 29372 16772 29428
rect 16828 31052 16996 31108
rect 17052 31388 17332 31444
rect 15708 26290 15764 26908
rect 15820 26852 15988 26908
rect 16044 26852 16212 26908
rect 16492 27074 16548 27086
rect 16492 27022 16494 27074
rect 16546 27022 16548 27074
rect 16380 26852 16436 26862
rect 15820 26516 15876 26852
rect 15820 26450 15876 26460
rect 15932 26740 15988 26750
rect 15708 26238 15710 26290
rect 15762 26238 15764 26290
rect 15708 26226 15764 26238
rect 15932 26068 15988 26684
rect 16044 26290 16100 26852
rect 16268 26850 16436 26852
rect 16268 26798 16382 26850
rect 16434 26798 16436 26850
rect 16268 26796 16436 26798
rect 16044 26238 16046 26290
rect 16098 26238 16100 26290
rect 16044 26226 16100 26238
rect 16156 26628 16212 26638
rect 16156 26292 16212 26572
rect 16156 26226 16212 26236
rect 15932 26012 16212 26068
rect 15484 25172 15540 25182
rect 15372 23826 15428 23838
rect 15372 23774 15374 23826
rect 15426 23774 15428 23826
rect 15372 22820 15428 23774
rect 15484 23826 15540 25116
rect 15932 24722 15988 24734
rect 15932 24670 15934 24722
rect 15986 24670 15988 24722
rect 15484 23774 15486 23826
rect 15538 23774 15540 23826
rect 15484 23762 15540 23774
rect 15596 24610 15652 24622
rect 15596 24558 15598 24610
rect 15650 24558 15652 24610
rect 15596 23828 15652 24558
rect 15596 23762 15652 23772
rect 15932 23828 15988 24670
rect 15932 23762 15988 23772
rect 16044 23938 16100 23950
rect 16044 23886 16046 23938
rect 16098 23886 16100 23938
rect 15708 23714 15764 23726
rect 15708 23662 15710 23714
rect 15762 23662 15764 23714
rect 15708 23604 15764 23662
rect 15708 23538 15764 23548
rect 15372 22754 15428 22764
rect 15484 23044 15540 23054
rect 15260 22430 15262 22482
rect 15314 22430 15316 22482
rect 15260 22418 15316 22430
rect 15372 22148 15428 22158
rect 15372 22054 15428 22092
rect 14924 21980 15092 22036
rect 14924 21812 14980 21822
rect 14924 21474 14980 21756
rect 14924 21422 14926 21474
rect 14978 21422 14980 21474
rect 14924 21140 14980 21422
rect 14924 21074 14980 21084
rect 14812 20402 14868 20412
rect 15036 20578 15092 21980
rect 15372 21476 15428 21486
rect 15036 20526 15038 20578
rect 15090 20526 15092 20578
rect 14588 18610 14644 18620
rect 13804 17390 13806 17442
rect 13858 17390 13860 17442
rect 13804 17220 13860 17390
rect 13804 17154 13860 17164
rect 13916 18450 13972 18462
rect 13916 18398 13918 18450
rect 13970 18398 13972 18450
rect 13804 16884 13860 16894
rect 13916 16884 13972 18398
rect 14588 18452 14644 18462
rect 14588 18358 14644 18396
rect 14588 18116 14644 18126
rect 14140 17780 14196 17790
rect 14140 17686 14196 17724
rect 14364 17780 14420 17790
rect 14364 17554 14420 17724
rect 14364 17502 14366 17554
rect 14418 17502 14420 17554
rect 14364 16996 14420 17502
rect 14588 17554 14644 18060
rect 14924 17668 14980 17678
rect 14924 17574 14980 17612
rect 14588 17502 14590 17554
rect 14642 17502 14644 17554
rect 14588 17490 14644 17502
rect 14700 17556 14756 17566
rect 14700 17462 14756 17500
rect 14364 16930 14420 16940
rect 14700 17220 14756 17230
rect 13860 16828 13972 16884
rect 13804 16790 13860 16828
rect 14588 16772 14644 16782
rect 14140 16324 14196 16334
rect 13916 16210 13972 16222
rect 13916 16158 13918 16210
rect 13970 16158 13972 16210
rect 13580 15988 13636 15998
rect 13468 15204 13524 15214
rect 13468 14754 13524 15148
rect 13468 14702 13470 14754
rect 13522 14702 13524 14754
rect 13468 14690 13524 14702
rect 13580 14642 13636 15932
rect 13580 14590 13582 14642
rect 13634 14590 13636 14642
rect 13580 14578 13636 14590
rect 13916 15316 13972 16158
rect 13804 14530 13860 14542
rect 13804 14478 13806 14530
rect 13858 14478 13860 14530
rect 13804 14084 13860 14478
rect 13804 14018 13860 14028
rect 13916 13748 13972 15260
rect 13356 12338 13412 12348
rect 13468 13634 13524 13646
rect 13468 13582 13470 13634
rect 13522 13582 13524 13634
rect 13468 12180 13524 13582
rect 13804 13634 13860 13646
rect 13804 13582 13806 13634
rect 13858 13582 13860 13634
rect 13804 13300 13860 13582
rect 13804 13234 13860 13244
rect 13916 12962 13972 13692
rect 13916 12910 13918 12962
rect 13970 12910 13972 12962
rect 13916 12852 13972 12910
rect 13468 12114 13524 12124
rect 13692 12796 13972 12852
rect 14028 13412 14084 13422
rect 13356 11954 13412 11966
rect 13356 11902 13358 11954
rect 13410 11902 13412 11954
rect 13356 10948 13412 11902
rect 13692 11620 13748 12796
rect 13916 12628 13972 12638
rect 13804 12516 13860 12526
rect 13804 11732 13860 12460
rect 13804 11666 13860 11676
rect 13916 12290 13972 12572
rect 14028 12402 14084 13356
rect 14028 12350 14030 12402
rect 14082 12350 14084 12402
rect 14028 12338 14084 12350
rect 13916 12238 13918 12290
rect 13970 12238 13972 12290
rect 13356 10882 13412 10892
rect 13580 11564 13748 11620
rect 13580 11394 13636 11564
rect 13580 11342 13582 11394
rect 13634 11342 13636 11394
rect 13244 10670 13246 10722
rect 13298 10670 13300 10722
rect 13244 10658 13300 10670
rect 13356 10724 13412 10734
rect 13580 10724 13636 11342
rect 13916 11060 13972 12238
rect 14028 12180 14084 12190
rect 14028 11284 14084 12124
rect 14140 11956 14196 16268
rect 14252 14420 14308 14430
rect 14252 14326 14308 14364
rect 14476 14418 14532 14430
rect 14476 14366 14478 14418
rect 14530 14366 14532 14418
rect 14476 14196 14532 14366
rect 14588 14306 14644 16716
rect 14588 14254 14590 14306
rect 14642 14254 14644 14306
rect 14588 14242 14644 14254
rect 14700 16436 14756 17164
rect 14812 16996 14868 17006
rect 14812 16882 14868 16940
rect 14812 16830 14814 16882
rect 14866 16830 14868 16882
rect 14812 16818 14868 16830
rect 14476 14130 14532 14140
rect 14700 14084 14756 16380
rect 15036 15764 15092 20526
rect 15260 21028 15316 21038
rect 15260 19234 15316 20972
rect 15372 20690 15428 21420
rect 15372 20638 15374 20690
rect 15426 20638 15428 20690
rect 15372 20626 15428 20638
rect 15260 19182 15262 19234
rect 15314 19182 15316 19234
rect 15260 19170 15316 19182
rect 15484 20244 15540 22988
rect 16044 22932 16100 23886
rect 15932 22876 16044 22932
rect 15932 22370 15988 22876
rect 16044 22866 16100 22876
rect 15932 22318 15934 22370
rect 15986 22318 15988 22370
rect 15932 22306 15988 22318
rect 15484 19122 15540 20188
rect 15484 19070 15486 19122
rect 15538 19070 15540 19122
rect 15484 19058 15540 19070
rect 15596 22148 15652 22158
rect 15596 20916 15652 22092
rect 15708 21588 15764 21598
rect 15708 21586 15876 21588
rect 15708 21534 15710 21586
rect 15762 21534 15876 21586
rect 15708 21532 15876 21534
rect 15708 21522 15764 21532
rect 15708 20916 15764 20926
rect 15596 20914 15764 20916
rect 15596 20862 15710 20914
rect 15762 20862 15764 20914
rect 15596 20860 15764 20862
rect 15596 19684 15652 20860
rect 15708 20850 15764 20860
rect 15820 20916 15876 21532
rect 15820 20850 15876 20860
rect 15932 21028 15988 21038
rect 15708 20692 15764 20702
rect 15708 20244 15764 20636
rect 15708 20150 15764 20188
rect 15932 20468 15988 20972
rect 15036 15698 15092 15708
rect 15148 18564 15204 18574
rect 15148 15428 15204 18508
rect 15372 17556 15428 17566
rect 15372 17554 15540 17556
rect 15372 17502 15374 17554
rect 15426 17502 15540 17554
rect 15372 17500 15540 17502
rect 15372 17490 15428 17500
rect 15372 16884 15428 16894
rect 15372 16770 15428 16828
rect 15372 16718 15374 16770
rect 15426 16718 15428 16770
rect 15372 16706 15428 16718
rect 15036 15372 15204 15428
rect 15036 14980 15092 15372
rect 15148 15202 15204 15214
rect 15148 15150 15150 15202
rect 15202 15150 15204 15202
rect 15148 15148 15204 15150
rect 15484 15148 15540 17500
rect 15148 15092 15316 15148
rect 15036 14924 15204 14980
rect 15036 14530 15092 14542
rect 15036 14478 15038 14530
rect 15090 14478 15092 14530
rect 14812 14420 14868 14430
rect 15036 14420 15092 14478
rect 14812 14418 15092 14420
rect 14812 14366 14814 14418
rect 14866 14366 15092 14418
rect 14812 14364 15092 14366
rect 14812 14308 14868 14364
rect 14812 14242 14868 14252
rect 14700 14028 14868 14084
rect 14364 13746 14420 13758
rect 14364 13694 14366 13746
rect 14418 13694 14420 13746
rect 14364 13636 14420 13694
rect 14364 13570 14420 13580
rect 14252 13300 14308 13310
rect 14252 12402 14308 13244
rect 14252 12350 14254 12402
rect 14306 12350 14308 12402
rect 14252 12338 14308 12350
rect 14364 13188 14420 13198
rect 14364 12180 14420 13132
rect 14588 12852 14644 12862
rect 14588 12758 14644 12796
rect 14588 12404 14644 12414
rect 14644 12348 14756 12404
rect 14588 12310 14644 12348
rect 14476 12292 14532 12302
rect 14476 12198 14532 12236
rect 14364 12114 14420 12124
rect 14588 11956 14644 11966
rect 14140 11954 14644 11956
rect 14140 11902 14590 11954
rect 14642 11902 14644 11954
rect 14140 11900 14644 11902
rect 14588 11890 14644 11900
rect 14364 11732 14420 11742
rect 14364 11506 14420 11676
rect 14364 11454 14366 11506
rect 14418 11454 14420 11506
rect 14364 11442 14420 11454
rect 14588 11620 14644 11630
rect 14028 11228 14420 11284
rect 13916 11004 14196 11060
rect 14028 10836 14084 10846
rect 14028 10742 14084 10780
rect 13356 10722 13524 10724
rect 13356 10670 13358 10722
rect 13410 10670 13524 10722
rect 13356 10668 13524 10670
rect 13356 10658 13412 10668
rect 13468 10500 13524 10668
rect 13468 10434 13524 10444
rect 13580 9042 13636 10668
rect 13804 10722 13860 10734
rect 13804 10670 13806 10722
rect 13858 10670 13860 10722
rect 13692 10610 13748 10622
rect 13692 10558 13694 10610
rect 13746 10558 13748 10610
rect 13692 10276 13748 10558
rect 13804 10500 13860 10670
rect 13804 10434 13860 10444
rect 14140 10388 14196 11004
rect 13916 10332 14196 10388
rect 14252 10722 14308 10734
rect 14252 10670 14254 10722
rect 14306 10670 14308 10722
rect 13916 10276 13972 10332
rect 13692 10220 13972 10276
rect 14252 9828 14308 10670
rect 14028 9772 14308 9828
rect 13580 8990 13582 9042
rect 13634 8990 13636 9042
rect 13580 8978 13636 8990
rect 13804 9714 13860 9726
rect 13804 9662 13806 9714
rect 13858 9662 13860 9714
rect 13804 8708 13860 9662
rect 13804 8642 13860 8652
rect 13916 9602 13972 9614
rect 13916 9550 13918 9602
rect 13970 9550 13972 9602
rect 13244 8596 13300 8606
rect 13020 6750 13022 6802
rect 13074 6750 13076 6802
rect 13020 6738 13076 6750
rect 13132 8540 13244 8596
rect 12908 6524 13076 6580
rect 12908 6132 12964 6142
rect 12908 5906 12964 6076
rect 12908 5854 12910 5906
rect 12962 5854 12964 5906
rect 12908 5842 12964 5854
rect 12124 4844 12740 4900
rect 11564 4610 11620 4620
rect 12236 4676 12292 4686
rect 11340 3666 11508 3668
rect 11340 3614 11342 3666
rect 11394 3614 11508 3666
rect 11340 3612 11508 3614
rect 12236 3666 12292 4620
rect 12684 4004 12740 4844
rect 12796 4834 12852 4844
rect 13020 4452 13076 6524
rect 13132 6020 13188 8540
rect 13244 8530 13300 8540
rect 13916 8484 13972 9550
rect 14028 9380 14084 9772
rect 14140 9604 14196 9614
rect 14140 9602 14308 9604
rect 14140 9550 14142 9602
rect 14194 9550 14308 9602
rect 14140 9548 14308 9550
rect 14140 9538 14196 9548
rect 14028 9324 14196 9380
rect 14028 9042 14084 9054
rect 14028 8990 14030 9042
rect 14082 8990 14084 9042
rect 14028 8820 14084 8990
rect 14028 8754 14084 8764
rect 13916 8418 13972 8428
rect 13468 8370 13524 8382
rect 13468 8318 13470 8370
rect 13522 8318 13524 8370
rect 13468 8148 13524 8318
rect 13468 7588 13524 8092
rect 13468 7522 13524 7532
rect 13804 8260 13860 8270
rect 13804 7586 13860 8204
rect 13804 7534 13806 7586
rect 13858 7534 13860 7586
rect 13804 7522 13860 7534
rect 14140 7364 14196 9324
rect 14252 9154 14308 9548
rect 14252 9102 14254 9154
rect 14306 9102 14308 9154
rect 14252 9090 14308 9102
rect 14364 7474 14420 11228
rect 14476 11060 14532 11070
rect 14476 10612 14532 11004
rect 14588 10836 14644 11564
rect 14588 10770 14644 10780
rect 14476 10518 14532 10556
rect 14700 10388 14756 12348
rect 14812 11284 14868 14028
rect 14812 11218 14868 11228
rect 14924 13858 14980 13870
rect 14924 13806 14926 13858
rect 14978 13806 14980 13858
rect 14924 11956 14980 13806
rect 15148 13076 15204 14924
rect 15260 14642 15316 15092
rect 15260 14590 15262 14642
rect 15314 14590 15316 14642
rect 15260 14578 15316 14590
rect 15372 15092 15540 15148
rect 15260 13972 15316 13982
rect 15260 13878 15316 13916
rect 15036 13020 15204 13076
rect 15036 12404 15092 13020
rect 15036 12338 15092 12348
rect 15148 12852 15204 12862
rect 15148 12402 15204 12796
rect 15372 12516 15428 15092
rect 15484 14418 15540 14430
rect 15484 14366 15486 14418
rect 15538 14366 15540 14418
rect 15484 13524 15540 14366
rect 15484 13458 15540 13468
rect 15148 12350 15150 12402
rect 15202 12350 15204 12402
rect 15148 12338 15204 12350
rect 15260 12460 15428 12516
rect 15036 12178 15092 12190
rect 15036 12126 15038 12178
rect 15090 12126 15092 12178
rect 15036 11956 15092 12126
rect 14924 11900 15036 11956
rect 14588 10332 14756 10388
rect 14812 11060 14868 11070
rect 14476 8932 14532 8942
rect 14476 8838 14532 8876
rect 14364 7422 14366 7474
rect 14418 7422 14420 7474
rect 14364 7410 14420 7422
rect 14252 7364 14308 7374
rect 14140 7308 14252 7364
rect 14588 7364 14644 10332
rect 14812 9940 14868 11004
rect 14924 10722 14980 11900
rect 15036 11890 15092 11900
rect 15036 11732 15092 11742
rect 15036 10834 15092 11676
rect 15260 11508 15316 12460
rect 15596 12404 15652 19628
rect 15932 19458 15988 20412
rect 15932 19406 15934 19458
rect 15986 19406 15988 19458
rect 15708 16772 15764 16782
rect 15708 14530 15764 16716
rect 15932 15876 15988 19406
rect 16156 17780 16212 26012
rect 16268 25394 16324 26796
rect 16380 26786 16436 26796
rect 16492 26628 16548 27022
rect 16604 26740 16660 29372
rect 16828 29316 16884 31052
rect 16604 26674 16660 26684
rect 16716 29260 16884 29316
rect 16940 30436 16996 30446
rect 16492 26562 16548 26572
rect 16268 25342 16270 25394
rect 16322 25342 16324 25394
rect 16268 25330 16324 25342
rect 16380 26516 16436 26526
rect 16380 26402 16436 26460
rect 16716 26404 16772 29260
rect 16940 29204 16996 30380
rect 16828 29148 16996 29204
rect 16828 27746 16884 29148
rect 16940 28980 16996 28990
rect 16940 28532 16996 28924
rect 17052 28756 17108 31388
rect 17164 31220 17220 31230
rect 17276 31220 17332 31388
rect 17388 31220 17444 31230
rect 17276 31218 17444 31220
rect 17276 31166 17390 31218
rect 17442 31166 17444 31218
rect 17276 31164 17444 31166
rect 17164 30434 17220 31164
rect 17388 31154 17444 31164
rect 17500 30884 17556 31726
rect 17500 30818 17556 30828
rect 17612 30994 17668 31006
rect 17612 30942 17614 30994
rect 17666 30942 17668 30994
rect 17276 30772 17332 30782
rect 17276 30678 17332 30716
rect 17164 30382 17166 30434
rect 17218 30382 17220 30434
rect 17164 30370 17220 30382
rect 17612 30324 17668 30942
rect 17948 30994 18004 37660
rect 18284 36482 18340 38108
rect 18396 38722 18452 38734
rect 18396 38670 18398 38722
rect 18450 38670 18452 38722
rect 18396 37716 18452 38670
rect 18956 38722 19012 38892
rect 19852 38882 19908 38892
rect 20076 38836 20132 38846
rect 18956 38670 18958 38722
rect 19010 38670 19012 38722
rect 18396 37650 18452 37660
rect 18508 38610 18564 38622
rect 18508 38558 18510 38610
rect 18562 38558 18564 38610
rect 18396 37154 18452 37166
rect 18396 37102 18398 37154
rect 18450 37102 18452 37154
rect 18396 37044 18452 37102
rect 18396 36978 18452 36988
rect 18284 36430 18286 36482
rect 18338 36430 18340 36482
rect 18284 36418 18340 36430
rect 18172 36260 18228 36270
rect 18172 35810 18228 36204
rect 18172 35758 18174 35810
rect 18226 35758 18228 35810
rect 18172 35746 18228 35758
rect 18284 35700 18340 35710
rect 18172 34914 18228 34926
rect 18172 34862 18174 34914
rect 18226 34862 18228 34914
rect 18060 34132 18116 34142
rect 18060 31892 18116 34076
rect 18172 33348 18228 34862
rect 18284 34468 18340 35644
rect 18284 34412 18452 34468
rect 18284 34132 18340 34142
rect 18284 34038 18340 34076
rect 18172 32004 18228 33292
rect 18172 31938 18228 31948
rect 18396 33346 18452 34412
rect 18508 34132 18564 38558
rect 18732 37266 18788 37278
rect 18732 37214 18734 37266
rect 18786 37214 18788 37266
rect 18732 37156 18788 37214
rect 18844 37156 18900 37166
rect 18732 37100 18844 37156
rect 18844 37090 18900 37100
rect 18620 36652 18900 36708
rect 18620 34914 18676 36652
rect 18732 36482 18788 36494
rect 18732 36430 18734 36482
rect 18786 36430 18788 36482
rect 18732 35026 18788 36430
rect 18844 36484 18900 36652
rect 18844 36390 18900 36428
rect 18956 35700 19012 38670
rect 19404 38722 19460 38734
rect 19404 38670 19406 38722
rect 19458 38670 19460 38722
rect 19404 38610 19460 38670
rect 19404 38558 19406 38610
rect 19458 38558 19460 38610
rect 19404 38546 19460 38558
rect 20076 38610 20132 38780
rect 20076 38558 20078 38610
rect 20130 38558 20132 38610
rect 20076 38164 20132 38558
rect 19628 38108 20132 38164
rect 19180 37378 19236 37390
rect 19180 37326 19182 37378
rect 19234 37326 19236 37378
rect 19068 37266 19124 37278
rect 19068 37214 19070 37266
rect 19122 37214 19124 37266
rect 19068 36820 19124 37214
rect 19068 36754 19124 36764
rect 19180 36596 19236 37326
rect 19404 37266 19460 37278
rect 19404 37214 19406 37266
rect 19458 37214 19460 37266
rect 19404 36708 19460 37214
rect 19628 37156 19684 38108
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19740 37156 19796 37166
rect 19628 37154 19796 37156
rect 19628 37102 19742 37154
rect 19794 37102 19796 37154
rect 19628 37100 19796 37102
rect 19740 37090 19796 37100
rect 19404 36642 19460 36652
rect 19852 37044 19908 37054
rect 20188 37044 20244 40124
rect 20524 39844 20580 39854
rect 20524 39506 20580 39788
rect 20636 39730 20692 40572
rect 20636 39678 20638 39730
rect 20690 39678 20692 39730
rect 20636 39666 20692 39678
rect 20972 40404 21028 40414
rect 20748 39620 20804 39630
rect 20748 39526 20804 39564
rect 20524 39454 20526 39506
rect 20578 39454 20580 39506
rect 20524 39442 20580 39454
rect 20972 39058 21028 40348
rect 21532 40404 21588 40910
rect 21532 40338 21588 40348
rect 21196 40290 21252 40302
rect 21196 40238 21198 40290
rect 21250 40238 21252 40290
rect 21196 39844 21252 40238
rect 21196 39778 21252 39788
rect 21420 40292 21476 40302
rect 21420 39842 21476 40236
rect 21420 39790 21422 39842
rect 21474 39790 21476 39842
rect 21420 39778 21476 39790
rect 21532 39508 21588 39518
rect 21644 39508 21700 42924
rect 21980 42754 22036 42766
rect 21980 42702 21982 42754
rect 22034 42702 22036 42754
rect 21756 42642 21812 42654
rect 21756 42590 21758 42642
rect 21810 42590 21812 42642
rect 21756 42532 21812 42590
rect 21756 42466 21812 42476
rect 21868 42084 21924 42094
rect 21980 42084 22036 42702
rect 21868 42082 22036 42084
rect 21868 42030 21870 42082
rect 21922 42030 22036 42082
rect 21868 42028 22036 42030
rect 21868 42018 21924 42028
rect 21868 41186 21924 41198
rect 21868 41134 21870 41186
rect 21922 41134 21924 41186
rect 21756 40626 21812 40638
rect 21756 40574 21758 40626
rect 21810 40574 21812 40626
rect 21756 39842 21812 40574
rect 21756 39790 21758 39842
rect 21810 39790 21812 39842
rect 21756 39778 21812 39790
rect 21868 39620 21924 41134
rect 21980 41188 22036 42028
rect 22092 41410 22148 43372
rect 22428 43334 22484 43372
rect 22316 42980 22372 42990
rect 22540 42980 22596 43708
rect 22764 43650 22820 43708
rect 24332 43762 24388 44268
rect 24556 44322 24612 45052
rect 24556 44270 24558 44322
rect 24610 44270 24612 44322
rect 24556 43764 24612 44270
rect 24332 43710 24334 43762
rect 24386 43710 24388 43762
rect 24332 43698 24388 43710
rect 24444 43762 24612 43764
rect 24444 43710 24558 43762
rect 24610 43710 24612 43762
rect 24444 43708 24612 43710
rect 22764 43598 22766 43650
rect 22818 43598 22820 43650
rect 22316 42978 22596 42980
rect 22316 42926 22318 42978
rect 22370 42926 22596 42978
rect 22316 42924 22596 42926
rect 22652 43538 22708 43550
rect 22652 43486 22654 43538
rect 22706 43486 22708 43538
rect 22316 42914 22372 42924
rect 22316 42532 22372 42542
rect 22316 42194 22372 42476
rect 22316 42142 22318 42194
rect 22370 42142 22372 42194
rect 22316 42130 22372 42142
rect 22540 42196 22596 42206
rect 22652 42196 22708 43486
rect 22540 42194 22708 42196
rect 22540 42142 22542 42194
rect 22594 42142 22708 42194
rect 22540 42140 22708 42142
rect 22540 42130 22596 42140
rect 22204 42082 22260 42094
rect 22204 42030 22206 42082
rect 22258 42030 22260 42082
rect 22204 41860 22260 42030
rect 22764 41970 22820 43598
rect 24220 43652 24276 43662
rect 24220 43558 24276 43596
rect 22988 43538 23044 43550
rect 22988 43486 22990 43538
rect 23042 43486 23044 43538
rect 22876 42866 22932 42878
rect 22876 42814 22878 42866
rect 22930 42814 22932 42866
rect 22876 42196 22932 42814
rect 22988 42754 23044 43486
rect 23772 43538 23828 43550
rect 23772 43486 23774 43538
rect 23826 43486 23828 43538
rect 23436 43428 23492 43438
rect 23772 43428 23828 43486
rect 24332 43540 24388 43550
rect 23436 43426 23828 43428
rect 23436 43374 23438 43426
rect 23490 43374 23828 43426
rect 23436 43372 23828 43374
rect 23996 43428 24052 43438
rect 23436 43316 23492 43372
rect 23436 43250 23492 43260
rect 23660 42868 23716 42878
rect 23660 42774 23716 42812
rect 22988 42702 22990 42754
rect 23042 42702 23044 42754
rect 22988 42196 23044 42702
rect 23100 42196 23156 42206
rect 22988 42194 23156 42196
rect 22988 42142 23102 42194
rect 23154 42142 23156 42194
rect 22988 42140 23156 42142
rect 22876 42130 22932 42140
rect 23100 42130 23156 42140
rect 23324 42196 23380 42206
rect 23324 42102 23380 42140
rect 22764 41918 22766 41970
rect 22818 41918 22820 41970
rect 22764 41906 22820 41918
rect 22204 41794 22260 41804
rect 23212 41860 23268 41870
rect 23212 41766 23268 41804
rect 23772 41858 23828 41870
rect 23772 41806 23774 41858
rect 23826 41806 23828 41858
rect 23772 41748 23828 41806
rect 23772 41682 23828 41692
rect 22092 41358 22094 41410
rect 22146 41358 22148 41410
rect 22092 41346 22148 41358
rect 22876 41410 22932 41422
rect 22876 41358 22878 41410
rect 22930 41358 22932 41410
rect 22876 41298 22932 41358
rect 22876 41246 22878 41298
rect 22930 41246 22932 41298
rect 22876 41234 22932 41246
rect 23324 41410 23380 41422
rect 23324 41358 23326 41410
rect 23378 41358 23380 41410
rect 23324 41298 23380 41358
rect 23324 41246 23326 41298
rect 23378 41246 23380 41298
rect 21980 41132 22148 41188
rect 21980 40404 22036 40414
rect 21980 40310 22036 40348
rect 21980 39620 22036 39630
rect 21868 39618 22036 39620
rect 21868 39566 21982 39618
rect 22034 39566 22036 39618
rect 21868 39564 22036 39566
rect 21980 39554 22036 39564
rect 20972 39006 20974 39058
rect 21026 39006 21028 39058
rect 20972 38994 21028 39006
rect 21196 39506 21700 39508
rect 21196 39454 21534 39506
rect 21586 39454 21700 39506
rect 21196 39452 21700 39454
rect 20300 38946 20356 38958
rect 20300 38894 20302 38946
rect 20354 38894 20356 38946
rect 20300 38612 20356 38894
rect 20748 38836 20804 38846
rect 20412 38724 20468 38762
rect 20748 38742 20804 38780
rect 20972 38834 21028 38846
rect 20972 38782 20974 38834
rect 21026 38782 21028 38834
rect 20412 38658 20468 38668
rect 20300 38162 20356 38556
rect 20972 38612 21028 38782
rect 20972 38546 21028 38556
rect 20300 38110 20302 38162
rect 20354 38110 20356 38162
rect 20300 37378 20356 38110
rect 21196 38052 21252 39452
rect 21532 39442 21588 39452
rect 21308 38948 21364 38958
rect 21756 38948 21812 38958
rect 21308 38946 21812 38948
rect 21308 38894 21310 38946
rect 21362 38894 21758 38946
rect 21810 38894 21812 38946
rect 21308 38892 21812 38894
rect 21308 38882 21364 38892
rect 21756 38882 21812 38892
rect 21868 38946 21924 38958
rect 21868 38894 21870 38946
rect 21922 38894 21924 38946
rect 21420 38724 21476 38734
rect 21644 38724 21700 38734
rect 21476 38722 21700 38724
rect 21476 38670 21646 38722
rect 21698 38670 21700 38722
rect 21476 38668 21700 38670
rect 21868 38668 21924 38894
rect 21420 38658 21476 38668
rect 21644 38658 21700 38668
rect 21756 38612 21924 38668
rect 21308 38052 21364 38062
rect 21196 38050 21364 38052
rect 21196 37998 21310 38050
rect 21362 37998 21364 38050
rect 21196 37996 21364 37998
rect 20300 37326 20302 37378
rect 20354 37326 20356 37378
rect 20300 37314 20356 37326
rect 20748 37828 20804 37838
rect 20748 37044 20804 37772
rect 20188 36988 20692 37044
rect 19180 36530 19236 36540
rect 19292 36428 19684 36484
rect 19180 36370 19236 36382
rect 19180 36318 19182 36370
rect 19234 36318 19236 36370
rect 19068 36260 19124 36270
rect 19068 36166 19124 36204
rect 18956 35634 19012 35644
rect 18732 34974 18734 35026
rect 18786 34974 18788 35026
rect 18732 34962 18788 34974
rect 19180 35588 19236 36318
rect 18620 34862 18622 34914
rect 18674 34862 18676 34914
rect 18620 34692 18676 34862
rect 18844 34916 18900 34926
rect 19180 34916 19236 35532
rect 18844 34914 19236 34916
rect 18844 34862 18846 34914
rect 18898 34862 19236 34914
rect 18844 34860 19236 34862
rect 18844 34850 18900 34860
rect 19292 34692 19348 36428
rect 19628 36314 19684 36428
rect 19404 36258 19460 36270
rect 19404 36206 19406 36258
rect 19458 36206 19460 36258
rect 19404 34858 19460 36206
rect 19516 36260 19572 36270
rect 19628 36262 19630 36314
rect 19682 36262 19684 36314
rect 19740 36372 19796 36382
rect 19740 36278 19796 36316
rect 19628 36250 19684 36262
rect 19852 36260 19908 36988
rect 20188 36820 20244 36830
rect 19964 36484 20020 36494
rect 19964 36390 20020 36428
rect 19516 35812 19572 36204
rect 19852 36194 19908 36204
rect 20188 36260 20244 36764
rect 20636 36708 20692 36988
rect 20748 36978 20804 36988
rect 20636 36652 20916 36708
rect 20412 36596 20468 36606
rect 20412 36484 20468 36540
rect 20188 36194 20244 36204
rect 20300 36482 20468 36484
rect 20300 36430 20414 36482
rect 20466 36430 20468 36482
rect 20300 36428 20468 36430
rect 19836 36092 20100 36102
rect 19628 36036 19684 36046
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19628 35924 19684 35980
rect 19628 35868 19796 35924
rect 19516 35756 19684 35812
rect 19516 35140 19572 35150
rect 19516 35046 19572 35084
rect 19404 34806 19406 34858
rect 19458 34806 19460 34858
rect 19404 34794 19460 34806
rect 18620 34636 19236 34692
rect 19292 34636 19460 34692
rect 19180 34580 19236 34636
rect 19180 34524 19348 34580
rect 19180 34356 19236 34366
rect 18956 34300 19180 34356
rect 18508 34066 18564 34076
rect 18732 34132 18788 34142
rect 18732 34020 18788 34076
rect 18732 34018 18900 34020
rect 18732 33966 18734 34018
rect 18786 33966 18900 34018
rect 18732 33964 18900 33966
rect 18732 33954 18788 33964
rect 18396 33294 18398 33346
rect 18450 33294 18452 33346
rect 18060 31556 18116 31836
rect 18172 31668 18228 31678
rect 18172 31574 18228 31612
rect 18060 31490 18116 31500
rect 17948 30942 17950 30994
rect 18002 30942 18004 30994
rect 17948 30772 18004 30942
rect 17948 30706 18004 30716
rect 18172 31444 18228 31454
rect 17276 30268 17668 30324
rect 17836 30324 17892 30334
rect 17052 28700 17220 28756
rect 17052 28532 17108 28542
rect 16940 28530 17108 28532
rect 16940 28478 17054 28530
rect 17106 28478 17108 28530
rect 16940 28476 17108 28478
rect 17052 28466 17108 28476
rect 17164 27972 17220 28700
rect 17276 28196 17332 30268
rect 17836 30210 17892 30268
rect 17836 30158 17838 30210
rect 17890 30158 17892 30210
rect 17836 30146 17892 30158
rect 18060 30210 18116 30222
rect 18060 30158 18062 30210
rect 18114 30158 18116 30210
rect 17500 30100 17556 30110
rect 17724 30100 17780 30110
rect 17556 30098 17780 30100
rect 17556 30046 17726 30098
rect 17778 30046 17780 30098
rect 17556 30044 17780 30046
rect 17388 29876 17444 29886
rect 17388 29426 17444 29820
rect 17388 29374 17390 29426
rect 17442 29374 17444 29426
rect 17388 29362 17444 29374
rect 17388 28644 17444 28654
rect 17500 28644 17556 30044
rect 17724 30034 17780 30044
rect 18060 29876 18116 30158
rect 17388 28642 17556 28644
rect 17388 28590 17390 28642
rect 17442 28590 17556 28642
rect 17388 28588 17556 28590
rect 17612 29820 18116 29876
rect 17612 29428 17668 29820
rect 18060 29652 18116 29662
rect 18172 29652 18228 31388
rect 18396 30884 18452 33294
rect 18732 32116 18788 32126
rect 18396 30818 18452 30828
rect 18620 32060 18732 32116
rect 18060 29650 18228 29652
rect 18060 29598 18062 29650
rect 18114 29598 18228 29650
rect 18060 29596 18228 29598
rect 18396 30660 18452 30670
rect 18060 29586 18116 29596
rect 17948 29540 18004 29550
rect 17948 29446 18004 29484
rect 17388 28578 17444 28588
rect 17276 28140 17556 28196
rect 17164 27906 17220 27916
rect 16828 27694 16830 27746
rect 16882 27694 16884 27746
rect 16828 26964 16884 27694
rect 17276 27748 17332 27758
rect 16828 26898 16884 26908
rect 16940 27636 16996 27646
rect 16380 26350 16382 26402
rect 16434 26350 16436 26402
rect 16268 25172 16324 25182
rect 16268 20018 16324 25116
rect 16380 24836 16436 26350
rect 16492 26348 16772 26404
rect 16492 26178 16548 26348
rect 16492 26126 16494 26178
rect 16546 26126 16548 26178
rect 16492 26114 16548 26126
rect 16940 25620 16996 27580
rect 17164 27074 17220 27086
rect 17164 27022 17166 27074
rect 17218 27022 17220 27074
rect 17052 26852 17108 26862
rect 17052 26758 17108 26796
rect 16828 25564 16996 25620
rect 17052 25844 17108 25854
rect 16828 25172 16884 25564
rect 17052 25508 17108 25788
rect 17052 25442 17108 25452
rect 16828 25106 16884 25116
rect 16940 25394 16996 25406
rect 16940 25342 16942 25394
rect 16994 25342 16996 25394
rect 16828 24948 16884 24958
rect 16828 24854 16884 24892
rect 16492 24836 16548 24846
rect 16380 24834 16548 24836
rect 16380 24782 16494 24834
rect 16546 24782 16548 24834
rect 16380 24780 16548 24782
rect 16492 24770 16548 24780
rect 16380 23828 16436 23838
rect 16380 23042 16436 23772
rect 16716 23826 16772 23838
rect 16716 23774 16718 23826
rect 16770 23774 16772 23826
rect 16380 22990 16382 23042
rect 16434 22990 16436 23042
rect 16380 22978 16436 22990
rect 16604 23492 16660 23502
rect 16604 23154 16660 23436
rect 16604 23102 16606 23154
rect 16658 23102 16660 23154
rect 16604 22596 16660 23102
rect 16604 22530 16660 22540
rect 16604 22258 16660 22270
rect 16604 22206 16606 22258
rect 16658 22206 16660 22258
rect 16604 21700 16660 22206
rect 16716 21812 16772 23774
rect 16716 21746 16772 21756
rect 16604 21634 16660 21644
rect 16492 21588 16548 21598
rect 16492 21364 16548 21532
rect 16492 21270 16548 21308
rect 16716 21588 16772 21598
rect 16268 19966 16270 20018
rect 16322 19966 16324 20018
rect 16268 19954 16324 19966
rect 16380 19236 16436 19246
rect 16380 19142 16436 19180
rect 16716 19234 16772 21532
rect 16940 21252 16996 25342
rect 17164 24052 17220 27022
rect 17276 26402 17332 27692
rect 17276 26350 17278 26402
rect 17330 26350 17332 26402
rect 17276 26338 17332 26350
rect 17388 27076 17444 28140
rect 17500 27858 17556 28140
rect 17500 27806 17502 27858
rect 17554 27806 17556 27858
rect 17500 27794 17556 27806
rect 17612 27636 17668 29372
rect 17836 29428 17892 29438
rect 17836 29334 17892 29372
rect 18396 29428 18452 30604
rect 18396 29362 18452 29372
rect 18508 30436 18564 30446
rect 18396 29204 18452 29214
rect 18508 29204 18564 30380
rect 18396 29202 18564 29204
rect 18396 29150 18398 29202
rect 18450 29150 18564 29202
rect 18396 29148 18564 29150
rect 18396 29138 18452 29148
rect 18172 28868 18228 28878
rect 18396 28868 18452 28878
rect 18060 28756 18116 28766
rect 18060 28662 18116 28700
rect 18060 28420 18116 28430
rect 17948 28308 18004 28318
rect 17836 28252 17948 28308
rect 17276 26068 17332 26078
rect 17276 24724 17332 26012
rect 17388 24948 17444 27020
rect 17500 27580 17668 27636
rect 17724 27972 17780 27982
rect 17500 26404 17556 27580
rect 17500 25506 17556 26348
rect 17724 27188 17780 27916
rect 17500 25454 17502 25506
rect 17554 25454 17556 25506
rect 17500 25442 17556 25454
rect 17612 26290 17668 26302
rect 17612 26238 17614 26290
rect 17666 26238 17668 26290
rect 17612 25060 17668 26238
rect 17724 25730 17780 27132
rect 17836 26962 17892 28252
rect 17948 28242 18004 28252
rect 17948 27748 18004 27758
rect 18060 27748 18116 28364
rect 17948 27746 18116 27748
rect 17948 27694 17950 27746
rect 18002 27694 18116 27746
rect 17948 27692 18116 27694
rect 17948 27682 18004 27692
rect 18172 27188 18228 28812
rect 18284 28812 18396 28868
rect 18284 28082 18340 28812
rect 18396 28802 18452 28812
rect 18620 28756 18676 32060
rect 18732 32050 18788 32060
rect 18732 30996 18788 31006
rect 18732 30902 18788 30940
rect 18844 30324 18900 33964
rect 18956 33458 19012 34300
rect 19180 34262 19236 34300
rect 19292 34354 19348 34524
rect 19292 34302 19294 34354
rect 19346 34302 19348 34354
rect 19292 34290 19348 34302
rect 19404 34132 19460 34636
rect 19292 34130 19460 34132
rect 19292 34078 19406 34130
rect 19458 34078 19460 34130
rect 19292 34076 19460 34078
rect 18956 33406 18958 33458
rect 19010 33406 19012 33458
rect 18956 33394 19012 33406
rect 19180 33908 19236 33918
rect 18508 28700 18620 28756
rect 18396 28644 18452 28654
rect 18396 28550 18452 28588
rect 18284 28030 18286 28082
rect 18338 28030 18340 28082
rect 18284 28018 18340 28030
rect 18508 28082 18564 28700
rect 18620 28690 18676 28700
rect 18732 30268 18900 30324
rect 19068 33348 19124 33358
rect 18732 29876 18788 30268
rect 18844 30100 18900 30110
rect 18844 30006 18900 30044
rect 19068 29876 19124 33292
rect 19180 32450 19236 33852
rect 19180 32398 19182 32450
rect 19234 32398 19236 32450
rect 19180 32386 19236 32398
rect 19292 33346 19348 34076
rect 19404 34066 19460 34076
rect 19516 34690 19572 34702
rect 19516 34638 19518 34690
rect 19570 34638 19572 34690
rect 19516 33572 19572 34638
rect 19628 33908 19684 35756
rect 19740 34916 19796 35868
rect 20300 35700 20356 36428
rect 20412 36418 20468 36428
rect 20524 36484 20580 36494
rect 20748 36484 20804 36494
rect 20524 36482 20748 36484
rect 20524 36430 20526 36482
rect 20578 36430 20748 36482
rect 20524 36428 20748 36430
rect 20524 36418 20580 36428
rect 20748 36418 20804 36428
rect 20636 36260 20692 36270
rect 20692 36204 20804 36260
rect 20636 36166 20692 36204
rect 20300 35586 20356 35644
rect 20748 35698 20804 36204
rect 20748 35646 20750 35698
rect 20802 35646 20804 35698
rect 20748 35634 20804 35646
rect 20300 35534 20302 35586
rect 20354 35534 20356 35586
rect 20300 35522 20356 35534
rect 20636 35588 20692 35598
rect 20636 35494 20692 35532
rect 20076 34916 20132 34926
rect 20860 34916 20916 36652
rect 21196 36260 21252 37996
rect 21308 37986 21364 37996
rect 21532 37940 21588 37950
rect 21532 37846 21588 37884
rect 21644 37938 21700 37950
rect 21644 37886 21646 37938
rect 21698 37886 21700 37938
rect 21644 37490 21700 37886
rect 21644 37438 21646 37490
rect 21698 37438 21700 37490
rect 21644 37426 21700 37438
rect 21532 37378 21588 37390
rect 21532 37326 21534 37378
rect 21586 37326 21588 37378
rect 21532 37268 21588 37326
rect 21756 37268 21812 38612
rect 21532 37212 21924 37268
rect 21308 36708 21364 36718
rect 21308 36594 21364 36652
rect 21308 36542 21310 36594
rect 21362 36542 21364 36594
rect 21308 36530 21364 36542
rect 21756 36708 21812 36718
rect 21532 36484 21588 36494
rect 21532 36390 21588 36428
rect 21196 36204 21476 36260
rect 21084 35700 21140 35710
rect 21084 35606 21140 35644
rect 21308 35028 21364 35038
rect 19740 34860 19908 34916
rect 19852 34692 19908 34860
rect 19964 34804 20020 34814
rect 19964 34710 20020 34748
rect 20076 34802 20132 34860
rect 20748 34860 20916 34916
rect 20972 35026 21364 35028
rect 20972 34974 21310 35026
rect 21362 34974 21364 35026
rect 20972 34972 21364 34974
rect 20076 34750 20078 34802
rect 20130 34750 20132 34802
rect 20076 34738 20132 34750
rect 20188 34804 20244 34814
rect 19852 34626 19908 34636
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19740 34132 19796 34142
rect 19740 34038 19796 34076
rect 20188 34130 20244 34748
rect 20524 34802 20580 34814
rect 20524 34750 20526 34802
rect 20578 34750 20580 34802
rect 20188 34078 20190 34130
rect 20242 34078 20244 34130
rect 20188 33908 20244 34078
rect 19628 33852 19908 33908
rect 19292 33294 19294 33346
rect 19346 33294 19348 33346
rect 19292 31556 19348 33294
rect 19404 33516 19572 33572
rect 19404 32452 19460 33516
rect 19740 33348 19796 33358
rect 19404 32386 19460 32396
rect 19516 33346 19796 33348
rect 19516 33294 19742 33346
rect 19794 33294 19796 33346
rect 19516 33292 19796 33294
rect 19292 31490 19348 31500
rect 19516 31780 19572 33292
rect 19740 33282 19796 33292
rect 19852 33124 19908 33852
rect 20188 33842 20244 33852
rect 20300 34690 20356 34702
rect 20300 34638 20302 34690
rect 20354 34638 20356 34690
rect 20300 33348 20356 34638
rect 20524 33460 20580 34750
rect 20636 34692 20692 34702
rect 20636 34598 20692 34636
rect 20748 33572 20804 34860
rect 20860 34690 20916 34702
rect 20860 34638 20862 34690
rect 20914 34638 20916 34690
rect 20860 33572 20916 34638
rect 20972 34242 21028 34972
rect 21308 34962 21364 34972
rect 21420 34916 21476 36204
rect 21420 34802 21476 34860
rect 21420 34750 21422 34802
rect 21474 34750 21476 34802
rect 21420 34738 21476 34750
rect 21644 34802 21700 34814
rect 21644 34750 21646 34802
rect 21698 34750 21700 34802
rect 20972 34190 20974 34242
rect 21026 34190 21028 34242
rect 20972 34178 21028 34190
rect 21532 33684 21588 33694
rect 20860 33516 21364 33572
rect 20748 33506 20804 33516
rect 20524 33394 20580 33404
rect 20300 33282 20356 33292
rect 19516 31444 19572 31724
rect 19516 31378 19572 31388
rect 19628 33068 19908 33124
rect 20412 33124 20468 33134
rect 20748 33124 20804 33134
rect 19628 32564 19684 33068
rect 20412 33030 20468 33068
rect 20524 33122 20804 33124
rect 20524 33070 20750 33122
rect 20802 33070 20804 33122
rect 20524 33068 20804 33070
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 20524 32900 20580 33068
rect 20748 33058 20804 33068
rect 19740 32564 19796 32574
rect 19628 32562 19796 32564
rect 19628 32510 19742 32562
rect 19794 32510 19796 32562
rect 19628 32508 19796 32510
rect 19628 30996 19684 32508
rect 19740 32498 19796 32508
rect 20300 31890 20356 31902
rect 20300 31838 20302 31890
rect 20354 31838 20356 31890
rect 20300 31444 20356 31838
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20300 31378 20356 31388
rect 19836 31322 20100 31332
rect 20524 31108 20580 32844
rect 21308 32562 21364 33516
rect 21308 32510 21310 32562
rect 21362 32510 21364 32562
rect 21308 32498 21364 32510
rect 20636 32450 20692 32462
rect 20636 32398 20638 32450
rect 20690 32398 20692 32450
rect 20636 32116 20692 32398
rect 20636 32050 20692 32060
rect 20860 32450 20916 32462
rect 20860 32398 20862 32450
rect 20914 32398 20916 32450
rect 20748 31666 20804 31678
rect 20748 31614 20750 31666
rect 20802 31614 20804 31666
rect 20636 31556 20692 31566
rect 20636 31462 20692 31500
rect 20748 31444 20804 31614
rect 20748 31378 20804 31388
rect 20412 31052 20580 31108
rect 19740 30996 19796 31006
rect 19628 30940 19740 30996
rect 19740 30930 19796 30940
rect 20076 30884 20132 30894
rect 19852 30324 19908 30334
rect 19852 30230 19908 30268
rect 20076 30212 20132 30828
rect 20412 30434 20468 31052
rect 20860 30996 20916 32398
rect 21196 31780 21252 31790
rect 21196 31686 21252 31724
rect 21420 31668 21476 31678
rect 21420 31574 21476 31612
rect 20412 30382 20414 30434
rect 20466 30382 20468 30434
rect 20412 30370 20468 30382
rect 20524 30940 20916 30996
rect 21532 30994 21588 33628
rect 21644 33122 21700 34750
rect 21644 33070 21646 33122
rect 21698 33070 21700 33122
rect 21644 33058 21700 33070
rect 21532 30942 21534 30994
rect 21586 30942 21588 30994
rect 20300 30324 20356 30334
rect 20300 30230 20356 30268
rect 20076 30156 20244 30212
rect 19404 30100 19460 30110
rect 18732 28420 18788 29820
rect 18844 29820 19124 29876
rect 19180 30098 19460 30100
rect 19180 30046 19406 30098
rect 19458 30046 19460 30098
rect 19180 30044 19460 30046
rect 18844 29538 18900 29820
rect 18844 29486 18846 29538
rect 18898 29486 18900 29538
rect 18844 29474 18900 29486
rect 18956 29428 19012 29438
rect 18956 29334 19012 29372
rect 19068 29426 19124 29438
rect 19068 29374 19070 29426
rect 19122 29374 19124 29426
rect 19068 28868 19124 29374
rect 19068 28802 19124 28812
rect 18732 28354 18788 28364
rect 19068 28418 19124 28430
rect 19068 28366 19070 28418
rect 19122 28366 19124 28418
rect 19068 28196 19124 28366
rect 19180 28308 19236 30044
rect 19404 30034 19460 30044
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20188 29764 20244 30156
rect 20188 29708 20356 29764
rect 19852 29426 19908 29438
rect 19852 29374 19854 29426
rect 19906 29374 19908 29426
rect 19852 29316 19908 29374
rect 19852 29250 19908 29260
rect 20188 29426 20244 29438
rect 20188 29374 20190 29426
rect 20242 29374 20244 29426
rect 19180 28242 19236 28252
rect 19292 29204 19348 29214
rect 19068 28130 19124 28140
rect 18508 28030 18510 28082
rect 18562 28030 18564 28082
rect 18508 27748 18564 28030
rect 19068 27972 19124 27982
rect 18620 27860 18676 27870
rect 18620 27766 18676 27804
rect 18844 27860 18900 27870
rect 18508 27682 18564 27692
rect 18172 27122 18228 27132
rect 18396 27186 18452 27198
rect 18396 27134 18398 27186
rect 18450 27134 18452 27186
rect 17836 26910 17838 26962
rect 17890 26910 17892 26962
rect 17836 26068 17892 26910
rect 18060 27074 18116 27086
rect 18060 27022 18062 27074
rect 18114 27022 18116 27074
rect 18060 26908 18116 27022
rect 18396 27076 18452 27134
rect 18508 27076 18564 27086
rect 18396 27020 18508 27076
rect 18508 27010 18564 27020
rect 18844 27076 18900 27804
rect 19068 27746 19124 27916
rect 19068 27694 19070 27746
rect 19122 27694 19124 27746
rect 18844 27010 18900 27020
rect 18956 27074 19012 27086
rect 18956 27022 18958 27074
rect 19010 27022 19012 27074
rect 18060 26852 18452 26908
rect 18396 26740 18452 26852
rect 18396 26684 18564 26740
rect 17836 26002 17892 26012
rect 18396 26516 18452 26526
rect 17724 25678 17726 25730
rect 17778 25678 17780 25730
rect 17724 25666 17780 25678
rect 18172 25506 18228 25518
rect 18172 25454 18174 25506
rect 18226 25454 18228 25506
rect 17836 25172 17892 25182
rect 17612 25004 17780 25060
rect 17500 24948 17556 24958
rect 17388 24946 17556 24948
rect 17388 24894 17502 24946
rect 17554 24894 17556 24946
rect 17388 24892 17556 24894
rect 17500 24882 17556 24892
rect 17612 24834 17668 24846
rect 17612 24782 17614 24834
rect 17666 24782 17668 24834
rect 17500 24724 17556 24734
rect 17276 24668 17500 24724
rect 17500 24630 17556 24668
rect 17164 23986 17220 23996
rect 17612 23828 17668 24782
rect 17612 23762 17668 23772
rect 17388 21924 17444 21934
rect 17724 21924 17780 25004
rect 17836 23154 17892 25116
rect 18172 25060 18228 25454
rect 18284 25284 18340 25294
rect 18284 25190 18340 25228
rect 18284 25060 18340 25070
rect 18172 25004 18284 25060
rect 18284 24994 18340 25004
rect 17836 23102 17838 23154
rect 17890 23102 17892 23154
rect 17836 23090 17892 23102
rect 17948 24836 18004 24846
rect 17948 23042 18004 24780
rect 18284 24836 18340 24846
rect 17948 22990 17950 23042
rect 18002 22990 18004 23042
rect 17948 22978 18004 22990
rect 18172 24612 18228 24622
rect 17724 21868 17892 21924
rect 17388 21810 17444 21868
rect 17388 21758 17390 21810
rect 17442 21758 17444 21810
rect 17388 21746 17444 21758
rect 17500 21812 17556 21822
rect 17500 21718 17556 21756
rect 16940 21186 16996 21196
rect 17612 21698 17668 21710
rect 17612 21646 17614 21698
rect 17666 21646 17668 21698
rect 16940 20692 16996 20702
rect 16828 20018 16884 20030
rect 16828 19966 16830 20018
rect 16882 19966 16884 20018
rect 16828 19796 16884 19966
rect 16828 19730 16884 19740
rect 16940 19236 16996 20636
rect 17500 20468 17556 20478
rect 17388 20018 17444 20030
rect 17388 19966 17390 20018
rect 17442 19966 17444 20018
rect 17388 19572 17444 19966
rect 17388 19506 17444 19516
rect 17500 19460 17556 20412
rect 17500 19394 17556 19404
rect 17164 19348 17220 19358
rect 17164 19254 17220 19292
rect 16716 19182 16718 19234
rect 16770 19182 16772 19234
rect 16716 19170 16772 19182
rect 16828 19234 16996 19236
rect 16828 19182 16942 19234
rect 16994 19182 16996 19234
rect 16828 19180 16996 19182
rect 16492 19012 16548 19022
rect 16492 18918 16548 18956
rect 16156 17714 16212 17724
rect 16716 18340 16772 18350
rect 16828 18340 16884 19180
rect 16940 19170 16996 19180
rect 17052 19236 17108 19246
rect 17052 19012 17108 19180
rect 17052 18956 17220 19012
rect 16716 18338 16884 18340
rect 16716 18286 16718 18338
rect 16770 18286 16884 18338
rect 16716 18284 16884 18286
rect 16716 17556 16772 18284
rect 16716 17490 16772 17500
rect 17052 17666 17108 17678
rect 17052 17614 17054 17666
rect 17106 17614 17108 17666
rect 16940 17444 16996 17454
rect 16828 17442 16996 17444
rect 16828 17390 16942 17442
rect 16994 17390 16996 17442
rect 16828 17388 16996 17390
rect 16044 16996 16100 17006
rect 16044 16098 16100 16940
rect 16044 16046 16046 16098
rect 16098 16046 16100 16098
rect 16044 16034 16100 16046
rect 16156 16884 16212 16894
rect 15932 15820 16100 15876
rect 15820 15316 15876 15326
rect 15820 15222 15876 15260
rect 15932 15204 15988 15214
rect 15708 14478 15710 14530
rect 15762 14478 15764 14530
rect 15708 14466 15764 14478
rect 15820 15092 15988 15148
rect 15708 13972 15764 13982
rect 15708 13746 15764 13916
rect 15708 13694 15710 13746
rect 15762 13694 15764 13746
rect 15708 13682 15764 13694
rect 15484 12348 15652 12404
rect 15260 11442 15316 11452
rect 15372 12292 15428 12302
rect 15372 12178 15428 12236
rect 15372 12126 15374 12178
rect 15426 12126 15428 12178
rect 15372 11284 15428 12126
rect 15260 11228 15428 11284
rect 15260 11172 15316 11228
rect 15484 11172 15540 12348
rect 15708 12292 15764 12302
rect 15596 12236 15708 12292
rect 15596 12178 15652 12236
rect 15708 12226 15764 12236
rect 15596 12126 15598 12178
rect 15650 12126 15652 12178
rect 15596 12114 15652 12126
rect 15036 10782 15038 10834
rect 15090 10782 15092 10834
rect 15036 10770 15092 10782
rect 15148 11116 15316 11172
rect 15372 11116 15540 11172
rect 14924 10670 14926 10722
rect 14978 10670 14980 10722
rect 14924 10658 14980 10670
rect 14812 9884 14980 9940
rect 14812 9716 14868 9726
rect 14700 9660 14812 9716
rect 14700 9268 14756 9660
rect 14812 9622 14868 9660
rect 14924 9268 14980 9884
rect 15148 9716 15204 11116
rect 15148 9650 15204 9660
rect 15260 10612 15316 10622
rect 14700 9202 14756 9212
rect 14812 9212 14980 9268
rect 15260 9268 15316 10556
rect 15372 9940 15428 11116
rect 15484 10722 15540 10734
rect 15484 10670 15486 10722
rect 15538 10670 15540 10722
rect 15484 10612 15540 10670
rect 15596 10612 15652 10622
rect 15484 10556 15596 10612
rect 15820 10612 15876 15092
rect 15932 13858 15988 13870
rect 15932 13806 15934 13858
rect 15986 13806 15988 13858
rect 15932 12404 15988 13806
rect 15932 12338 15988 12348
rect 16044 10834 16100 15820
rect 16044 10782 16046 10834
rect 16098 10782 16100 10834
rect 16044 10770 16100 10782
rect 15820 10556 16100 10612
rect 15596 10546 15652 10556
rect 15932 10052 15988 10062
rect 15372 9938 15652 9940
rect 15372 9886 15374 9938
rect 15426 9886 15652 9938
rect 15372 9884 15652 9886
rect 15372 9874 15428 9884
rect 15260 9212 15428 9268
rect 14700 9044 14756 9054
rect 14700 8950 14756 8988
rect 14812 8484 14868 9212
rect 15036 9154 15092 9166
rect 15036 9102 15038 9154
rect 15090 9102 15092 9154
rect 14924 9042 14980 9054
rect 14924 8990 14926 9042
rect 14978 8990 14980 9042
rect 14924 8596 14980 8990
rect 14924 8530 14980 8540
rect 14812 8418 14868 8428
rect 15036 8260 15092 9102
rect 15260 9044 15316 9054
rect 15260 8950 15316 8988
rect 14812 7588 14868 7598
rect 14812 7586 14980 7588
rect 14812 7534 14814 7586
rect 14866 7534 14980 7586
rect 14812 7532 14980 7534
rect 14812 7522 14868 7532
rect 14588 7308 14868 7364
rect 14252 7298 14308 7308
rect 14140 6802 14196 6814
rect 14140 6750 14142 6802
rect 14194 6750 14196 6802
rect 13692 6690 13748 6702
rect 13692 6638 13694 6690
rect 13746 6638 13748 6690
rect 13468 6468 13524 6478
rect 13468 6374 13524 6412
rect 13692 6244 13748 6638
rect 14140 6692 14196 6750
rect 14140 6626 14196 6636
rect 13692 6178 13748 6188
rect 13916 6468 13972 6478
rect 13468 6132 13524 6142
rect 13468 6038 13524 6076
rect 13132 5906 13188 5964
rect 13692 6020 13748 6030
rect 13692 5926 13748 5964
rect 13132 5854 13134 5906
rect 13186 5854 13188 5906
rect 13132 5842 13188 5854
rect 13580 5794 13636 5806
rect 13580 5742 13582 5794
rect 13634 5742 13636 5794
rect 13468 5348 13524 5358
rect 13580 5348 13636 5742
rect 13916 5460 13972 6412
rect 14588 6356 14644 6366
rect 14364 6244 14420 6254
rect 14140 5908 14196 5918
rect 14140 5814 14196 5852
rect 14252 5906 14308 5918
rect 14252 5854 14254 5906
rect 14306 5854 14308 5906
rect 14252 5460 14308 5854
rect 14364 5572 14420 6188
rect 14476 6132 14532 6142
rect 14476 6038 14532 6076
rect 14364 5506 14420 5516
rect 13916 5404 14196 5460
rect 13468 5346 13636 5348
rect 13468 5294 13470 5346
rect 13522 5294 13636 5346
rect 13468 5292 13636 5294
rect 13468 5282 13524 5292
rect 14028 5236 14084 5246
rect 13580 5124 13636 5134
rect 13580 5030 13636 5068
rect 13804 5012 13860 5022
rect 13804 4918 13860 4956
rect 13020 4386 13076 4396
rect 13244 4900 13300 4910
rect 12796 4228 12852 4238
rect 12796 4226 13188 4228
rect 12796 4174 12798 4226
rect 12850 4174 13188 4226
rect 12796 4172 13188 4174
rect 12796 4162 12852 4172
rect 12684 3948 12852 4004
rect 12236 3614 12238 3666
rect 12290 3614 12292 3666
rect 11340 3602 11396 3612
rect 12236 3602 12292 3614
rect 10892 3444 10948 3482
rect 10892 3378 10948 3388
rect 11788 3444 11844 3482
rect 11788 3378 11844 3388
rect 12684 3444 12740 3482
rect 12684 3378 12740 3388
rect 12796 1652 12852 3948
rect 13132 3778 13188 4172
rect 13132 3726 13134 3778
rect 13186 3726 13188 3778
rect 13132 3714 13188 3726
rect 13244 3666 13300 4844
rect 13244 3614 13246 3666
rect 13298 3614 13300 3666
rect 13244 3602 13300 3614
rect 13580 4564 13636 4574
rect 13580 4338 13636 4508
rect 13580 4286 13582 4338
rect 13634 4286 13636 4338
rect 13580 3668 13636 4286
rect 13916 4228 13972 4238
rect 14028 4228 14084 5180
rect 14140 5010 14196 5404
rect 14252 5394 14308 5404
rect 14364 5348 14420 5358
rect 14364 5122 14420 5292
rect 14364 5070 14366 5122
rect 14418 5070 14420 5122
rect 14364 5058 14420 5070
rect 14140 4958 14142 5010
rect 14194 4958 14196 5010
rect 14140 4946 14196 4958
rect 14252 4900 14308 4910
rect 14252 4806 14308 4844
rect 13916 4226 14084 4228
rect 13916 4174 13918 4226
rect 13970 4174 14084 4226
rect 13916 4172 14084 4174
rect 14140 4228 14196 4238
rect 13916 4162 13972 4172
rect 13580 3602 13636 3612
rect 14140 3666 14196 4172
rect 14140 3614 14142 3666
rect 14194 3614 14196 3666
rect 14140 3602 14196 3614
rect 14588 3666 14644 6300
rect 14700 5908 14756 5918
rect 14700 5814 14756 5852
rect 14588 3614 14590 3666
rect 14642 3614 14644 3666
rect 14588 3602 14644 3614
rect 14812 3668 14868 7308
rect 14924 6244 14980 7532
rect 14924 6178 14980 6188
rect 14924 5906 14980 5918
rect 14924 5854 14926 5906
rect 14978 5854 14980 5906
rect 14924 5348 14980 5854
rect 14924 5282 14980 5292
rect 15036 5124 15092 8204
rect 14924 5068 15092 5124
rect 15148 8484 15204 8494
rect 15148 7698 15204 8428
rect 15148 7646 15150 7698
rect 15202 7646 15204 7698
rect 14924 4676 14980 5068
rect 14924 4610 14980 4620
rect 15036 4898 15092 4910
rect 15036 4846 15038 4898
rect 15090 4846 15092 4898
rect 15036 4564 15092 4846
rect 15036 4498 15092 4508
rect 15148 3892 15204 7646
rect 15036 3668 15092 3678
rect 14812 3666 15092 3668
rect 14812 3614 15038 3666
rect 15090 3614 15092 3666
rect 14812 3612 15092 3614
rect 15036 3602 15092 3612
rect 15148 3444 15204 3836
rect 12796 1586 12852 1596
rect 15036 3388 15204 3444
rect 15260 5124 15316 5134
rect 15260 3444 15316 5068
rect 15372 4564 15428 9212
rect 15596 8820 15652 9884
rect 15708 9828 15764 9838
rect 15708 9734 15764 9772
rect 15820 8820 15876 8830
rect 15596 8818 15876 8820
rect 15596 8766 15822 8818
rect 15874 8766 15876 8818
rect 15596 8764 15876 8766
rect 15820 8754 15876 8764
rect 15932 8596 15988 9996
rect 16044 9940 16100 10556
rect 16044 9266 16100 9884
rect 16044 9214 16046 9266
rect 16098 9214 16100 9266
rect 16044 9202 16100 9214
rect 15708 8540 15988 8596
rect 15596 8148 15652 8158
rect 15596 8054 15652 8092
rect 15484 5908 15540 5918
rect 15484 5814 15540 5852
rect 15596 5908 15652 5918
rect 15708 5908 15764 8540
rect 15932 8036 15988 8046
rect 15932 7698 15988 7980
rect 15932 7646 15934 7698
rect 15986 7646 15988 7698
rect 15932 7634 15988 7646
rect 16156 7700 16212 16828
rect 16492 16324 16548 16334
rect 16492 16230 16548 16268
rect 16604 16212 16660 16222
rect 16380 15986 16436 15998
rect 16380 15934 16382 15986
rect 16434 15934 16436 15986
rect 16380 15764 16436 15934
rect 16492 15988 16548 15998
rect 16604 15988 16660 16156
rect 16492 15986 16660 15988
rect 16492 15934 16494 15986
rect 16546 15934 16660 15986
rect 16492 15932 16660 15934
rect 16716 15988 16772 15998
rect 16492 15922 16548 15932
rect 16380 15708 16548 15764
rect 16268 15540 16324 15550
rect 16268 15446 16324 15484
rect 16492 15204 16548 15708
rect 16492 15138 16548 15148
rect 16716 15202 16772 15932
rect 16828 15876 16884 17388
rect 16940 17378 16996 17388
rect 17052 16098 17108 17614
rect 17052 16046 17054 16098
rect 17106 16046 17108 16098
rect 16828 15820 16996 15876
rect 16716 15150 16718 15202
rect 16770 15150 16772 15202
rect 16492 14756 16548 14766
rect 16492 14662 16548 14700
rect 16604 14532 16660 14542
rect 16604 14438 16660 14476
rect 16492 14308 16548 14318
rect 16268 13860 16324 13870
rect 16268 13766 16324 13804
rect 16492 13748 16548 14252
rect 16604 14196 16660 14206
rect 16604 13858 16660 14140
rect 16604 13806 16606 13858
rect 16658 13806 16660 13858
rect 16604 13794 16660 13806
rect 16492 13682 16548 13692
rect 16380 13634 16436 13646
rect 16380 13582 16382 13634
rect 16434 13582 16436 13634
rect 16380 13076 16436 13582
rect 16716 13412 16772 15150
rect 16940 14530 16996 15820
rect 17052 15652 17108 16046
rect 17052 15316 17108 15596
rect 17052 15250 17108 15260
rect 17164 15148 17220 18956
rect 17500 19010 17556 19022
rect 17500 18958 17502 19010
rect 17554 18958 17556 19010
rect 17388 18676 17444 18686
rect 17388 18452 17444 18620
rect 17388 18386 17444 18396
rect 17388 18228 17444 18238
rect 17276 18172 17388 18228
rect 17276 17108 17332 18172
rect 17388 18162 17444 18172
rect 17388 18004 17444 18014
rect 17388 17666 17444 17948
rect 17388 17614 17390 17666
rect 17442 17614 17444 17666
rect 17388 17602 17444 17614
rect 17388 17108 17444 17118
rect 17332 17106 17444 17108
rect 17332 17054 17390 17106
rect 17442 17054 17444 17106
rect 17332 17052 17444 17054
rect 17276 17014 17332 17052
rect 17388 17042 17444 17052
rect 17500 17108 17556 18958
rect 17612 18788 17668 21646
rect 17724 21698 17780 21710
rect 17724 21646 17726 21698
rect 17778 21646 17780 21698
rect 17724 20356 17780 21646
rect 17836 21364 17892 21868
rect 17836 21298 17892 21308
rect 17948 21812 18004 21822
rect 17948 21252 18004 21756
rect 17948 21186 18004 21196
rect 18060 21586 18116 21598
rect 18060 21534 18062 21586
rect 18114 21534 18116 21586
rect 18060 20804 18116 21534
rect 18172 21476 18228 24556
rect 18284 21588 18340 24780
rect 18396 23266 18452 26460
rect 18396 23214 18398 23266
rect 18450 23214 18452 23266
rect 18396 23202 18452 23214
rect 18508 21924 18564 26684
rect 18956 25172 19012 27022
rect 19068 26852 19124 27694
rect 19180 27188 19236 27198
rect 19180 27074 19236 27132
rect 19180 27022 19182 27074
rect 19234 27022 19236 27074
rect 19180 27010 19236 27022
rect 19068 26796 19236 26852
rect 19068 26628 19124 26638
rect 19068 26290 19124 26572
rect 19068 26238 19070 26290
rect 19122 26238 19124 26290
rect 19068 25396 19124 26238
rect 19180 26068 19236 26796
rect 19180 26002 19236 26012
rect 19180 25396 19236 25406
rect 19068 25394 19236 25396
rect 19068 25342 19182 25394
rect 19234 25342 19236 25394
rect 19068 25340 19236 25342
rect 19180 25330 19236 25340
rect 18732 25116 19012 25172
rect 18620 25060 18676 25070
rect 18620 23828 18676 25004
rect 18620 23762 18676 23772
rect 18732 22484 18788 25116
rect 18956 24892 19236 24948
rect 18844 24836 18900 24846
rect 18844 24050 18900 24780
rect 18956 24834 19012 24892
rect 18956 24782 18958 24834
rect 19010 24782 19012 24834
rect 18956 24770 19012 24782
rect 19068 24722 19124 24734
rect 19068 24670 19070 24722
rect 19122 24670 19124 24722
rect 18956 24500 19012 24510
rect 18956 24406 19012 24444
rect 18844 23998 18846 24050
rect 18898 23998 18900 24050
rect 18844 23548 18900 23998
rect 19068 24052 19124 24670
rect 18844 23492 19012 23548
rect 18844 23154 18900 23166
rect 18844 23102 18846 23154
rect 18898 23102 18900 23154
rect 18844 22932 18900 23102
rect 18844 22866 18900 22876
rect 18396 21868 18564 21924
rect 18620 22428 18732 22484
rect 18396 21810 18452 21868
rect 18396 21758 18398 21810
rect 18450 21758 18452 21810
rect 18396 21746 18452 21758
rect 18508 21698 18564 21710
rect 18508 21646 18510 21698
rect 18562 21646 18564 21698
rect 18508 21588 18564 21646
rect 18284 21532 18564 21588
rect 18620 21588 18676 22428
rect 18732 22390 18788 22428
rect 18956 22372 19012 23492
rect 19068 23044 19124 23996
rect 19180 23492 19236 24892
rect 19180 23426 19236 23436
rect 19068 22978 19124 22988
rect 19292 22932 19348 29148
rect 19516 29092 19572 29102
rect 19404 28532 19460 28542
rect 19404 28438 19460 28476
rect 19516 28308 19572 29036
rect 20188 29092 20244 29374
rect 20300 29204 20356 29708
rect 20300 29138 20356 29148
rect 20412 29540 20468 29550
rect 20412 29314 20468 29484
rect 20412 29262 20414 29314
rect 20466 29262 20468 29314
rect 20188 29026 20244 29036
rect 19964 28756 20020 28766
rect 19964 28662 20020 28700
rect 20076 28532 20132 28542
rect 20300 28532 20356 28542
rect 20132 28530 20356 28532
rect 20132 28478 20302 28530
rect 20354 28478 20356 28530
rect 20132 28476 20356 28478
rect 20076 28466 20132 28476
rect 20300 28466 20356 28476
rect 19404 28252 19572 28308
rect 19836 28252 20100 28262
rect 19404 26516 19460 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19516 27858 19572 27870
rect 19516 27806 19518 27858
rect 19570 27806 19572 27858
rect 19516 26908 19572 27806
rect 19852 27468 20244 27524
rect 19852 27074 19908 27468
rect 19852 27022 19854 27074
rect 19906 27022 19908 27074
rect 19852 27010 19908 27022
rect 19964 27186 20020 27198
rect 19964 27134 19966 27186
rect 20018 27134 20020 27186
rect 19516 26852 19684 26908
rect 19628 26516 19684 26852
rect 19964 26852 20020 27134
rect 20076 27076 20132 27114
rect 20188 27076 20244 27468
rect 20412 27298 20468 29262
rect 20524 28644 20580 30940
rect 21196 30884 21252 30894
rect 20748 30882 21252 30884
rect 20748 30830 21198 30882
rect 21250 30830 21252 30882
rect 20748 30828 21252 30830
rect 20748 30434 20804 30828
rect 21196 30818 21252 30828
rect 21532 30772 21588 30942
rect 21532 30706 21588 30716
rect 21644 32452 21700 32462
rect 21644 31666 21700 32396
rect 21644 31614 21646 31666
rect 21698 31614 21700 31666
rect 21644 30660 21700 31614
rect 21644 30594 21700 30604
rect 21756 30436 21812 36652
rect 21868 36706 21924 37212
rect 21868 36654 21870 36706
rect 21922 36654 21924 36706
rect 21868 36642 21924 36654
rect 21980 34916 22036 34926
rect 21980 34802 22036 34860
rect 21980 34750 21982 34802
rect 22034 34750 22036 34802
rect 21980 34738 22036 34750
rect 22092 34580 22148 41132
rect 22316 40964 22372 40974
rect 22316 40852 22372 40908
rect 22316 40796 22596 40852
rect 22204 39844 22260 39854
rect 22204 39506 22260 39788
rect 22316 39620 22372 39630
rect 22316 39526 22372 39564
rect 22204 39454 22206 39506
rect 22258 39454 22260 39506
rect 22204 39442 22260 39454
rect 22428 39508 22484 39518
rect 22428 39172 22484 39452
rect 22316 39116 22484 39172
rect 22316 38946 22372 39116
rect 22316 38894 22318 38946
rect 22370 38894 22372 38946
rect 22204 38836 22260 38846
rect 22204 37940 22260 38780
rect 22316 38724 22372 38894
rect 22428 38948 22484 38958
rect 22428 38854 22484 38892
rect 22316 38658 22372 38668
rect 22316 37940 22372 37950
rect 22204 37938 22372 37940
rect 22204 37886 22318 37938
rect 22370 37886 22372 37938
rect 22204 37884 22372 37886
rect 22316 37874 22372 37884
rect 22316 37156 22372 37166
rect 22540 37156 22596 40796
rect 23324 40628 23380 41246
rect 23996 41300 24052 43372
rect 24332 43426 24388 43484
rect 24332 43374 24334 43426
rect 24386 43374 24388 43426
rect 24332 43362 24388 43374
rect 24444 42980 24500 43708
rect 24556 43698 24612 43708
rect 24668 45106 24724 45118
rect 24668 45054 24670 45106
rect 24722 45054 24724 45106
rect 24668 43540 24724 45054
rect 25228 44100 25284 44110
rect 25340 44100 25396 45164
rect 25452 45154 25508 45164
rect 25564 45106 25620 45118
rect 25564 45054 25566 45106
rect 25618 45054 25620 45106
rect 25452 44882 25508 44894
rect 25452 44830 25454 44882
rect 25506 44830 25508 44882
rect 25452 44322 25508 44830
rect 25452 44270 25454 44322
rect 25506 44270 25508 44322
rect 25452 44258 25508 44270
rect 25284 44044 25396 44100
rect 25228 43762 25284 44044
rect 25228 43710 25230 43762
rect 25282 43710 25284 43762
rect 25228 43698 25284 43710
rect 25116 43652 25172 43662
rect 25564 43652 25620 45054
rect 26348 45108 26404 45146
rect 26348 45042 26404 45052
rect 27468 45108 27524 45118
rect 26124 44996 26180 45006
rect 26124 44902 26180 44940
rect 27132 44994 27188 45006
rect 27132 44942 27134 44994
rect 27186 44942 27188 44994
rect 26012 44882 26068 44894
rect 26012 44830 26014 44882
rect 26066 44830 26068 44882
rect 26012 44434 26068 44830
rect 26012 44382 26014 44434
rect 26066 44382 26068 44434
rect 26012 44370 26068 44382
rect 26908 44324 26964 44334
rect 26460 44100 26516 44110
rect 26908 44100 26964 44268
rect 26460 44098 26964 44100
rect 26460 44046 26462 44098
rect 26514 44046 26964 44098
rect 26460 44044 26964 44046
rect 27132 44322 27188 44942
rect 27132 44270 27134 44322
rect 27186 44270 27188 44322
rect 27132 44212 27188 44270
rect 25676 43652 25732 43662
rect 25564 43596 25676 43652
rect 25116 43558 25172 43596
rect 25676 43558 25732 43596
rect 24668 43474 24724 43484
rect 25452 43540 25508 43550
rect 25452 43446 25508 43484
rect 26460 43538 26516 44044
rect 27132 43764 27188 44156
rect 26684 43708 27188 43764
rect 27468 43876 27524 45052
rect 29932 45106 29988 45118
rect 29932 45054 29934 45106
rect 29986 45054 29988 45106
rect 29260 44994 29316 45006
rect 29260 44942 29262 44994
rect 29314 44942 29316 44994
rect 28364 44324 28420 44334
rect 28364 44230 28420 44268
rect 26572 43652 26628 43662
rect 26572 43558 26628 43596
rect 26684 43650 26740 43708
rect 26684 43598 26686 43650
rect 26738 43598 26740 43650
rect 26684 43586 26740 43598
rect 27468 43650 27524 43820
rect 27468 43598 27470 43650
rect 27522 43598 27524 43650
rect 27468 43586 27524 43598
rect 27804 44210 27860 44222
rect 27804 44158 27806 44210
rect 27858 44158 27860 44210
rect 27804 43762 27860 44158
rect 28252 44212 28308 44222
rect 28252 44118 28308 44156
rect 28028 44100 28084 44110
rect 28028 44006 28084 44044
rect 28364 43876 28420 43886
rect 28252 43764 28308 43774
rect 27804 43710 27806 43762
rect 27858 43710 27860 43762
rect 26460 43486 26462 43538
rect 26514 43486 26516 43538
rect 26124 43428 26180 43438
rect 26460 43428 26516 43486
rect 23996 41234 24052 41244
rect 24108 42924 24500 42980
rect 26012 43426 26516 43428
rect 26012 43374 26126 43426
rect 26178 43374 26516 43426
rect 26012 43372 26516 43374
rect 27020 43538 27076 43550
rect 27020 43486 27022 43538
rect 27074 43486 27076 43538
rect 23884 41076 23940 41086
rect 23884 40982 23940 41020
rect 24108 41074 24164 42924
rect 24332 42642 24388 42654
rect 24332 42590 24334 42642
rect 24386 42590 24388 42642
rect 24220 41970 24276 41982
rect 24220 41918 24222 41970
rect 24274 41918 24276 41970
rect 24220 41300 24276 41918
rect 24332 41748 24388 42590
rect 25340 42644 25396 42654
rect 25340 42550 25396 42588
rect 25788 42644 25844 42654
rect 26012 42644 26068 43372
rect 26124 43362 26180 43372
rect 27020 43092 27076 43486
rect 26684 43036 27076 43092
rect 26460 42756 26516 42766
rect 26684 42756 26740 43036
rect 26460 42754 26684 42756
rect 26460 42702 26462 42754
rect 26514 42702 26684 42754
rect 26460 42700 26684 42702
rect 26460 42690 26516 42700
rect 26684 42690 26740 42700
rect 27692 42756 27748 42766
rect 27804 42756 27860 43710
rect 27916 43708 28196 43764
rect 27916 43650 27972 43708
rect 27916 43598 27918 43650
rect 27970 43598 27972 43650
rect 27916 43586 27972 43598
rect 28028 43538 28084 43550
rect 28028 43486 28030 43538
rect 28082 43486 28084 43538
rect 27692 42754 27860 42756
rect 27692 42702 27694 42754
rect 27746 42702 27860 42754
rect 27692 42700 27860 42702
rect 27916 42756 27972 42766
rect 28028 42756 28084 43486
rect 27972 42700 28084 42756
rect 28140 42754 28196 43708
rect 28140 42702 28142 42754
rect 28194 42702 28196 42754
rect 27692 42690 27748 42700
rect 27916 42662 27972 42700
rect 28140 42690 28196 42702
rect 25844 42588 26068 42644
rect 26124 42644 26180 42654
rect 25788 42550 25844 42588
rect 26124 42550 26180 42588
rect 26796 42644 26852 42654
rect 26796 42550 26852 42588
rect 24332 41682 24388 41692
rect 24444 42530 24500 42542
rect 24444 42478 24446 42530
rect 24498 42478 24500 42530
rect 24444 41300 24500 42478
rect 24668 42532 24724 42542
rect 25228 42532 25284 42542
rect 24668 42530 25172 42532
rect 24668 42478 24670 42530
rect 24722 42478 25172 42530
rect 24668 42476 25172 42478
rect 24668 42466 24724 42476
rect 25116 42084 25172 42476
rect 25228 42438 25284 42476
rect 26236 42532 26292 42542
rect 26236 42530 26404 42532
rect 26236 42478 26238 42530
rect 26290 42478 26404 42530
rect 26236 42476 26404 42478
rect 26236 42466 26292 42476
rect 26236 42308 26292 42318
rect 26124 42252 26236 42308
rect 25228 42084 25284 42094
rect 25116 42082 25284 42084
rect 25116 42030 25230 42082
rect 25282 42030 25284 42082
rect 25116 42028 25284 42030
rect 25228 42018 25284 42028
rect 25340 42082 25396 42094
rect 25340 42030 25342 42082
rect 25394 42030 25396 42082
rect 24668 41972 24724 41982
rect 24668 41878 24724 41916
rect 25340 41860 25396 42030
rect 26124 42082 26180 42252
rect 26236 42242 26292 42252
rect 26348 42196 26404 42476
rect 26684 42530 26740 42542
rect 26684 42478 26686 42530
rect 26738 42478 26740 42530
rect 26684 42308 26740 42478
rect 26684 42242 26740 42252
rect 26908 42530 26964 42542
rect 26908 42478 26910 42530
rect 26962 42478 26964 42530
rect 26460 42196 26516 42206
rect 26348 42194 26516 42196
rect 26348 42142 26462 42194
rect 26514 42142 26516 42194
rect 26348 42140 26516 42142
rect 26460 42130 26516 42140
rect 26124 42030 26126 42082
rect 26178 42030 26180 42082
rect 25116 41804 25396 41860
rect 25564 41970 25620 41982
rect 25564 41918 25566 41970
rect 25618 41918 25620 41970
rect 24220 41244 24612 41300
rect 24108 41022 24110 41074
rect 24162 41022 24164 41074
rect 24108 40964 24164 41022
rect 24444 40964 24500 40974
rect 24108 40898 24164 40908
rect 24220 40962 24500 40964
rect 24220 40910 24446 40962
rect 24498 40910 24500 40962
rect 24220 40908 24500 40910
rect 23324 40562 23380 40572
rect 22988 40516 23044 40526
rect 22988 40402 23044 40460
rect 22988 40350 22990 40402
rect 23042 40350 23044 40402
rect 22876 39732 22932 39742
rect 22876 39620 22932 39676
rect 22764 39618 22932 39620
rect 22764 39566 22878 39618
rect 22930 39566 22932 39618
rect 22764 39564 22932 39566
rect 22652 39508 22708 39518
rect 22652 39058 22708 39452
rect 22652 39006 22654 39058
rect 22706 39006 22708 39058
rect 22652 38994 22708 39006
rect 22652 37828 22708 37838
rect 22652 37734 22708 37772
rect 22316 37154 22596 37156
rect 22316 37102 22318 37154
rect 22370 37102 22596 37154
rect 22316 37100 22596 37102
rect 22204 36482 22260 36494
rect 22204 36430 22206 36482
rect 22258 36430 22260 36482
rect 22204 36260 22260 36430
rect 22204 36194 22260 36204
rect 22316 35588 22372 37100
rect 22764 36708 22820 39564
rect 22876 39554 22932 39564
rect 22988 39620 23044 40350
rect 23100 40514 23156 40526
rect 23100 40462 23102 40514
rect 23154 40462 23156 40514
rect 23100 39844 23156 40462
rect 24108 40514 24164 40526
rect 24108 40462 24110 40514
rect 24162 40462 24164 40514
rect 24108 40292 24164 40462
rect 24108 40226 24164 40236
rect 23100 39778 23156 39788
rect 22988 39508 23044 39564
rect 24108 39620 24164 39630
rect 24220 39620 24276 40908
rect 24444 40898 24500 40908
rect 24108 39618 24276 39620
rect 24108 39566 24110 39618
rect 24162 39566 24276 39618
rect 24108 39564 24276 39566
rect 24108 39554 24164 39564
rect 23212 39508 23268 39518
rect 22988 39506 23268 39508
rect 22988 39454 23214 39506
rect 23266 39454 23268 39506
rect 22988 39452 23268 39454
rect 23212 39442 23268 39452
rect 23212 39060 23268 39070
rect 23212 38966 23268 39004
rect 22988 38946 23044 38958
rect 22988 38894 22990 38946
rect 23042 38894 23044 38946
rect 22876 38836 22932 38846
rect 22876 38742 22932 38780
rect 22988 38612 23044 38894
rect 23660 38948 23716 38958
rect 23660 38834 23716 38892
rect 23660 38782 23662 38834
rect 23714 38782 23716 38834
rect 23660 38668 23716 38782
rect 24108 38724 24164 38762
rect 23660 38612 24052 38668
rect 24108 38658 24164 38668
rect 22988 38546 23044 38556
rect 23996 38162 24052 38612
rect 23996 38110 23998 38162
rect 24050 38110 24052 38162
rect 23996 38098 24052 38110
rect 24220 38164 24276 39564
rect 24220 38098 24276 38108
rect 24444 40402 24500 40414
rect 24444 40350 24446 40402
rect 24498 40350 24500 40402
rect 24444 39618 24500 40350
rect 24556 39730 24612 41244
rect 25116 41186 25172 41804
rect 25564 41636 25620 41918
rect 25564 41570 25620 41580
rect 26124 41300 26180 42030
rect 26236 42082 26292 42094
rect 26908 42084 26964 42478
rect 26236 42030 26238 42082
rect 26290 42030 26292 42082
rect 26236 41972 26292 42030
rect 26684 42028 26964 42084
rect 27132 42530 27188 42542
rect 27132 42478 27134 42530
rect 27186 42478 27188 42530
rect 26684 41972 26740 42028
rect 26236 41916 26740 41972
rect 26684 41858 26740 41916
rect 26684 41806 26686 41858
rect 26738 41806 26740 41858
rect 26236 41300 26292 41310
rect 26124 41298 26292 41300
rect 26124 41246 26238 41298
rect 26290 41246 26292 41298
rect 26124 41244 26292 41246
rect 25116 41134 25118 41186
rect 25170 41134 25172 41186
rect 25116 41122 25172 41134
rect 24780 41074 24836 41086
rect 24780 41022 24782 41074
rect 24834 41022 24836 41074
rect 24780 40292 24836 41022
rect 24892 40964 24948 40974
rect 24892 40870 24948 40908
rect 25788 40964 25844 40974
rect 25788 40870 25844 40908
rect 25340 40628 25396 40638
rect 25116 40292 25172 40302
rect 24780 40226 24836 40236
rect 25004 40236 25116 40292
rect 25004 39842 25060 40236
rect 25116 40226 25172 40236
rect 25004 39790 25006 39842
rect 25058 39790 25060 39842
rect 25004 39778 25060 39790
rect 24556 39678 24558 39730
rect 24610 39678 24612 39730
rect 24556 39666 24612 39678
rect 24444 39566 24446 39618
rect 24498 39566 24500 39618
rect 23548 38052 23604 38062
rect 23212 37266 23268 37278
rect 23212 37214 23214 37266
rect 23266 37214 23268 37266
rect 22764 36642 22820 36652
rect 22988 37154 23044 37166
rect 22988 37102 22990 37154
rect 23042 37102 23044 37154
rect 22428 36482 22484 36494
rect 22428 36430 22430 36482
rect 22482 36430 22484 36482
rect 22428 35924 22484 36430
rect 22764 36484 22820 36494
rect 22988 36484 23044 37102
rect 23100 36484 23156 36494
rect 22988 36482 23156 36484
rect 22988 36430 23102 36482
rect 23154 36430 23156 36482
rect 22988 36428 23156 36430
rect 22764 36390 22820 36428
rect 22428 35858 22484 35868
rect 22652 36260 22708 36270
rect 22204 35532 22372 35588
rect 22204 34804 22260 35532
rect 22316 35028 22372 35038
rect 22316 34914 22372 34972
rect 22316 34862 22318 34914
rect 22370 34862 22372 34914
rect 22316 34850 22372 34862
rect 22204 34738 22260 34748
rect 22652 34802 22708 36204
rect 23100 36036 23156 36428
rect 23212 36372 23268 37214
rect 23548 36372 23604 37996
rect 23884 38050 23940 38062
rect 23884 37998 23886 38050
rect 23938 37998 23940 38050
rect 23884 37828 23940 37998
rect 24332 38052 24388 38062
rect 24332 37958 24388 37996
rect 23772 37604 23828 37614
rect 23772 37378 23828 37548
rect 23772 37326 23774 37378
rect 23826 37326 23828 37378
rect 23772 37314 23828 37326
rect 23772 36596 23828 36606
rect 23772 36502 23828 36540
rect 23212 36370 23380 36372
rect 23212 36318 23214 36370
rect 23266 36318 23380 36370
rect 23212 36316 23380 36318
rect 23548 36316 23828 36372
rect 23212 36306 23268 36316
rect 23100 35970 23156 35980
rect 23324 35810 23380 36316
rect 23660 35924 23716 35934
rect 23660 35830 23716 35868
rect 23324 35758 23326 35810
rect 23378 35758 23380 35810
rect 23324 35746 23380 35758
rect 22652 34750 22654 34802
rect 22706 34750 22708 34802
rect 22652 34738 22708 34750
rect 22876 35698 22932 35710
rect 22876 35646 22878 35698
rect 22930 35646 22932 35698
rect 22876 34914 22932 35646
rect 23212 35700 23268 35710
rect 23212 35606 23268 35644
rect 22876 34862 22878 34914
rect 22930 34862 22932 34914
rect 22092 34524 22260 34580
rect 21980 33796 22036 33806
rect 21868 31666 21924 31678
rect 21868 31614 21870 31666
rect 21922 31614 21924 31666
rect 21868 30548 21924 31614
rect 21868 30482 21924 30492
rect 20748 30382 20750 30434
rect 20802 30382 20804 30434
rect 20748 30370 20804 30382
rect 21420 30380 21812 30436
rect 21420 30322 21476 30380
rect 21420 30270 21422 30322
rect 21474 30270 21476 30322
rect 21420 30258 21476 30270
rect 20636 30210 20692 30222
rect 20636 30158 20638 30210
rect 20690 30158 20692 30210
rect 20636 29876 20692 30158
rect 21308 30212 21364 30222
rect 21308 30118 21364 30156
rect 21532 30212 21588 30222
rect 21532 30210 21700 30212
rect 21532 30158 21534 30210
rect 21586 30158 21700 30210
rect 21532 30156 21700 30158
rect 21532 30146 21588 30156
rect 20636 29316 20692 29820
rect 20860 29988 20916 29998
rect 20860 29650 20916 29932
rect 21532 29988 21588 29998
rect 21644 29988 21700 30156
rect 21980 30210 22036 33740
rect 22092 33346 22148 33358
rect 22092 33294 22094 33346
rect 22146 33294 22148 33346
rect 22092 32564 22148 33294
rect 22092 32498 22148 32508
rect 22092 32004 22148 32014
rect 22204 32004 22260 34524
rect 22876 33684 22932 34862
rect 23548 34914 23604 34926
rect 23548 34862 23550 34914
rect 23602 34862 23604 34914
rect 23548 34804 23604 34862
rect 23548 34738 23604 34748
rect 22092 32002 22260 32004
rect 22092 31950 22094 32002
rect 22146 31950 22260 32002
rect 22092 31948 22260 31950
rect 22316 33628 22932 33684
rect 23100 34692 23156 34702
rect 23100 34018 23156 34636
rect 23548 34242 23604 34254
rect 23548 34190 23550 34242
rect 23602 34190 23604 34242
rect 23100 33966 23102 34018
rect 23154 33966 23156 34018
rect 22092 31938 22148 31948
rect 22316 31780 22372 33628
rect 22876 33460 22932 33470
rect 22876 33346 22932 33404
rect 22876 33294 22878 33346
rect 22930 33294 22932 33346
rect 22876 33282 22932 33294
rect 23100 33236 23156 33966
rect 23324 34132 23380 34142
rect 23548 34132 23604 34190
rect 23100 33234 23268 33236
rect 23100 33182 23102 33234
rect 23154 33182 23268 33234
rect 23100 33180 23268 33182
rect 23100 33170 23156 33180
rect 23212 32786 23268 33180
rect 23212 32734 23214 32786
rect 23266 32734 23268 32786
rect 23212 32722 23268 32734
rect 22428 32564 22484 32574
rect 22484 32508 22596 32564
rect 22428 32470 22484 32508
rect 22092 31724 22372 31780
rect 22092 31106 22148 31724
rect 22092 31054 22094 31106
rect 22146 31054 22148 31106
rect 22092 31042 22148 31054
rect 22204 31554 22260 31566
rect 22204 31502 22206 31554
rect 22258 31502 22260 31554
rect 21980 30158 21982 30210
rect 22034 30158 22036 30210
rect 21980 30146 22036 30158
rect 22092 30434 22148 30446
rect 22092 30382 22094 30434
rect 22146 30382 22148 30434
rect 21588 29932 21924 29988
rect 21532 29922 21588 29932
rect 20860 29598 20862 29650
rect 20914 29598 20916 29650
rect 20860 29586 20916 29598
rect 21308 29876 21364 29886
rect 21196 29538 21252 29550
rect 21196 29486 21198 29538
rect 21250 29486 21252 29538
rect 20748 29428 20804 29438
rect 20804 29372 20916 29428
rect 20748 29362 20804 29372
rect 20636 29250 20692 29260
rect 20860 28866 20916 29372
rect 21196 29092 21252 29486
rect 21196 29026 21252 29036
rect 21308 29426 21364 29820
rect 21308 29374 21310 29426
rect 21362 29374 21364 29426
rect 20860 28814 20862 28866
rect 20914 28814 20916 28866
rect 20860 28802 20916 28814
rect 20524 28588 20692 28644
rect 20524 28420 20580 28430
rect 20524 28326 20580 28364
rect 20524 28196 20580 28206
rect 20636 28196 20692 28588
rect 20748 28420 20804 28430
rect 21084 28420 21140 28430
rect 20748 28418 20916 28420
rect 20748 28366 20750 28418
rect 20802 28366 20916 28418
rect 20748 28364 20916 28366
rect 20748 28354 20804 28364
rect 20636 28140 20804 28196
rect 20524 28082 20580 28140
rect 20524 28030 20526 28082
rect 20578 28030 20580 28082
rect 20524 28018 20580 28030
rect 20636 27748 20692 27758
rect 20636 27654 20692 27692
rect 20412 27246 20414 27298
rect 20466 27246 20468 27298
rect 20412 27234 20468 27246
rect 20636 27524 20692 27534
rect 20188 27020 20356 27076
rect 20076 27010 20132 27020
rect 19964 26796 20244 26852
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19628 26460 20020 26516
rect 19404 26450 19460 26460
rect 19516 26404 19572 26414
rect 19516 26310 19572 26348
rect 19404 26290 19460 26302
rect 19404 26238 19406 26290
rect 19458 26238 19460 26290
rect 19404 25956 19460 26238
rect 19404 25890 19460 25900
rect 19740 26290 19796 26302
rect 19740 26238 19742 26290
rect 19794 26238 19796 26290
rect 19628 25844 19684 25854
rect 19516 25732 19572 25742
rect 19516 25508 19572 25676
rect 19292 22866 19348 22876
rect 19404 25284 19460 25294
rect 18956 22306 19012 22316
rect 19068 22820 19124 22830
rect 19068 22258 19124 22764
rect 19404 22820 19460 25228
rect 19516 24946 19572 25452
rect 19516 24894 19518 24946
rect 19570 24894 19572 24946
rect 19516 24882 19572 24894
rect 19628 24162 19684 25788
rect 19740 25508 19796 26238
rect 19964 25732 20020 26460
rect 20076 26068 20132 26078
rect 20188 26068 20244 26796
rect 20132 26012 20244 26068
rect 20300 26290 20356 27020
rect 20636 26908 20692 27468
rect 20524 26852 20692 26908
rect 20524 26516 20580 26852
rect 20300 26238 20302 26290
rect 20354 26238 20356 26290
rect 20076 25974 20132 26012
rect 19964 25676 20244 25732
rect 19740 25442 19796 25452
rect 19964 25506 20020 25518
rect 19964 25454 19966 25506
rect 20018 25454 20020 25506
rect 19964 25284 20020 25454
rect 19964 25218 20020 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20188 24948 20244 25676
rect 20300 25172 20356 26238
rect 20300 25106 20356 25116
rect 20412 26460 20580 26516
rect 19964 24892 20356 24948
rect 19964 24834 20020 24892
rect 19964 24782 19966 24834
rect 20018 24782 20020 24834
rect 19964 24770 20020 24782
rect 19628 24110 19630 24162
rect 19682 24110 19684 24162
rect 19628 24098 19684 24110
rect 20076 24724 20132 24734
rect 19740 23940 19796 23950
rect 19740 23846 19796 23884
rect 20076 23938 20132 24668
rect 20076 23886 20078 23938
rect 20130 23886 20132 23938
rect 20076 23874 20132 23886
rect 20188 24050 20244 24062
rect 20188 23998 20190 24050
rect 20242 23998 20244 24050
rect 20188 23716 20244 23998
rect 20188 23650 20244 23660
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20076 23380 20132 23390
rect 19964 23324 20076 23380
rect 19404 22754 19460 22764
rect 19516 23042 19572 23054
rect 19516 22990 19518 23042
rect 19570 22990 19572 23042
rect 19516 22596 19572 22990
rect 19516 22530 19572 22540
rect 19628 22484 19684 22494
rect 19684 22428 19796 22484
rect 19628 22418 19684 22428
rect 19740 22370 19796 22428
rect 19964 22482 20020 23324
rect 20076 23314 20132 23324
rect 20300 23044 20356 24892
rect 20412 23380 20468 26460
rect 20524 26292 20580 26302
rect 20524 26198 20580 26236
rect 20636 26290 20692 26302
rect 20636 26238 20638 26290
rect 20690 26238 20692 26290
rect 20636 25284 20692 26238
rect 20748 25620 20804 28140
rect 20860 27748 20916 28364
rect 20860 27682 20916 27692
rect 21084 27524 21140 28364
rect 21084 27458 21140 27468
rect 21196 27748 21252 27758
rect 21196 27076 21252 27692
rect 20748 25554 20804 25564
rect 20860 26852 20916 26862
rect 20860 26066 20916 26796
rect 21196 26740 21252 27020
rect 20860 26014 20862 26066
rect 20914 26014 20916 26066
rect 20860 25396 20916 26014
rect 21084 26684 21252 26740
rect 21084 26180 21140 26684
rect 21084 25508 21140 26124
rect 20860 25330 20916 25340
rect 20972 25452 21140 25508
rect 20636 25218 20692 25228
rect 20748 25172 20804 25182
rect 20412 23314 20468 23324
rect 20524 23940 20580 23950
rect 20300 22988 20468 23044
rect 20076 22820 20132 22830
rect 20132 22764 20244 22820
rect 20076 22754 20132 22764
rect 19964 22430 19966 22482
rect 20018 22430 20020 22482
rect 19964 22418 20020 22430
rect 19740 22318 19742 22370
rect 19794 22318 19796 22370
rect 19740 22306 19796 22318
rect 20076 22372 20132 22382
rect 20076 22278 20132 22316
rect 19068 22206 19070 22258
rect 19122 22206 19124 22258
rect 18732 21812 18788 21822
rect 18732 21718 18788 21756
rect 18620 21532 18788 21588
rect 18172 21420 18452 21476
rect 18284 20804 18340 20814
rect 18060 20748 18228 20804
rect 17724 20290 17780 20300
rect 17836 20690 17892 20702
rect 17836 20638 17838 20690
rect 17890 20638 17892 20690
rect 17724 20018 17780 20030
rect 17724 19966 17726 20018
rect 17778 19966 17780 20018
rect 17724 19460 17780 19966
rect 17836 19906 17892 20638
rect 18172 20188 18228 20748
rect 17836 19854 17838 19906
rect 17890 19854 17892 19906
rect 17836 19842 17892 19854
rect 17948 20130 18004 20142
rect 17948 20078 17950 20130
rect 18002 20078 18004 20130
rect 17724 19394 17780 19404
rect 17612 18722 17668 18732
rect 17948 18564 18004 20078
rect 18060 20132 18228 20188
rect 18060 19572 18116 20132
rect 18172 20018 18228 20030
rect 18172 19966 18174 20018
rect 18226 19966 18228 20018
rect 18172 19908 18228 19966
rect 18172 19842 18228 19852
rect 18172 19572 18228 19582
rect 18060 19516 18172 19572
rect 18172 19506 18228 19516
rect 18284 19236 18340 20748
rect 18396 20356 18452 21420
rect 18396 20290 18452 20300
rect 18508 20916 18564 20926
rect 18508 20356 18564 20860
rect 18620 20802 18676 20814
rect 18620 20750 18622 20802
rect 18674 20750 18676 20802
rect 18620 20580 18676 20750
rect 18620 20514 18676 20524
rect 18732 20468 18788 21532
rect 18956 21586 19012 21598
rect 18956 21534 18958 21586
rect 19010 21534 19012 21586
rect 18956 21252 19012 21534
rect 18956 21186 19012 21196
rect 19068 20916 19124 22206
rect 19404 22148 19460 22158
rect 19404 22146 19684 22148
rect 19404 22094 19406 22146
rect 19458 22094 19684 22146
rect 19404 22092 19684 22094
rect 19404 22082 19460 22092
rect 19068 20850 19124 20860
rect 19292 21924 19348 21934
rect 19292 21586 19348 21868
rect 19404 21700 19460 21710
rect 19404 21606 19460 21644
rect 19516 21698 19572 21710
rect 19516 21646 19518 21698
rect 19570 21646 19572 21698
rect 19292 21534 19294 21586
rect 19346 21534 19348 21586
rect 19292 20916 19348 21534
rect 19292 20850 19348 20860
rect 18956 20804 19012 20814
rect 19516 20804 19572 21646
rect 19628 21140 19684 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20188 21700 20244 22764
rect 20412 22708 20468 22988
rect 20412 22370 20468 22652
rect 20412 22318 20414 22370
rect 20466 22318 20468 22370
rect 20412 22306 20468 22318
rect 20524 22148 20580 23884
rect 20188 21634 20244 21644
rect 20300 22092 20580 22148
rect 20636 23828 20692 23838
rect 19740 21588 19796 21598
rect 19740 21494 19796 21532
rect 20076 21588 20132 21598
rect 20076 21494 20132 21532
rect 19628 21074 19684 21084
rect 18956 20710 19012 20748
rect 19404 20748 19684 20804
rect 19068 20692 19124 20702
rect 19068 20598 19124 20636
rect 19292 20692 19348 20702
rect 18732 20412 18900 20468
rect 18508 20300 18788 20356
rect 18396 20018 18452 20030
rect 18396 19966 18398 20018
rect 18450 19966 18452 20018
rect 18396 19460 18452 19966
rect 18396 19394 18452 19404
rect 17948 18498 18004 18508
rect 18060 19180 18340 19236
rect 18508 19236 18564 20300
rect 18620 20130 18676 20142
rect 18620 20078 18622 20130
rect 18674 20078 18676 20130
rect 18620 19684 18676 20078
rect 18732 20130 18788 20300
rect 18732 20078 18734 20130
rect 18786 20078 18788 20130
rect 18732 20066 18788 20078
rect 18620 19618 18676 19628
rect 18844 19572 18900 20412
rect 19292 20186 19348 20636
rect 19404 20468 19460 20748
rect 19404 20402 19460 20412
rect 19516 20578 19572 20590
rect 19516 20526 19518 20578
rect 19570 20526 19572 20578
rect 19180 20132 19236 20170
rect 19292 20134 19294 20186
rect 19346 20134 19348 20186
rect 19292 20122 19348 20134
rect 19404 20130 19460 20142
rect 19180 20066 19236 20076
rect 19404 20078 19406 20130
rect 19458 20078 19460 20130
rect 19068 20018 19124 20030
rect 19068 19966 19070 20018
rect 19122 19966 19124 20018
rect 19068 19908 19124 19966
rect 19292 20020 19348 20030
rect 19404 20020 19460 20078
rect 19348 19964 19460 20020
rect 19292 19954 19348 19964
rect 19068 19842 19124 19852
rect 19292 19684 19348 19694
rect 19516 19684 19572 20526
rect 19628 19796 19684 20748
rect 20188 20802 20244 20814
rect 20188 20750 20190 20802
rect 20242 20750 20244 20802
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20188 20244 20244 20750
rect 20188 20178 20244 20188
rect 20300 20242 20356 22092
rect 20524 21700 20580 21710
rect 20524 21606 20580 21644
rect 20300 20190 20302 20242
rect 20354 20190 20356 20242
rect 20300 20178 20356 20190
rect 20412 21028 20468 21038
rect 19852 20018 19908 20030
rect 20188 20020 20244 20030
rect 19852 19966 19854 20018
rect 19906 19966 19908 20018
rect 19628 19740 19796 19796
rect 19516 19628 19684 19684
rect 18844 19516 19124 19572
rect 18844 19348 18900 19358
rect 18732 19346 18900 19348
rect 18732 19294 18846 19346
rect 18898 19294 18900 19346
rect 18732 19292 18900 19294
rect 18060 18676 18116 19180
rect 18508 19170 18564 19180
rect 18620 19234 18676 19246
rect 18620 19182 18622 19234
rect 18674 19182 18676 19234
rect 17612 18450 17668 18462
rect 17612 18398 17614 18450
rect 17666 18398 17668 18450
rect 17612 18340 17668 18398
rect 18060 18450 18116 18620
rect 18060 18398 18062 18450
rect 18114 18398 18116 18450
rect 18060 18386 18116 18398
rect 18172 19010 18228 19022
rect 18172 18958 18174 19010
rect 18226 18958 18228 19010
rect 17612 18274 17668 18284
rect 18060 18228 18116 18238
rect 18060 18134 18116 18172
rect 18172 17668 18228 18958
rect 18284 19010 18340 19022
rect 18284 18958 18286 19010
rect 18338 18958 18340 19010
rect 18284 18900 18340 18958
rect 18284 18834 18340 18844
rect 18396 19010 18452 19022
rect 18396 18958 18398 19010
rect 18450 18958 18452 19010
rect 18396 18564 18452 18958
rect 18508 19012 18564 19022
rect 18508 18674 18564 18956
rect 18508 18622 18510 18674
rect 18562 18622 18564 18674
rect 18508 18610 18564 18622
rect 17500 17042 17556 17052
rect 17948 17554 18004 17566
rect 17948 17502 17950 17554
rect 18002 17502 18004 17554
rect 17948 17108 18004 17502
rect 17612 16882 17668 16894
rect 17612 16830 17614 16882
rect 17666 16830 17668 16882
rect 17500 16772 17556 16782
rect 17500 16678 17556 16716
rect 17500 16436 17556 16446
rect 16940 14478 16942 14530
rect 16994 14478 16996 14530
rect 16940 13972 16996 14478
rect 16940 13906 16996 13916
rect 17052 15092 17220 15148
rect 17388 16380 17500 16436
rect 16716 13346 16772 13356
rect 16828 13746 16884 13758
rect 16828 13694 16830 13746
rect 16882 13694 16884 13746
rect 16716 13076 16772 13086
rect 16380 13010 16436 13020
rect 16492 13074 16772 13076
rect 16492 13022 16718 13074
rect 16770 13022 16772 13074
rect 16492 13020 16772 13022
rect 16268 12404 16324 12414
rect 16268 12310 16324 12348
rect 16492 12402 16548 13020
rect 16716 13010 16772 13020
rect 16828 12628 16884 13694
rect 16828 12562 16884 12572
rect 16940 13188 16996 13198
rect 16492 12350 16494 12402
rect 16546 12350 16548 12402
rect 16380 12292 16436 12302
rect 16380 12198 16436 12236
rect 16492 11732 16548 12350
rect 16716 12516 16772 12526
rect 16716 12404 16772 12460
rect 16940 12404 16996 13132
rect 17052 12962 17108 15092
rect 17276 14306 17332 14318
rect 17276 14254 17278 14306
rect 17330 14254 17332 14306
rect 17276 13860 17332 14254
rect 17276 13794 17332 13804
rect 17052 12910 17054 12962
rect 17106 12910 17108 12962
rect 17052 12898 17108 12910
rect 17388 12962 17444 16380
rect 17500 16370 17556 16380
rect 17612 15988 17668 16830
rect 17612 15894 17668 15932
rect 17500 15540 17556 15550
rect 17500 15446 17556 15484
rect 17948 15426 18004 17052
rect 18060 16884 18116 16894
rect 18060 16790 18116 16828
rect 17948 15374 17950 15426
rect 18002 15374 18004 15426
rect 17948 15362 18004 15374
rect 18172 15148 18228 17612
rect 18284 18508 18452 18564
rect 18284 17108 18340 18508
rect 18284 17042 18340 17052
rect 18396 18340 18452 18350
rect 18396 16882 18452 18284
rect 18620 17332 18676 19182
rect 18732 18228 18788 19292
rect 18844 19282 18900 19292
rect 19068 19124 19124 19516
rect 19292 19346 19348 19628
rect 19292 19294 19294 19346
rect 19346 19294 19348 19346
rect 19292 19282 19348 19294
rect 18844 19068 19124 19124
rect 18844 18450 18900 19068
rect 19628 18676 19684 19628
rect 19740 19460 19796 19740
rect 19852 19572 19908 19966
rect 19852 19506 19908 19516
rect 20076 19964 20188 20020
rect 19740 19394 19796 19404
rect 19740 19236 19796 19246
rect 19740 19142 19796 19180
rect 20076 19012 20132 19964
rect 20188 19926 20244 19964
rect 20188 19236 20244 19246
rect 20412 19236 20468 20972
rect 20524 21028 20580 21038
rect 20636 21028 20692 23772
rect 20524 21026 20692 21028
rect 20524 20974 20526 21026
rect 20578 20974 20692 21026
rect 20524 20972 20692 20974
rect 20524 20962 20580 20972
rect 20748 20804 20804 25116
rect 20860 24722 20916 24734
rect 20860 24670 20862 24722
rect 20914 24670 20916 24722
rect 20860 23940 20916 24670
rect 20860 23874 20916 23884
rect 20972 23716 21028 25452
rect 20636 20748 20804 20804
rect 20860 23660 21028 23716
rect 21084 25284 21140 25294
rect 20636 20020 20692 20748
rect 20636 19954 20692 19964
rect 20748 20580 20804 20590
rect 20748 20132 20804 20524
rect 20748 20018 20804 20076
rect 20748 19966 20750 20018
rect 20802 19966 20804 20018
rect 20524 19348 20580 19358
rect 20524 19254 20580 19292
rect 20188 19234 20468 19236
rect 20188 19182 20190 19234
rect 20242 19182 20468 19234
rect 20188 19180 20468 19182
rect 20188 19170 20244 19180
rect 20076 18946 20132 18956
rect 20524 18900 20580 18910
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 18844 18398 18846 18450
rect 18898 18398 18900 18450
rect 18844 18386 18900 18398
rect 19516 18620 19684 18676
rect 19404 18340 19460 18350
rect 19404 18246 19460 18284
rect 19180 18228 19236 18238
rect 18732 18172 18900 18228
rect 18620 17276 18788 17332
rect 18620 17108 18676 17118
rect 18620 17014 18676 17052
rect 18396 16830 18398 16882
rect 18450 16830 18452 16882
rect 18284 15652 18340 15662
rect 18396 15652 18452 16830
rect 18340 15596 18452 15652
rect 18508 16770 18564 16782
rect 18508 16718 18510 16770
rect 18562 16718 18564 16770
rect 18284 15586 18340 15596
rect 17948 15092 18004 15102
rect 17948 14532 18004 15036
rect 17836 14530 18004 14532
rect 17836 14478 17950 14530
rect 18002 14478 18004 14530
rect 17836 14476 18004 14478
rect 17724 14420 17780 14430
rect 17724 13970 17780 14364
rect 17724 13918 17726 13970
rect 17778 13918 17780 13970
rect 17724 13906 17780 13918
rect 17388 12910 17390 12962
rect 17442 12910 17444 12962
rect 17388 12898 17444 12910
rect 17500 13860 17556 13870
rect 17500 13746 17556 13804
rect 17500 13694 17502 13746
rect 17554 13694 17556 13746
rect 17164 12852 17220 12862
rect 17164 12758 17220 12796
rect 17500 12740 17556 13694
rect 16716 12402 16996 12404
rect 16716 12350 16718 12402
rect 16770 12350 16996 12402
rect 16716 12348 16996 12350
rect 17388 12684 17556 12740
rect 17724 13748 17780 13758
rect 16716 12338 16772 12348
rect 17164 12068 17220 12078
rect 16492 11666 16548 11676
rect 16940 11844 16996 11854
rect 16492 11506 16548 11518
rect 16492 11454 16494 11506
rect 16546 11454 16548 11506
rect 16268 10836 16324 10846
rect 16268 10742 16324 10780
rect 16380 10612 16436 10622
rect 16380 10518 16436 10556
rect 16492 10612 16548 11454
rect 16828 11284 16884 11294
rect 16828 11190 16884 11228
rect 16492 10610 16660 10612
rect 16492 10558 16494 10610
rect 16546 10558 16660 10610
rect 16492 10556 16660 10558
rect 16492 10546 16548 10556
rect 16380 9940 16436 9950
rect 16380 9846 16436 9884
rect 16268 9828 16324 9838
rect 16268 8258 16324 9772
rect 16492 8930 16548 8942
rect 16492 8878 16494 8930
rect 16546 8878 16548 8930
rect 16492 8818 16548 8878
rect 16492 8766 16494 8818
rect 16546 8766 16548 8818
rect 16492 8754 16548 8766
rect 16268 8206 16270 8258
rect 16322 8206 16324 8258
rect 16268 8194 16324 8206
rect 16380 7700 16436 7710
rect 16156 7698 16436 7700
rect 16156 7646 16382 7698
rect 16434 7646 16436 7698
rect 16156 7644 16436 7646
rect 16380 7634 16436 7644
rect 15820 7588 15876 7598
rect 15820 7494 15876 7532
rect 16268 7364 16324 7374
rect 16156 7252 16212 7262
rect 15596 5906 15764 5908
rect 15596 5854 15598 5906
rect 15650 5854 15764 5906
rect 15596 5852 15764 5854
rect 16044 7250 16212 7252
rect 16044 7198 16158 7250
rect 16210 7198 16212 7250
rect 16044 7196 16212 7198
rect 16044 5906 16100 7196
rect 16156 7186 16212 7196
rect 16268 6690 16324 7308
rect 16604 6916 16660 10556
rect 16940 10610 16996 11788
rect 17164 11284 17220 12012
rect 17164 11190 17220 11228
rect 17276 10836 17332 10846
rect 17388 10836 17444 12684
rect 17612 12178 17668 12190
rect 17612 12126 17614 12178
rect 17666 12126 17668 12178
rect 17612 11956 17668 12126
rect 17724 12180 17780 13692
rect 17836 12962 17892 14476
rect 17948 14466 18004 14476
rect 18060 15092 18228 15148
rect 17948 13746 18004 13758
rect 17948 13694 17950 13746
rect 18002 13694 18004 13746
rect 17948 13524 18004 13694
rect 17948 13458 18004 13468
rect 18060 13300 18116 15092
rect 18508 14532 18564 16718
rect 18732 16772 18788 17276
rect 18844 17220 18900 18172
rect 19068 18226 19236 18228
rect 19068 18174 19182 18226
rect 19234 18174 19236 18226
rect 19068 18172 19236 18174
rect 19068 18004 19124 18172
rect 19180 18162 19236 18172
rect 19516 18004 19572 18620
rect 19068 17948 19572 18004
rect 19628 18450 19684 18462
rect 19628 18398 19630 18450
rect 19682 18398 19684 18450
rect 18844 17154 18900 17164
rect 19404 17666 19460 17948
rect 19628 17892 19684 18398
rect 19852 18450 19908 18462
rect 19852 18398 19854 18450
rect 19906 18398 19908 18450
rect 19740 18340 19796 18350
rect 19740 18246 19796 18284
rect 19404 17614 19406 17666
rect 19458 17614 19460 17666
rect 19068 17108 19124 17118
rect 19068 16882 19124 17052
rect 19068 16830 19070 16882
rect 19122 16830 19124 16882
rect 19068 16818 19124 16830
rect 18844 16772 18900 16782
rect 18732 16770 18900 16772
rect 18732 16718 18846 16770
rect 18898 16718 18900 16770
rect 18732 16716 18900 16718
rect 18732 16324 18788 16716
rect 18844 16706 18900 16716
rect 18732 16258 18788 16268
rect 19404 15988 19460 17614
rect 19516 17836 19684 17892
rect 19852 17892 19908 18398
rect 20300 18452 20356 18462
rect 20300 18358 20356 18396
rect 19516 17444 19572 17836
rect 19852 17826 19908 17836
rect 19628 17668 19684 17678
rect 19628 17574 19684 17612
rect 19964 17668 20020 17678
rect 19964 17666 20468 17668
rect 19964 17614 19966 17666
rect 20018 17614 20468 17666
rect 19964 17612 20468 17614
rect 19964 17602 20020 17612
rect 19852 17554 19908 17566
rect 19852 17502 19854 17554
rect 19906 17502 19908 17554
rect 19852 17444 19908 17502
rect 19516 17378 19572 17388
rect 19628 17388 19908 17444
rect 20076 17444 20132 17482
rect 20132 17388 20244 17444
rect 19628 17220 19684 17388
rect 20076 17378 20132 17388
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19628 17154 19684 17164
rect 20076 16996 20132 17006
rect 20076 16882 20132 16940
rect 20076 16830 20078 16882
rect 20130 16830 20132 16882
rect 20076 16818 20132 16830
rect 19628 15988 19684 15998
rect 19404 15986 19684 15988
rect 19404 15934 19630 15986
rect 19682 15934 19684 15986
rect 19404 15932 19684 15934
rect 19628 15922 19684 15932
rect 19740 15876 19796 15914
rect 19740 15810 19796 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19068 15540 19124 15550
rect 19068 15314 19124 15484
rect 19068 15262 19070 15314
rect 19122 15262 19124 15314
rect 19068 15250 19124 15262
rect 19404 15316 19460 15326
rect 19404 15222 19460 15260
rect 18508 14466 18564 14476
rect 19628 14868 19684 14878
rect 18620 14420 18676 14430
rect 18620 14326 18676 14364
rect 19628 14196 19684 14812
rect 20188 14308 20244 17388
rect 20300 14308 20356 14318
rect 20188 14252 20300 14308
rect 20300 14242 20356 14252
rect 19628 14130 19684 14140
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20412 14084 20468 17612
rect 20524 17666 20580 18844
rect 20636 17892 20692 17902
rect 20636 17798 20692 17836
rect 20524 17614 20526 17666
rect 20578 17614 20580 17666
rect 20524 17602 20580 17614
rect 20636 17444 20692 17454
rect 20636 17350 20692 17388
rect 20636 16996 20692 17006
rect 20524 15988 20580 15998
rect 20524 15426 20580 15932
rect 20524 15374 20526 15426
rect 20578 15374 20580 15426
rect 20524 15362 20580 15374
rect 20412 14018 20468 14028
rect 19740 13972 19796 13982
rect 18060 13234 18116 13244
rect 18172 13746 18228 13758
rect 18172 13694 18174 13746
rect 18226 13694 18228 13746
rect 17836 12910 17838 12962
rect 17890 12910 17892 12962
rect 17836 12898 17892 12910
rect 18060 12964 18116 12974
rect 17836 12404 17892 12414
rect 18060 12404 18116 12908
rect 18172 12628 18228 13694
rect 19404 13634 19460 13646
rect 19404 13582 19406 13634
rect 19458 13582 19460 13634
rect 19180 13188 19236 13198
rect 18508 13076 18564 13086
rect 18732 13076 18788 13086
rect 18564 13020 18676 13076
rect 18508 13010 18564 13020
rect 18620 12962 18676 13020
rect 18620 12910 18622 12962
rect 18674 12910 18676 12962
rect 18620 12898 18676 12910
rect 18172 12562 18228 12572
rect 18620 12740 18676 12750
rect 18508 12404 18564 12442
rect 17836 12402 18004 12404
rect 17836 12350 17838 12402
rect 17890 12350 18004 12402
rect 17836 12348 18004 12350
rect 18060 12348 18228 12404
rect 17836 12338 17892 12348
rect 17836 12180 17892 12190
rect 17724 12178 17892 12180
rect 17724 12126 17838 12178
rect 17890 12126 17892 12178
rect 17724 12124 17892 12126
rect 17612 11890 17668 11900
rect 17836 11620 17892 12124
rect 17332 10780 17444 10836
rect 17500 11564 17892 11620
rect 17276 10770 17332 10780
rect 16940 10558 16942 10610
rect 16994 10558 16996 10610
rect 16940 10546 16996 10558
rect 17500 9716 17556 11564
rect 17948 11508 18004 12348
rect 18172 12290 18228 12348
rect 18508 12338 18564 12348
rect 18620 12402 18676 12684
rect 18620 12350 18622 12402
rect 18674 12350 18676 12402
rect 18620 12338 18676 12350
rect 18732 12402 18788 13020
rect 18732 12350 18734 12402
rect 18786 12350 18788 12402
rect 18732 12338 18788 12350
rect 18172 12238 18174 12290
rect 18226 12238 18228 12290
rect 18172 12226 18228 12238
rect 18620 12180 18676 12190
rect 18508 11956 18564 11966
rect 17948 11442 18004 11452
rect 18060 11844 18116 11854
rect 17612 11394 17668 11406
rect 17612 11342 17614 11394
rect 17666 11342 17668 11394
rect 17612 9828 17668 11342
rect 17724 10836 17780 10846
rect 18060 10836 18116 11788
rect 18396 11844 18452 11854
rect 18396 11620 18452 11788
rect 18396 11554 18452 11564
rect 18284 11508 18340 11518
rect 18284 11396 18340 11452
rect 18396 11396 18452 11406
rect 18284 11394 18452 11396
rect 18284 11342 18398 11394
rect 18450 11342 18452 11394
rect 18284 11340 18452 11342
rect 18396 11330 18452 11340
rect 18172 10836 18228 10846
rect 18060 10834 18228 10836
rect 18060 10782 18174 10834
rect 18226 10782 18228 10834
rect 18060 10780 18228 10782
rect 17724 10742 17780 10780
rect 18172 10770 18228 10780
rect 17836 10612 17892 10622
rect 17836 10518 17892 10556
rect 17948 10610 18004 10622
rect 17948 10558 17950 10610
rect 18002 10558 18004 10610
rect 17948 9940 18004 10558
rect 18508 10610 18564 11900
rect 18620 10948 18676 12124
rect 19068 12180 19124 12190
rect 18956 11956 19012 11966
rect 18956 11788 19012 11900
rect 18620 10882 18676 10892
rect 18844 11732 19012 11788
rect 18508 10558 18510 10610
rect 18562 10558 18564 10610
rect 18508 10546 18564 10558
rect 18732 10498 18788 10510
rect 18732 10446 18734 10498
rect 18786 10446 18788 10498
rect 18508 9940 18564 9950
rect 17948 9938 18564 9940
rect 17948 9886 18510 9938
rect 18562 9886 18564 9938
rect 17948 9884 18564 9886
rect 17724 9828 17780 9838
rect 17612 9772 17724 9828
rect 17724 9762 17780 9772
rect 17500 9660 17668 9716
rect 16828 9268 16884 9278
rect 16884 9212 16996 9268
rect 16828 9202 16884 9212
rect 16940 9154 16996 9212
rect 17388 9156 17444 9166
rect 16940 9102 16942 9154
rect 16994 9102 16996 9154
rect 16940 9090 16996 9102
rect 17276 9154 17444 9156
rect 17276 9102 17390 9154
rect 17442 9102 17444 9154
rect 17276 9100 17444 9102
rect 16828 8148 16884 8158
rect 16828 8054 16884 8092
rect 17052 8148 17108 8158
rect 17052 8054 17108 8092
rect 16716 8034 16772 8046
rect 16716 7982 16718 8034
rect 16770 7982 16772 8034
rect 16716 7476 16772 7982
rect 16940 8036 16996 8046
rect 16940 7942 16996 7980
rect 16940 7700 16996 7710
rect 16940 7606 16996 7644
rect 16716 7250 16772 7420
rect 17276 7476 17332 9100
rect 17388 9090 17444 9100
rect 17500 8258 17556 8270
rect 17500 8206 17502 8258
rect 17554 8206 17556 8258
rect 17500 7588 17556 8206
rect 17276 7382 17332 7420
rect 17388 7532 17500 7588
rect 16716 7198 16718 7250
rect 16770 7198 16772 7250
rect 16716 7186 16772 7198
rect 16716 6916 16772 6926
rect 16604 6860 16716 6916
rect 16716 6850 16772 6860
rect 16268 6638 16270 6690
rect 16322 6638 16324 6690
rect 16268 6626 16324 6638
rect 16380 6692 16436 6702
rect 16380 6130 16436 6636
rect 17052 6690 17108 6702
rect 17052 6638 17054 6690
rect 17106 6638 17108 6690
rect 16380 6078 16382 6130
rect 16434 6078 16436 6130
rect 16380 6066 16436 6078
rect 16716 6580 16772 6590
rect 16716 6130 16772 6524
rect 16716 6078 16718 6130
rect 16770 6078 16772 6130
rect 16716 6066 16772 6078
rect 16828 6132 16884 6142
rect 16828 6038 16884 6076
rect 16044 5854 16046 5906
rect 16098 5854 16100 5906
rect 15484 5124 15540 5134
rect 15484 5030 15540 5068
rect 15596 4788 15652 5852
rect 16044 5842 16100 5854
rect 16604 5906 16660 5918
rect 16604 5854 16606 5906
rect 16658 5854 16660 5906
rect 15820 5794 15876 5806
rect 15820 5742 15822 5794
rect 15874 5742 15876 5794
rect 15820 5348 15876 5742
rect 15820 5292 16212 5348
rect 16156 5234 16212 5292
rect 16156 5182 16158 5234
rect 16210 5182 16212 5234
rect 16156 5170 16212 5182
rect 16604 5236 16660 5854
rect 16604 5170 16660 5180
rect 17052 5124 17108 6638
rect 17388 6244 17444 7532
rect 17500 7522 17556 7532
rect 17500 7364 17556 7374
rect 17500 7270 17556 7308
rect 17500 6692 17556 6702
rect 17500 6578 17556 6636
rect 17500 6526 17502 6578
rect 17554 6526 17556 6578
rect 17500 6514 17556 6526
rect 15596 4722 15652 4732
rect 16044 5012 16100 5022
rect 15372 4508 15876 4564
rect 15820 3666 15876 4508
rect 16044 4450 16100 4956
rect 16044 4398 16046 4450
rect 16098 4398 16100 4450
rect 16044 4386 16100 4398
rect 16492 4788 16548 4798
rect 15820 3614 15822 3666
rect 15874 3614 15876 3666
rect 15820 3602 15876 3614
rect 16492 3666 16548 4732
rect 16828 4340 16884 4350
rect 17052 4340 17108 5068
rect 17276 6188 17444 6244
rect 17612 6244 17668 9660
rect 17724 9604 17780 9614
rect 17724 9266 17780 9548
rect 17724 9214 17726 9266
rect 17778 9214 17780 9266
rect 17724 9202 17780 9214
rect 18172 9604 18228 9614
rect 18172 8258 18228 9548
rect 18284 9268 18340 9278
rect 18284 9174 18340 9212
rect 18508 8820 18564 9884
rect 18732 9940 18788 10446
rect 18844 10500 18900 11732
rect 18956 10724 19012 10734
rect 18956 10630 19012 10668
rect 18844 10444 19012 10500
rect 18732 9874 18788 9884
rect 18620 9828 18676 9838
rect 18620 9042 18676 9772
rect 18620 8990 18622 9042
rect 18674 8990 18676 9042
rect 18620 8978 18676 8990
rect 18508 8764 18788 8820
rect 18172 8206 18174 8258
rect 18226 8206 18228 8258
rect 18172 8194 18228 8206
rect 18620 8484 18676 8494
rect 18508 8146 18564 8158
rect 18508 8094 18510 8146
rect 18562 8094 18564 8146
rect 17836 8036 17892 8046
rect 18508 8036 18564 8094
rect 17892 7980 18004 8036
rect 17836 7942 17892 7980
rect 17724 7474 17780 7486
rect 17724 7422 17726 7474
rect 17778 7422 17780 7474
rect 17724 7028 17780 7422
rect 17724 6962 17780 6972
rect 17836 7474 17892 7486
rect 17836 7422 17838 7474
rect 17890 7422 17892 7474
rect 17836 6802 17892 7422
rect 17836 6750 17838 6802
rect 17890 6750 17892 6802
rect 17836 6738 17892 6750
rect 17948 6690 18004 7980
rect 18508 7970 18564 7980
rect 18620 8034 18676 8428
rect 18620 7982 18622 8034
rect 18674 7982 18676 8034
rect 18620 7812 18676 7982
rect 18620 7746 18676 7756
rect 18620 7588 18676 7598
rect 18172 7476 18228 7486
rect 17948 6638 17950 6690
rect 18002 6638 18004 6690
rect 17724 6468 17780 6478
rect 17724 6374 17780 6412
rect 17612 6188 17892 6244
rect 17276 4788 17332 6188
rect 17500 6132 17556 6142
rect 17500 6038 17556 6076
rect 17612 5908 17668 5918
rect 17612 5814 17668 5852
rect 17724 5906 17780 5918
rect 17724 5854 17726 5906
rect 17778 5854 17780 5906
rect 17724 5796 17780 5854
rect 17724 5730 17780 5740
rect 17276 4722 17332 4732
rect 17612 4340 17668 4350
rect 16828 4338 17668 4340
rect 16828 4286 16830 4338
rect 16882 4286 17614 4338
rect 17666 4286 17668 4338
rect 16828 4284 17668 4286
rect 16828 4274 16884 4284
rect 17612 3778 17668 4284
rect 17612 3726 17614 3778
rect 17666 3726 17668 3778
rect 17612 3714 17668 3726
rect 16492 3614 16494 3666
rect 16546 3614 16548 3666
rect 16492 3602 16548 3614
rect 17724 3668 17780 3678
rect 17724 3574 17780 3612
rect 10780 1362 10836 1372
rect 15036 1316 15092 3388
rect 15260 3378 15316 3388
rect 17388 3444 17444 3454
rect 17836 3444 17892 6188
rect 17948 6132 18004 6638
rect 17948 6066 18004 6076
rect 18060 6692 18116 6702
rect 18060 5906 18116 6636
rect 18172 6690 18228 7420
rect 18508 7364 18564 7374
rect 18508 7270 18564 7308
rect 18172 6638 18174 6690
rect 18226 6638 18228 6690
rect 18172 6626 18228 6638
rect 18284 7028 18340 7038
rect 18620 7028 18676 7532
rect 18732 7140 18788 8764
rect 18844 8148 18900 8158
rect 18844 8054 18900 8092
rect 18844 7700 18900 7710
rect 18844 7606 18900 7644
rect 18844 7140 18900 7150
rect 18732 7084 18844 7140
rect 18844 7074 18900 7084
rect 18620 6972 18788 7028
rect 18284 6020 18340 6972
rect 18620 6578 18676 6590
rect 18620 6526 18622 6578
rect 18674 6526 18676 6578
rect 18060 5854 18062 5906
rect 18114 5854 18116 5906
rect 18060 5842 18116 5854
rect 18172 5964 18340 6020
rect 18396 6466 18452 6478
rect 18396 6414 18398 6466
rect 18450 6414 18452 6466
rect 18172 5460 18228 5964
rect 18060 5404 18228 5460
rect 18284 5796 18340 5806
rect 18060 4228 18116 5404
rect 18060 4162 18116 4172
rect 18172 5236 18228 5246
rect 18172 3668 18228 5180
rect 18284 5234 18340 5740
rect 18284 5182 18286 5234
rect 18338 5182 18340 5234
rect 18284 5170 18340 5182
rect 18396 5012 18452 6414
rect 18620 6468 18676 6526
rect 18620 6402 18676 6412
rect 18620 6020 18676 6030
rect 18620 5906 18676 5964
rect 18620 5854 18622 5906
rect 18674 5854 18676 5906
rect 18620 5842 18676 5854
rect 18396 4946 18452 4956
rect 18508 5572 18564 5582
rect 18284 4228 18340 4238
rect 18284 4134 18340 4172
rect 18396 3668 18452 3678
rect 18172 3666 18452 3668
rect 18172 3614 18398 3666
rect 18450 3614 18452 3666
rect 18172 3612 18452 3614
rect 18396 3602 18452 3612
rect 17388 3442 17892 3444
rect 17388 3390 17390 3442
rect 17442 3390 17892 3442
rect 17388 3388 17892 3390
rect 17388 3378 17444 3388
rect 18508 2548 18564 5516
rect 18732 5346 18788 6972
rect 18844 6580 18900 6590
rect 18844 6486 18900 6524
rect 18956 6356 19012 10444
rect 19068 9938 19124 12124
rect 19180 12180 19236 13132
rect 19292 12180 19348 12190
rect 19180 12178 19348 12180
rect 19180 12126 19182 12178
rect 19234 12126 19294 12178
rect 19346 12126 19348 12178
rect 19180 12124 19348 12126
rect 19180 12114 19236 12124
rect 19292 12114 19348 12124
rect 19180 10612 19236 10622
rect 19180 10518 19236 10556
rect 19068 9886 19070 9938
rect 19122 9886 19124 9938
rect 19068 9874 19124 9886
rect 19404 9828 19460 13582
rect 19740 12740 19796 13916
rect 20636 13746 20692 16940
rect 20748 16772 20804 19966
rect 20860 19684 20916 23660
rect 21084 21700 21140 25228
rect 21196 24610 21252 24622
rect 21196 24558 21198 24610
rect 21250 24558 21252 24610
rect 21196 22596 21252 24558
rect 21308 23826 21364 29374
rect 21756 29316 21812 29326
rect 21756 29222 21812 29260
rect 21868 29314 21924 29932
rect 21868 29262 21870 29314
rect 21922 29262 21924 29314
rect 21868 29250 21924 29262
rect 21420 29204 21476 29214
rect 21420 28754 21476 29148
rect 21420 28702 21422 28754
rect 21474 28702 21476 28754
rect 21420 28690 21476 28702
rect 21644 28868 21700 28878
rect 21980 28868 22036 28878
rect 22092 28868 22148 30382
rect 21700 28866 22148 28868
rect 21700 28814 21982 28866
rect 22034 28814 22148 28866
rect 21700 28812 22148 28814
rect 21420 27972 21476 27982
rect 21420 27878 21476 27916
rect 21644 26908 21700 28812
rect 21980 28802 22036 28812
rect 21756 28644 21812 28654
rect 21756 28642 21924 28644
rect 21756 28590 21758 28642
rect 21810 28590 21924 28642
rect 21756 28588 21924 28590
rect 21756 28578 21812 28588
rect 21868 27076 21924 28588
rect 22204 28420 22260 31502
rect 22428 31554 22484 31566
rect 22428 31502 22430 31554
rect 22482 31502 22484 31554
rect 22316 31332 22372 31342
rect 22428 31332 22484 31502
rect 22540 31556 22596 32508
rect 22652 32562 22708 32574
rect 23324 32564 23380 34076
rect 23436 34076 23604 34132
rect 23660 34244 23716 34254
rect 23436 33684 23492 34076
rect 23660 34020 23716 34188
rect 23436 33618 23492 33628
rect 23548 33964 23716 34020
rect 23436 33460 23492 33470
rect 23436 32788 23492 33404
rect 23436 32674 23492 32732
rect 23436 32622 23438 32674
rect 23490 32622 23492 32674
rect 23436 32610 23492 32622
rect 22652 32510 22654 32562
rect 22706 32510 22708 32562
rect 22652 32452 22708 32510
rect 23212 32508 23380 32564
rect 23100 32452 23156 32462
rect 22652 32450 23156 32452
rect 22652 32398 23102 32450
rect 23154 32398 23156 32450
rect 22652 32396 23156 32398
rect 23100 32386 23156 32396
rect 22988 32004 23044 32014
rect 22652 31892 22708 31902
rect 22652 31556 22708 31836
rect 22764 31780 22820 31790
rect 22764 31778 22932 31780
rect 22764 31726 22766 31778
rect 22818 31726 22932 31778
rect 22764 31724 22932 31726
rect 22764 31714 22820 31724
rect 22652 31500 22820 31556
rect 22540 31490 22596 31500
rect 22428 31276 22708 31332
rect 22316 30434 22372 31276
rect 22428 31108 22484 31146
rect 22428 31042 22484 31052
rect 22316 30382 22318 30434
rect 22370 30382 22372 30434
rect 22316 30370 22372 30382
rect 22652 30324 22708 31276
rect 22764 31218 22820 31500
rect 22876 31332 22932 31724
rect 22876 31266 22932 31276
rect 22764 31166 22766 31218
rect 22818 31166 22820 31218
rect 22764 30772 22820 31166
rect 22988 31108 23044 31948
rect 23100 31892 23156 31902
rect 23100 31798 23156 31836
rect 23212 31332 23268 32508
rect 23324 32340 23380 32350
rect 23324 31778 23380 32284
rect 23324 31726 23326 31778
rect 23378 31726 23380 31778
rect 23324 31714 23380 31726
rect 22988 31042 23044 31052
rect 23100 31276 23268 31332
rect 22764 30716 23044 30772
rect 22316 30212 22372 30222
rect 22316 29426 22372 30156
rect 22652 30100 22708 30268
rect 22764 30100 22820 30110
rect 22652 30098 22820 30100
rect 22652 30046 22766 30098
rect 22818 30046 22820 30098
rect 22652 30044 22820 30046
rect 22316 29374 22318 29426
rect 22370 29374 22372 29426
rect 22316 28866 22372 29374
rect 22316 28814 22318 28866
rect 22370 28814 22372 28866
rect 22316 28802 22372 28814
rect 22428 29986 22484 29998
rect 22428 29934 22430 29986
rect 22482 29934 22484 29986
rect 22428 28644 22484 29934
rect 22764 28756 22820 30044
rect 22652 28644 22708 28654
rect 22428 28642 22708 28644
rect 22428 28590 22654 28642
rect 22706 28590 22708 28642
rect 22428 28588 22708 28590
rect 22204 28354 22260 28364
rect 22428 28420 22484 28430
rect 22428 27858 22484 28364
rect 22428 27806 22430 27858
rect 22482 27806 22484 27858
rect 22428 27748 22484 27806
rect 22428 27682 22484 27692
rect 22540 28196 22596 28206
rect 22204 27412 22260 27422
rect 22092 27076 22148 27086
rect 21868 27020 22092 27076
rect 22092 26982 22148 27020
rect 21532 26852 21588 26862
rect 21644 26852 21812 26908
rect 21532 26758 21588 26796
rect 21532 26290 21588 26302
rect 21532 26238 21534 26290
rect 21586 26238 21588 26290
rect 21420 26180 21476 26190
rect 21420 26086 21476 26124
rect 21532 25732 21588 26238
rect 21756 25844 21812 26852
rect 21532 25666 21588 25676
rect 21644 25788 21812 25844
rect 22092 26180 22148 26190
rect 21644 24388 21700 25788
rect 21868 25620 21924 25630
rect 21756 25506 21812 25518
rect 21756 25454 21758 25506
rect 21810 25454 21812 25506
rect 21756 25284 21812 25454
rect 21756 25218 21812 25228
rect 21644 24332 21812 24388
rect 21420 23940 21476 23950
rect 21420 23846 21476 23884
rect 21308 23774 21310 23826
rect 21362 23774 21364 23826
rect 21308 23762 21364 23774
rect 21644 23042 21700 23054
rect 21644 22990 21646 23042
rect 21698 22990 21700 23042
rect 21644 22596 21700 22990
rect 21196 22540 21700 22596
rect 21196 21700 21252 21710
rect 21084 21644 21196 21700
rect 20860 19618 20916 19628
rect 20860 18788 20916 18798
rect 20860 18562 20916 18732
rect 20860 18510 20862 18562
rect 20914 18510 20916 18562
rect 20860 18498 20916 18510
rect 21196 18562 21252 21644
rect 21308 20580 21364 22540
rect 21532 22370 21588 22382
rect 21532 22318 21534 22370
rect 21586 22318 21588 22370
rect 21420 21812 21476 21822
rect 21420 21586 21476 21756
rect 21420 21534 21422 21586
rect 21474 21534 21476 21586
rect 21420 21252 21476 21534
rect 21420 21186 21476 21196
rect 21532 21028 21588 22318
rect 21644 21700 21700 21710
rect 21756 21700 21812 24332
rect 21868 23938 21924 25564
rect 21868 23886 21870 23938
rect 21922 23886 21924 23938
rect 21868 23874 21924 23886
rect 22092 22260 22148 26124
rect 22204 24948 22260 27356
rect 22540 27074 22596 28140
rect 22540 27022 22542 27074
rect 22594 27022 22596 27074
rect 22540 27010 22596 27022
rect 22652 26908 22708 28588
rect 22764 27858 22820 28700
rect 22988 28530 23044 30716
rect 23100 29652 23156 31276
rect 23212 30882 23268 30894
rect 23212 30830 23214 30882
rect 23266 30830 23268 30882
rect 23212 30772 23268 30830
rect 23548 30772 23604 33964
rect 23772 33684 23828 36316
rect 23884 35476 23940 37772
rect 23996 36484 24052 36522
rect 23996 36418 24052 36428
rect 24444 35812 24500 39566
rect 24892 39508 24948 39518
rect 24892 39414 24948 39452
rect 25004 39394 25060 39406
rect 25004 39342 25006 39394
rect 25058 39342 25060 39394
rect 25004 39060 25060 39342
rect 25004 38994 25060 39004
rect 24556 38948 24612 38958
rect 24556 38946 24724 38948
rect 24556 38894 24558 38946
rect 24610 38894 24724 38946
rect 24556 38892 24724 38894
rect 24556 38882 24612 38892
rect 24668 38836 24724 38892
rect 24668 38770 24724 38780
rect 24668 38612 24724 38622
rect 24668 37938 24724 38556
rect 25228 38612 25284 38622
rect 25228 38518 25284 38556
rect 24668 37886 24670 37938
rect 24722 37886 24724 37938
rect 24668 37874 24724 37886
rect 25228 37828 25284 37838
rect 25340 37828 25396 40572
rect 25564 40628 25620 40638
rect 25564 40534 25620 40572
rect 26236 40626 26292 41244
rect 26684 41186 26740 41806
rect 27132 41524 27188 42478
rect 27916 42532 27972 42542
rect 28252 42532 28308 43708
rect 27916 42530 28308 42532
rect 27916 42478 27918 42530
rect 27970 42478 28308 42530
rect 27916 42476 28308 42478
rect 27916 42466 27972 42476
rect 26684 41134 26686 41186
rect 26738 41134 26740 41186
rect 26684 41122 26740 41134
rect 26908 41468 27188 41524
rect 27916 41860 27972 41870
rect 26236 40574 26238 40626
rect 26290 40574 26292 40626
rect 25788 40516 25844 40526
rect 25788 40422 25844 40460
rect 25900 40514 25956 40526
rect 25900 40462 25902 40514
rect 25954 40462 25956 40514
rect 25900 40404 25956 40462
rect 26236 40404 26292 40574
rect 25900 40348 26292 40404
rect 26460 40402 26516 40414
rect 26460 40350 26462 40402
rect 26514 40350 26516 40402
rect 26012 39730 26068 39742
rect 26012 39678 26014 39730
rect 26066 39678 26068 39730
rect 26012 39396 26068 39678
rect 26124 39732 26180 39742
rect 26124 39618 26180 39676
rect 26124 39566 26126 39618
rect 26178 39566 26180 39618
rect 26124 39554 26180 39566
rect 26460 39396 26516 40350
rect 26908 40404 26964 41468
rect 27132 41300 27188 41310
rect 27020 41298 27860 41300
rect 27020 41246 27134 41298
rect 27186 41246 27860 41298
rect 27020 41244 27860 41246
rect 27020 40626 27076 41244
rect 27132 41234 27188 41244
rect 27468 41076 27524 41086
rect 27244 41074 27524 41076
rect 27244 41022 27470 41074
rect 27522 41022 27524 41074
rect 27244 41020 27524 41022
rect 27020 40574 27022 40626
rect 27074 40574 27076 40626
rect 27020 40562 27076 40574
rect 27132 40628 27188 40638
rect 27244 40628 27300 41020
rect 27468 41010 27524 41020
rect 27692 41074 27748 41086
rect 27692 41022 27694 41074
rect 27746 41022 27748 41074
rect 27132 40626 27300 40628
rect 27132 40574 27134 40626
rect 27186 40574 27300 40626
rect 27132 40572 27300 40574
rect 27468 40628 27524 40638
rect 27132 40562 27188 40572
rect 27468 40534 27524 40572
rect 27244 40404 27300 40414
rect 27692 40404 27748 41022
rect 27804 41076 27860 41244
rect 27916 41298 27972 41804
rect 27916 41246 27918 41298
rect 27970 41246 27972 41298
rect 27916 41234 27972 41246
rect 28028 41076 28084 41086
rect 27804 41074 28084 41076
rect 27804 41022 28030 41074
rect 28082 41022 28084 41074
rect 27804 41020 28084 41022
rect 28028 41010 28084 41020
rect 26908 40402 27748 40404
rect 26908 40350 27246 40402
rect 27298 40350 27748 40402
rect 26908 40348 27748 40350
rect 27804 40628 27860 40638
rect 26796 39508 26852 39518
rect 26796 39414 26852 39452
rect 26012 39340 26516 39396
rect 25452 38946 25508 38958
rect 25452 38894 25454 38946
rect 25506 38894 25508 38946
rect 25452 38612 25508 38894
rect 26012 38836 26068 38846
rect 25564 38834 26068 38836
rect 25564 38782 26014 38834
rect 26066 38782 26068 38834
rect 25564 38780 26068 38782
rect 25564 38722 25620 38780
rect 26012 38770 26068 38780
rect 25564 38670 25566 38722
rect 25618 38670 25620 38722
rect 25564 38658 25620 38670
rect 25452 38546 25508 38556
rect 26012 38612 26068 38622
rect 25676 38500 25732 38510
rect 25676 38162 25732 38444
rect 25676 38110 25678 38162
rect 25730 38110 25732 38162
rect 25676 38098 25732 38110
rect 26012 37938 26068 38556
rect 26012 37886 26014 37938
rect 26066 37886 26068 37938
rect 26012 37874 26068 37886
rect 25228 37826 25396 37828
rect 25228 37774 25230 37826
rect 25282 37774 25396 37826
rect 25228 37772 25396 37774
rect 25228 36932 25284 37772
rect 26124 37492 26180 39340
rect 26236 38834 26292 38846
rect 26236 38782 26238 38834
rect 26290 38782 26292 38834
rect 26236 38668 26292 38782
rect 27020 38722 27076 40348
rect 27244 40338 27300 40348
rect 27356 39732 27412 39742
rect 27356 39638 27412 39676
rect 27804 39732 27860 40572
rect 27916 40404 27972 40414
rect 27916 40310 27972 40348
rect 28252 39844 28308 39854
rect 28252 39750 28308 39788
rect 27804 39730 27972 39732
rect 27804 39678 27806 39730
rect 27858 39678 27972 39730
rect 27804 39676 27972 39678
rect 27804 39666 27860 39676
rect 27692 38946 27748 38958
rect 27692 38894 27694 38946
rect 27746 38894 27748 38946
rect 27244 38836 27300 38846
rect 27468 38836 27524 38846
rect 27244 38834 27524 38836
rect 27244 38782 27246 38834
rect 27298 38782 27470 38834
rect 27522 38782 27524 38834
rect 27244 38780 27524 38782
rect 27244 38770 27300 38780
rect 27468 38770 27524 38780
rect 27020 38670 27022 38722
rect 27074 38670 27076 38722
rect 26236 38612 26404 38668
rect 27020 38658 27076 38670
rect 27692 38668 27748 38894
rect 27804 38836 27860 38846
rect 27804 38742 27860 38780
rect 26348 37940 26404 38612
rect 27132 38612 27748 38668
rect 26348 37874 26404 37884
rect 27020 38164 27076 38174
rect 25228 36866 25284 36876
rect 26012 37436 26180 37492
rect 25900 36708 25956 36718
rect 24220 35756 24500 35812
rect 24668 36258 24724 36270
rect 24668 36206 24670 36258
rect 24722 36206 24724 36258
rect 23996 35700 24052 35710
rect 23996 35606 24052 35644
rect 23884 35420 24052 35476
rect 23884 34580 23940 34590
rect 23884 34242 23940 34524
rect 23996 34468 24052 35420
rect 23996 34402 24052 34412
rect 24108 34916 24164 34926
rect 23884 34190 23886 34242
rect 23938 34190 23940 34242
rect 23884 34178 23940 34190
rect 24108 34356 24164 34860
rect 24108 34130 24164 34300
rect 24108 34078 24110 34130
rect 24162 34078 24164 34130
rect 24108 34066 24164 34078
rect 23212 30716 23604 30772
rect 23660 33628 23828 33684
rect 23212 30210 23268 30222
rect 23212 30158 23214 30210
rect 23266 30158 23268 30210
rect 23212 29988 23268 30158
rect 23436 29988 23492 30716
rect 23548 30212 23604 30222
rect 23548 30118 23604 30156
rect 23436 29932 23604 29988
rect 23212 29922 23268 29932
rect 23436 29764 23492 29774
rect 23324 29652 23380 29662
rect 23100 29650 23380 29652
rect 23100 29598 23326 29650
rect 23378 29598 23380 29650
rect 23100 29596 23380 29598
rect 23324 29586 23380 29596
rect 23436 29650 23492 29708
rect 23436 29598 23438 29650
rect 23490 29598 23492 29650
rect 23436 29586 23492 29598
rect 23548 29652 23604 29932
rect 23660 29764 23716 33628
rect 24108 32788 24164 32798
rect 24108 32694 24164 32732
rect 23772 32562 23828 32574
rect 23772 32510 23774 32562
rect 23826 32510 23828 32562
rect 23772 30882 23828 32510
rect 23996 31890 24052 31902
rect 23996 31838 23998 31890
rect 24050 31838 24052 31890
rect 23996 31668 24052 31838
rect 24108 31780 24164 31790
rect 24108 31686 24164 31724
rect 23996 31220 24052 31612
rect 23996 31154 24052 31164
rect 23772 30830 23774 30882
rect 23826 30830 23828 30882
rect 23772 30548 23828 30830
rect 24108 30994 24164 31006
rect 24108 30942 24110 30994
rect 24162 30942 24164 30994
rect 23772 30482 23828 30492
rect 23996 30772 24052 30782
rect 23772 30324 23828 30334
rect 23772 29986 23828 30268
rect 23772 29934 23774 29986
rect 23826 29934 23828 29986
rect 23772 29922 23828 29934
rect 23996 29986 24052 30716
rect 24108 30660 24164 30942
rect 24108 30594 24164 30604
rect 24220 30436 24276 35756
rect 24444 35586 24500 35598
rect 24444 35534 24446 35586
rect 24498 35534 24500 35586
rect 24332 35028 24388 35038
rect 24332 34934 24388 34972
rect 24332 34244 24388 34254
rect 24444 34244 24500 35534
rect 24388 34188 24500 34244
rect 24668 35140 24724 36206
rect 25116 36258 25172 36270
rect 25116 36206 25118 36258
rect 25170 36206 25172 36258
rect 24332 34178 24388 34188
rect 24556 34132 24612 34142
rect 24556 34038 24612 34076
rect 24668 33684 24724 35084
rect 24668 33618 24724 33628
rect 25004 35700 25060 35710
rect 24892 33346 24948 33358
rect 24892 33294 24894 33346
rect 24946 33294 24948 33346
rect 24444 33236 24500 33246
rect 24332 33180 24444 33236
rect 24332 30770 24388 33180
rect 24444 33142 24500 33180
rect 24444 32900 24500 32910
rect 24444 32674 24500 32844
rect 24444 32622 24446 32674
rect 24498 32622 24500 32674
rect 24444 32610 24500 32622
rect 24556 32676 24612 32686
rect 24556 32674 24724 32676
rect 24556 32622 24558 32674
rect 24610 32622 24724 32674
rect 24556 32620 24724 32622
rect 24556 32610 24612 32620
rect 24556 32340 24612 32350
rect 24332 30718 24334 30770
rect 24386 30718 24388 30770
rect 24332 30706 24388 30718
rect 24444 32338 24612 32340
rect 24444 32286 24558 32338
rect 24610 32286 24612 32338
rect 24444 32284 24612 32286
rect 24444 30772 24500 32284
rect 24556 32274 24612 32284
rect 24444 30706 24500 30716
rect 24444 30436 24500 30446
rect 24220 30434 24500 30436
rect 24220 30382 24446 30434
rect 24498 30382 24500 30434
rect 24220 30380 24500 30382
rect 24444 30370 24500 30380
rect 24668 30324 24724 32620
rect 24892 32228 24948 33294
rect 24892 32162 24948 32172
rect 24780 31892 24836 31902
rect 24780 31666 24836 31836
rect 24780 31614 24782 31666
rect 24834 31614 24836 31666
rect 24780 31602 24836 31614
rect 24556 30268 24724 30324
rect 24780 30322 24836 30334
rect 24780 30270 24782 30322
rect 24834 30270 24836 30322
rect 24556 30100 24612 30268
rect 24780 30100 24836 30270
rect 24332 30098 24612 30100
rect 24332 30046 24558 30098
rect 24610 30046 24612 30098
rect 24332 30044 24612 30046
rect 23996 29934 23998 29986
rect 24050 29934 24052 29986
rect 23996 29922 24052 29934
rect 24220 29988 24276 29998
rect 24108 29764 24164 29774
rect 23660 29708 23940 29764
rect 23548 29596 23716 29652
rect 23212 29428 23268 29438
rect 22988 28478 22990 28530
rect 23042 28478 23044 28530
rect 22988 28466 23044 28478
rect 23100 29426 23268 29428
rect 23100 29374 23214 29426
rect 23266 29374 23268 29426
rect 23100 29372 23268 29374
rect 23100 29092 23156 29372
rect 23212 29362 23268 29372
rect 22764 27806 22766 27858
rect 22818 27806 22820 27858
rect 22764 27794 22820 27806
rect 23100 27076 23156 29036
rect 23436 29204 23492 29214
rect 23436 28642 23492 29148
rect 23436 28590 23438 28642
rect 23490 28590 23492 28642
rect 23436 28578 23492 28590
rect 23100 27010 23156 27020
rect 23212 27860 23268 27870
rect 23212 27074 23268 27804
rect 23548 27858 23604 27870
rect 23548 27806 23550 27858
rect 23602 27806 23604 27858
rect 23212 27022 23214 27074
rect 23266 27022 23268 27074
rect 23212 27010 23268 27022
rect 23324 27746 23380 27758
rect 23324 27694 23326 27746
rect 23378 27694 23380 27746
rect 23324 27186 23380 27694
rect 23324 27134 23326 27186
rect 23378 27134 23380 27186
rect 23324 26908 23380 27134
rect 22540 26852 22708 26908
rect 22876 26852 22932 26862
rect 22316 26292 22372 26302
rect 22316 26198 22372 26236
rect 22204 24882 22260 24892
rect 22540 24276 22596 26852
rect 22764 26290 22820 26302
rect 22764 26238 22766 26290
rect 22818 26238 22820 26290
rect 22764 25844 22820 26238
rect 22876 26066 22932 26796
rect 22876 26014 22878 26066
rect 22930 26014 22932 26066
rect 22876 26002 22932 26014
rect 23212 26852 23380 26908
rect 23212 26290 23268 26852
rect 23212 26238 23214 26290
rect 23266 26238 23268 26290
rect 22764 25778 22820 25788
rect 23212 25730 23268 26238
rect 23212 25678 23214 25730
rect 23266 25678 23268 25730
rect 23212 25666 23268 25678
rect 23324 26404 23380 26414
rect 22764 25284 22820 25294
rect 22540 24210 22596 24220
rect 22652 25228 22764 25284
rect 22652 24722 22708 25228
rect 22764 25218 22820 25228
rect 22652 24670 22654 24722
rect 22706 24670 22708 24722
rect 22652 23940 22708 24670
rect 22092 22194 22148 22204
rect 22204 23938 22708 23940
rect 22204 23886 22654 23938
rect 22706 23886 22708 23938
rect 22204 23884 22708 23886
rect 22204 22036 22260 23884
rect 22652 23874 22708 23884
rect 22764 24724 22820 24734
rect 23100 24724 23156 24734
rect 22764 23378 22820 24668
rect 22764 23326 22766 23378
rect 22818 23326 22820 23378
rect 22764 23314 22820 23326
rect 22988 24722 23156 24724
rect 22988 24670 23102 24722
rect 23154 24670 23156 24722
rect 22988 24668 23156 24670
rect 22428 23266 22484 23278
rect 22428 23214 22430 23266
rect 22482 23214 22484 23266
rect 21868 21980 22260 22036
rect 22316 22258 22372 22270
rect 22316 22206 22318 22258
rect 22370 22206 22372 22258
rect 21868 21812 21924 21980
rect 21868 21746 21924 21756
rect 21980 21868 22260 21924
rect 21644 21698 21812 21700
rect 21644 21646 21646 21698
rect 21698 21646 21812 21698
rect 21644 21644 21812 21646
rect 21644 21634 21700 21644
rect 21868 21586 21924 21598
rect 21868 21534 21870 21586
rect 21922 21534 21924 21586
rect 21532 20972 21700 21028
rect 21532 20804 21588 20814
rect 21532 20710 21588 20748
rect 21308 20524 21588 20580
rect 21420 19908 21476 19918
rect 21308 19906 21476 19908
rect 21308 19854 21422 19906
rect 21474 19854 21476 19906
rect 21308 19852 21476 19854
rect 21308 19346 21364 19852
rect 21420 19842 21476 19852
rect 21532 19796 21588 20524
rect 21644 20132 21700 20972
rect 21756 20916 21812 20926
rect 21756 20822 21812 20860
rect 21644 20066 21700 20076
rect 21308 19294 21310 19346
rect 21362 19294 21364 19346
rect 21308 19282 21364 19294
rect 21420 19684 21476 19694
rect 21420 19234 21476 19628
rect 21420 19182 21422 19234
rect 21474 19182 21476 19234
rect 21420 19170 21476 19182
rect 21532 19012 21588 19740
rect 21868 19236 21924 21534
rect 21868 19170 21924 19180
rect 21756 19124 21812 19134
rect 21756 19030 21812 19068
rect 21196 18510 21198 18562
rect 21250 18510 21252 18562
rect 21196 18498 21252 18510
rect 21420 18956 21588 19012
rect 21644 19012 21700 19022
rect 21420 18450 21476 18956
rect 21420 18398 21422 18450
rect 21474 18398 21476 18450
rect 21420 18386 21476 18398
rect 21532 18340 21588 18350
rect 20972 16772 21028 16782
rect 20748 16770 21028 16772
rect 20748 16718 20974 16770
rect 21026 16718 21028 16770
rect 20748 16716 21028 16718
rect 20748 16098 20804 16110
rect 20748 16046 20750 16098
rect 20802 16046 20804 16098
rect 20748 15988 20804 16046
rect 20748 15540 20804 15932
rect 20748 15474 20804 15484
rect 20860 15316 20916 15326
rect 20748 14644 20804 14654
rect 20748 13972 20804 14588
rect 20748 13906 20804 13916
rect 20636 13694 20638 13746
rect 20690 13694 20692 13746
rect 19516 12684 19796 12740
rect 20412 12964 20468 12974
rect 19516 12180 19572 12684
rect 19836 12572 20100 12582
rect 19628 12516 19684 12526
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19628 12404 19684 12460
rect 19852 12404 19908 12414
rect 19628 12402 19908 12404
rect 19628 12350 19854 12402
rect 19906 12350 19908 12402
rect 19628 12348 19908 12350
rect 19852 12338 19908 12348
rect 19964 12404 20020 12414
rect 20300 12404 20356 12414
rect 20020 12402 20356 12404
rect 20020 12350 20302 12402
rect 20354 12350 20356 12402
rect 20020 12348 20356 12350
rect 19964 12310 20020 12348
rect 20300 12338 20356 12348
rect 20412 12402 20468 12908
rect 20412 12350 20414 12402
rect 20466 12350 20468 12402
rect 20412 12338 20468 12350
rect 19740 12180 19796 12190
rect 19516 12178 19796 12180
rect 19516 12126 19742 12178
rect 19794 12126 19796 12178
rect 19516 12124 19796 12126
rect 19740 12114 19796 12124
rect 20524 12178 20580 12190
rect 20524 12126 20526 12178
rect 20578 12126 20580 12178
rect 19628 11956 19684 11966
rect 19404 9762 19460 9772
rect 19516 10948 19572 10958
rect 19516 10610 19572 10892
rect 19628 10724 19684 11900
rect 20300 11620 20356 11630
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19852 10724 19908 10734
rect 19628 10722 19908 10724
rect 19628 10670 19854 10722
rect 19906 10670 19908 10722
rect 19628 10668 19908 10670
rect 19516 10558 19518 10610
rect 19570 10558 19572 10610
rect 19404 9604 19460 9614
rect 19516 9604 19572 10558
rect 19852 10052 19908 10668
rect 20300 10612 20356 11564
rect 20524 11506 20580 12126
rect 20524 11454 20526 11506
rect 20578 11454 20580 11506
rect 20524 10948 20580 11454
rect 20636 11508 20692 13694
rect 20860 13524 20916 15260
rect 20972 15092 21028 16716
rect 21420 16436 21476 16446
rect 21420 16322 21476 16380
rect 21420 16270 21422 16322
rect 21474 16270 21476 16322
rect 21420 16258 21476 16270
rect 21308 15988 21364 15998
rect 20972 15026 21028 15036
rect 21084 15986 21364 15988
rect 21084 15934 21310 15986
rect 21362 15934 21364 15986
rect 21084 15932 21364 15934
rect 20860 13458 20916 13468
rect 20748 13076 20804 13086
rect 20748 12982 20804 13020
rect 20636 11442 20692 11452
rect 20748 12628 20804 12638
rect 20748 10948 20804 12572
rect 20972 12180 21028 12190
rect 20972 12086 21028 12124
rect 20524 10892 20692 10948
rect 20412 10836 20468 10846
rect 20412 10742 20468 10780
rect 20300 10556 20468 10612
rect 19852 9986 19908 9996
rect 19852 9604 19908 9614
rect 19404 9602 19908 9604
rect 19404 9550 19406 9602
rect 19458 9550 19854 9602
rect 19906 9550 19908 9602
rect 19404 9548 19908 9550
rect 19404 9380 19460 9548
rect 19852 9538 19908 9548
rect 20188 9604 20244 9614
rect 20188 9602 20356 9604
rect 20188 9550 20190 9602
rect 20242 9550 20356 9602
rect 20188 9548 20356 9550
rect 20188 9538 20244 9548
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19292 8932 19348 8942
rect 19292 8838 19348 8876
rect 19180 8372 19236 8382
rect 19180 8278 19236 8316
rect 19068 8146 19124 8158
rect 19068 8094 19070 8146
rect 19122 8094 19124 8146
rect 19068 7588 19124 8094
rect 19292 7700 19348 7710
rect 19292 7606 19348 7644
rect 19068 7522 19124 7532
rect 19404 6468 19460 9324
rect 20300 9268 20356 9548
rect 19516 8932 19572 8942
rect 19516 8258 19572 8876
rect 19516 8206 19518 8258
rect 19570 8206 19572 8258
rect 19516 7476 19572 8206
rect 19852 8372 19908 8382
rect 19852 8258 19908 8316
rect 19852 8206 19854 8258
rect 19906 8206 19908 8258
rect 19852 8194 19908 8206
rect 20188 8258 20244 8270
rect 20188 8206 20190 8258
rect 20242 8206 20244 8258
rect 19628 8034 19684 8046
rect 19628 7982 19630 8034
rect 19682 7982 19684 8034
rect 19628 7700 19684 7982
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19852 7700 19908 7710
rect 19628 7698 19908 7700
rect 19628 7646 19854 7698
rect 19906 7646 19908 7698
rect 19628 7644 19908 7646
rect 19628 7476 19684 7486
rect 19516 7474 19684 7476
rect 19516 7422 19630 7474
rect 19682 7422 19684 7474
rect 19516 7420 19684 7422
rect 19628 7410 19684 7420
rect 19740 6804 19796 7644
rect 19852 7634 19908 7644
rect 19964 7252 20020 7262
rect 19964 7158 20020 7196
rect 19628 6748 19796 6804
rect 19852 7140 19908 7150
rect 19516 6692 19572 6702
rect 19516 6598 19572 6636
rect 19404 6412 19572 6468
rect 18732 5294 18734 5346
rect 18786 5294 18788 5346
rect 18732 5282 18788 5294
rect 18844 6300 19012 6356
rect 18844 5234 18900 6300
rect 19292 6132 19348 6142
rect 19292 6038 19348 6076
rect 19068 5908 19124 5918
rect 18956 5906 19124 5908
rect 18956 5854 19070 5906
rect 19122 5854 19124 5906
rect 18956 5852 19124 5854
rect 18956 5796 19012 5852
rect 19068 5842 19124 5852
rect 18956 5730 19012 5740
rect 19180 5794 19236 5806
rect 19180 5742 19182 5794
rect 19234 5742 19236 5794
rect 19180 5348 19236 5742
rect 19180 5282 19236 5292
rect 19292 5346 19348 5358
rect 19292 5294 19294 5346
rect 19346 5294 19348 5346
rect 18844 5182 18846 5234
rect 18898 5182 18900 5234
rect 18844 5170 18900 5182
rect 19292 5234 19348 5294
rect 19292 5182 19294 5234
rect 19346 5182 19348 5234
rect 19292 5170 19348 5182
rect 19292 4788 19348 4798
rect 18844 3778 18900 3790
rect 18844 3726 18846 3778
rect 18898 3726 18900 3778
rect 18844 3668 18900 3726
rect 18844 3574 18900 3612
rect 19292 3666 19348 4732
rect 19516 4564 19572 6412
rect 19628 5796 19684 6748
rect 19852 6690 19908 7084
rect 20188 6804 20244 8206
rect 20300 7812 20356 9212
rect 20412 8148 20468 10556
rect 20636 9156 20692 10892
rect 20748 10882 20804 10892
rect 20860 11844 20916 11854
rect 20748 10724 20804 10734
rect 20748 10630 20804 10668
rect 20748 9716 20804 9726
rect 20748 9622 20804 9660
rect 20636 9090 20692 9100
rect 20860 8708 20916 11788
rect 21084 11060 21140 15932
rect 21308 15922 21364 15932
rect 21420 15764 21476 15774
rect 21420 14754 21476 15708
rect 21420 14702 21422 14754
rect 21474 14702 21476 14754
rect 21420 14690 21476 14702
rect 21196 14532 21252 14542
rect 21196 14308 21252 14476
rect 21308 14532 21364 14542
rect 21532 14532 21588 18284
rect 21644 17666 21700 18956
rect 21868 19010 21924 19022
rect 21868 18958 21870 19010
rect 21922 18958 21924 19010
rect 21868 18564 21924 18958
rect 21868 18498 21924 18508
rect 21980 17892 22036 21868
rect 22092 21698 22148 21710
rect 22092 21646 22094 21698
rect 22146 21646 22148 21698
rect 22092 20692 22148 21646
rect 22204 21698 22260 21868
rect 22204 21646 22206 21698
rect 22258 21646 22260 21698
rect 22204 21634 22260 21646
rect 22204 21476 22260 21486
rect 22316 21476 22372 22206
rect 22204 21474 22372 21476
rect 22204 21422 22206 21474
rect 22258 21422 22372 21474
rect 22204 21420 22372 21422
rect 22204 21410 22260 21420
rect 22204 21252 22260 21262
rect 22204 20802 22260 21196
rect 22204 20750 22206 20802
rect 22258 20750 22260 20802
rect 22204 20738 22260 20750
rect 22316 21140 22372 21150
rect 22092 20626 22148 20636
rect 22204 19908 22260 19918
rect 21980 17826 22036 17836
rect 22092 19236 22148 19246
rect 22092 18564 22148 19180
rect 22092 17668 22148 18508
rect 21644 17614 21646 17666
rect 21698 17614 21700 17666
rect 21644 15764 21700 17614
rect 21868 17612 22148 17668
rect 21868 17554 21924 17612
rect 21868 17502 21870 17554
rect 21922 17502 21924 17554
rect 21868 17490 21924 17502
rect 22204 17554 22260 19852
rect 22204 17502 22206 17554
rect 22258 17502 22260 17554
rect 22204 17490 22260 17502
rect 22316 17668 22372 21084
rect 22428 19460 22484 23214
rect 22876 23268 22932 23278
rect 22876 23174 22932 23212
rect 22652 23156 22708 23166
rect 22652 23154 22820 23156
rect 22652 23102 22654 23154
rect 22706 23102 22820 23154
rect 22652 23100 22820 23102
rect 22652 23090 22708 23100
rect 22764 21924 22820 23100
rect 22764 21858 22820 21868
rect 22988 22596 23044 24668
rect 23100 24658 23156 24668
rect 23324 24052 23380 26348
rect 23548 25844 23604 27806
rect 23660 26908 23716 29596
rect 23772 29426 23828 29438
rect 23772 29374 23774 29426
rect 23826 29374 23828 29426
rect 23772 27188 23828 29374
rect 23772 27122 23828 27132
rect 23660 26852 23828 26908
rect 23772 26180 23828 26852
rect 23772 26086 23828 26124
rect 23548 25778 23604 25788
rect 23436 25506 23492 25518
rect 23436 25454 23438 25506
rect 23490 25454 23492 25506
rect 23436 25284 23492 25454
rect 23436 25218 23492 25228
rect 23772 25284 23828 25294
rect 23660 24834 23716 24846
rect 23660 24782 23662 24834
rect 23714 24782 23716 24834
rect 23548 24724 23604 24734
rect 23548 24630 23604 24668
rect 23324 23996 23604 24052
rect 23100 23940 23156 23950
rect 23100 23846 23156 23884
rect 23436 23828 23492 23838
rect 23436 23734 23492 23772
rect 23324 23714 23380 23726
rect 23324 23662 23326 23714
rect 23378 23662 23380 23714
rect 23212 23380 23268 23390
rect 23212 23286 23268 23324
rect 22540 21588 22596 21598
rect 22540 19684 22596 21532
rect 22764 21476 22820 21486
rect 22764 20914 22820 21420
rect 22764 20862 22766 20914
rect 22818 20862 22820 20914
rect 22764 20850 22820 20862
rect 22540 19618 22596 19628
rect 22428 19404 22708 19460
rect 22428 19012 22484 19022
rect 22428 18918 22484 18956
rect 22540 18338 22596 18350
rect 22540 18286 22542 18338
rect 22594 18286 22596 18338
rect 22540 18116 22596 18286
rect 22540 18050 22596 18060
rect 22428 17668 22484 17678
rect 22316 17666 22484 17668
rect 22316 17614 22430 17666
rect 22482 17614 22484 17666
rect 22316 17612 22484 17614
rect 22316 16212 22372 17612
rect 22428 17602 22484 17612
rect 22428 17108 22484 17118
rect 22652 17108 22708 19404
rect 22764 19236 22820 19246
rect 22764 19122 22820 19180
rect 22764 19070 22766 19122
rect 22818 19070 22820 19122
rect 22764 18900 22820 19070
rect 22764 18834 22820 18844
rect 22876 18562 22932 18574
rect 22876 18510 22878 18562
rect 22930 18510 22932 18562
rect 22764 18450 22820 18462
rect 22764 18398 22766 18450
rect 22818 18398 22820 18450
rect 22764 18228 22820 18398
rect 22764 17668 22820 18172
rect 22764 17602 22820 17612
rect 22764 17108 22820 17118
rect 22652 17052 22764 17108
rect 22428 17014 22484 17052
rect 22764 17042 22820 17052
rect 22540 16884 22596 16894
rect 22540 16790 22596 16828
rect 22876 16772 22932 18510
rect 22988 16884 23044 22540
rect 23324 21588 23380 23662
rect 23548 23604 23604 23996
rect 23212 21532 23380 21588
rect 23436 23548 23604 23604
rect 23212 20804 23268 21532
rect 23324 21364 23380 21374
rect 23324 20914 23380 21308
rect 23324 20862 23326 20914
rect 23378 20862 23380 20914
rect 23324 20850 23380 20862
rect 23100 19684 23156 19694
rect 23100 19122 23156 19628
rect 23212 19460 23268 20748
rect 23436 20188 23492 23548
rect 23660 23380 23716 24782
rect 23660 23314 23716 23324
rect 23772 23938 23828 25228
rect 23884 24610 23940 29708
rect 24108 29650 24164 29708
rect 24108 29598 24110 29650
rect 24162 29598 24164 29650
rect 24108 29586 24164 29598
rect 24220 29650 24276 29932
rect 24220 29598 24222 29650
rect 24274 29598 24276 29650
rect 24220 29586 24276 29598
rect 24332 29650 24388 30044
rect 24332 29598 24334 29650
rect 24386 29598 24388 29650
rect 24332 29586 24388 29598
rect 24220 28868 24276 28878
rect 23996 28756 24052 28766
rect 23996 27300 24052 28700
rect 24108 28644 24164 28654
rect 24108 28550 24164 28588
rect 24108 27972 24164 27982
rect 24108 27878 24164 27916
rect 24220 27748 24276 28812
rect 24556 28082 24612 30044
rect 24668 30044 24836 30100
rect 24668 29092 24724 30044
rect 24668 29026 24724 29036
rect 24780 29426 24836 29438
rect 24780 29374 24782 29426
rect 24834 29374 24836 29426
rect 24556 28030 24558 28082
rect 24610 28030 24612 28082
rect 24444 27860 24500 27870
rect 24444 27766 24500 27804
rect 24220 27682 24276 27692
rect 24556 27636 24612 28030
rect 24780 28082 24836 29374
rect 24780 28030 24782 28082
rect 24834 28030 24836 28082
rect 24780 28018 24836 28030
rect 23996 26290 24052 27244
rect 24444 27580 24612 27636
rect 24332 26516 24388 26526
rect 24332 26422 24388 26460
rect 23996 26238 23998 26290
rect 24050 26238 24052 26290
rect 23996 26226 24052 26238
rect 24444 24948 24500 27580
rect 25004 26908 25060 35644
rect 25116 35588 25172 36206
rect 25900 35924 25956 36652
rect 25900 35858 25956 35868
rect 25340 35588 25396 35598
rect 25116 35586 25396 35588
rect 25116 35534 25342 35586
rect 25394 35534 25396 35586
rect 25116 35532 25396 35534
rect 25116 34804 25172 35532
rect 25340 35522 25396 35532
rect 25788 35588 25844 35598
rect 25788 35586 25956 35588
rect 25788 35534 25790 35586
rect 25842 35534 25956 35586
rect 25788 35532 25956 35534
rect 25788 35522 25844 35532
rect 25116 34738 25172 34748
rect 25228 34130 25284 34142
rect 25228 34078 25230 34130
rect 25282 34078 25284 34130
rect 25228 32674 25284 34078
rect 25340 34132 25396 34142
rect 25340 34038 25396 34076
rect 25452 34130 25508 34142
rect 25452 34078 25454 34130
rect 25506 34078 25508 34130
rect 25452 33236 25508 34078
rect 25788 34130 25844 34142
rect 25788 34078 25790 34130
rect 25842 34078 25844 34130
rect 25676 33348 25732 33358
rect 25452 33170 25508 33180
rect 25564 33346 25732 33348
rect 25564 33294 25678 33346
rect 25730 33294 25732 33346
rect 25564 33292 25732 33294
rect 25452 33012 25508 33022
rect 25228 32622 25230 32674
rect 25282 32622 25284 32674
rect 25228 32610 25284 32622
rect 25340 32956 25452 33012
rect 25228 31556 25284 31566
rect 25228 30434 25284 31500
rect 25340 31108 25396 32956
rect 25452 32946 25508 32956
rect 25452 32788 25508 32798
rect 25452 31778 25508 32732
rect 25564 32450 25620 33292
rect 25676 33282 25732 33292
rect 25564 32398 25566 32450
rect 25618 32398 25620 32450
rect 25564 31892 25620 32398
rect 25676 32562 25732 32574
rect 25676 32510 25678 32562
rect 25730 32510 25732 32562
rect 25676 32228 25732 32510
rect 25676 32162 25732 32172
rect 25564 31826 25620 31836
rect 25452 31726 25454 31778
rect 25506 31726 25508 31778
rect 25452 31714 25508 31726
rect 25788 31778 25844 34078
rect 25788 31726 25790 31778
rect 25842 31726 25844 31778
rect 25788 31714 25844 31726
rect 25564 31554 25620 31566
rect 25564 31502 25566 31554
rect 25618 31502 25620 31554
rect 25564 31444 25620 31502
rect 25620 31388 25732 31444
rect 25564 31378 25620 31388
rect 25676 31218 25732 31388
rect 25676 31166 25678 31218
rect 25730 31166 25732 31218
rect 25676 31154 25732 31166
rect 25340 31052 25508 31108
rect 25340 30884 25396 30922
rect 25340 30818 25396 30828
rect 25228 30382 25230 30434
rect 25282 30382 25284 30434
rect 25228 30370 25284 30382
rect 25340 30660 25396 30670
rect 25340 29652 25396 30604
rect 25228 29596 25396 29652
rect 25116 27188 25172 27198
rect 25116 27094 25172 27132
rect 24556 26852 25060 26908
rect 24556 25618 24612 26852
rect 24556 25566 24558 25618
rect 24610 25566 24612 25618
rect 24556 25554 24612 25566
rect 25004 25956 25060 25966
rect 23884 24558 23886 24610
rect 23938 24558 23940 24610
rect 23884 24546 23940 24558
rect 23996 24892 24500 24948
rect 24668 25506 24724 25518
rect 24668 25454 24670 25506
rect 24722 25454 24724 25506
rect 23772 23886 23774 23938
rect 23826 23886 23828 23938
rect 23772 23268 23828 23886
rect 23772 23202 23828 23212
rect 23772 23044 23828 23054
rect 23772 22950 23828 22988
rect 23548 22930 23604 22942
rect 23548 22878 23550 22930
rect 23602 22878 23604 22930
rect 23548 21588 23604 22878
rect 23772 22148 23828 22158
rect 23660 21700 23716 21710
rect 23660 21606 23716 21644
rect 23548 21522 23604 21532
rect 23772 20804 23828 22092
rect 23996 21698 24052 24892
rect 24444 24722 24500 24734
rect 24444 24670 24446 24722
rect 24498 24670 24500 24722
rect 24444 24050 24500 24670
rect 24444 23998 24446 24050
rect 24498 23998 24500 24050
rect 24444 23986 24500 23998
rect 24556 24050 24612 24062
rect 24556 23998 24558 24050
rect 24610 23998 24612 24050
rect 24220 23826 24276 23838
rect 24220 23774 24222 23826
rect 24274 23774 24276 23826
rect 24108 23380 24164 23390
rect 24108 23154 24164 23324
rect 24108 23102 24110 23154
rect 24162 23102 24164 23154
rect 24108 23090 24164 23102
rect 24220 21924 24276 23774
rect 24556 23380 24612 23998
rect 24556 23314 24612 23324
rect 24332 23268 24388 23278
rect 24332 23154 24388 23212
rect 24668 23266 24724 25454
rect 25004 25506 25060 25900
rect 25004 25454 25006 25506
rect 25058 25454 25060 25506
rect 25004 25442 25060 25454
rect 25228 25172 25284 29596
rect 25340 29314 25396 29326
rect 25340 29262 25342 29314
rect 25394 29262 25396 29314
rect 25340 28756 25396 29262
rect 25340 28690 25396 28700
rect 25340 28308 25396 28318
rect 25340 27860 25396 28252
rect 25340 27794 25396 27804
rect 25340 27076 25396 27086
rect 25340 26982 25396 27020
rect 25452 26908 25508 31052
rect 25900 30436 25956 35532
rect 26012 33012 26068 37436
rect 26124 37268 26180 37278
rect 26124 33684 26180 37212
rect 26348 37156 26404 37166
rect 26796 37156 26852 37166
rect 26348 37154 26852 37156
rect 26348 37102 26350 37154
rect 26402 37102 26798 37154
rect 26850 37102 26852 37154
rect 26348 37100 26852 37102
rect 26348 36932 26404 37100
rect 26348 36866 26404 36876
rect 26572 36484 26628 36494
rect 26236 36428 26572 36484
rect 26236 35812 26292 36428
rect 26572 36390 26628 36428
rect 26684 36260 26740 37100
rect 26796 37090 26852 37100
rect 26796 36708 26852 36718
rect 26796 36482 26852 36652
rect 27020 36596 27076 38108
rect 27132 37154 27188 38556
rect 27916 38164 27972 39676
rect 28140 39508 28196 39518
rect 28140 39414 28196 39452
rect 28364 39060 28420 43820
rect 29260 43764 29316 44942
rect 29932 44996 29988 45054
rect 29260 43698 29316 43708
rect 29596 44324 29652 44334
rect 29932 44324 29988 44940
rect 29596 44322 29988 44324
rect 29596 44270 29598 44322
rect 29650 44270 29988 44322
rect 29596 44268 29988 44270
rect 30492 44994 30548 45006
rect 30492 44942 30494 44994
rect 30546 44942 30548 44994
rect 30492 44324 30548 44942
rect 28476 43538 28532 43550
rect 28476 43486 28478 43538
rect 28530 43486 28532 43538
rect 28476 41300 28532 43486
rect 29036 43538 29092 43550
rect 29036 43486 29038 43538
rect 29090 43486 29092 43538
rect 28700 43204 28756 43214
rect 28588 41300 28644 41310
rect 28476 41298 28644 41300
rect 28476 41246 28590 41298
rect 28642 41246 28644 41298
rect 28476 41244 28644 41246
rect 28476 40628 28532 41244
rect 28588 41234 28644 41244
rect 28476 40562 28532 40572
rect 28588 40402 28644 40414
rect 28588 40350 28590 40402
rect 28642 40350 28644 40402
rect 28588 39396 28644 40350
rect 28588 39330 28644 39340
rect 28588 39060 28644 39070
rect 28364 39058 28644 39060
rect 28364 39006 28590 39058
rect 28642 39006 28644 39058
rect 28364 39004 28644 39006
rect 28364 38724 28420 39004
rect 28588 38994 28644 39004
rect 28364 38612 28532 38668
rect 27916 38098 27972 38108
rect 28476 38050 28532 38612
rect 28476 37998 28478 38050
rect 28530 37998 28532 38050
rect 28476 37986 28532 37998
rect 27132 37102 27134 37154
rect 27186 37102 27188 37154
rect 27132 37090 27188 37102
rect 27580 37940 27636 37950
rect 27580 37156 27636 37884
rect 27804 37940 27860 37950
rect 28140 37940 28196 37950
rect 27804 37938 28196 37940
rect 27804 37886 27806 37938
rect 27858 37886 28142 37938
rect 28194 37886 28196 37938
rect 27804 37884 28196 37886
rect 27804 37874 27860 37884
rect 28140 37874 28196 37884
rect 28252 37826 28308 37838
rect 28252 37774 28254 37826
rect 28306 37774 28308 37826
rect 28252 37380 28308 37774
rect 28252 37314 28308 37324
rect 28476 37716 28532 37726
rect 27580 37100 28196 37156
rect 27580 36708 27636 36718
rect 27580 36614 27636 36652
rect 27020 36540 27188 36596
rect 26796 36430 26798 36482
rect 26850 36430 26852 36482
rect 26796 36418 26852 36430
rect 27020 36372 27076 36382
rect 26796 36260 26852 36270
rect 26684 36204 26796 36260
rect 26796 36194 26852 36204
rect 26460 35924 26516 35934
rect 26236 35810 26404 35812
rect 26236 35758 26238 35810
rect 26290 35758 26404 35810
rect 26236 35756 26404 35758
rect 26236 35746 26292 35756
rect 26348 35028 26404 35756
rect 26460 35698 26516 35868
rect 26460 35646 26462 35698
rect 26514 35646 26516 35698
rect 26460 35634 26516 35646
rect 27020 35698 27076 36316
rect 27020 35646 27022 35698
rect 27074 35646 27076 35698
rect 27020 35634 27076 35646
rect 26796 35588 26852 35598
rect 26796 35494 26852 35532
rect 26460 35028 26516 35038
rect 26348 35026 26516 35028
rect 26348 34974 26462 35026
rect 26514 34974 26516 35026
rect 26348 34972 26516 34974
rect 26460 34962 26516 34972
rect 26572 34130 26628 34142
rect 26572 34078 26574 34130
rect 26626 34078 26628 34130
rect 26572 34020 26628 34078
rect 26572 33954 26628 33964
rect 26796 34018 26852 34030
rect 26796 33966 26798 34018
rect 26850 33966 26852 34018
rect 26236 33684 26292 33694
rect 26124 33628 26236 33684
rect 26236 33618 26292 33628
rect 26348 33234 26404 33246
rect 26348 33182 26350 33234
rect 26402 33182 26404 33234
rect 26348 33124 26404 33182
rect 26348 33058 26404 33068
rect 26796 33122 26852 33966
rect 26796 33070 26798 33122
rect 26850 33070 26852 33122
rect 26012 32946 26068 32956
rect 26684 32788 26740 32798
rect 26796 32788 26852 33070
rect 26740 32732 26852 32788
rect 27132 32788 27188 36540
rect 27356 36484 27412 36494
rect 27356 36390 27412 36428
rect 27916 36260 27972 36270
rect 27916 36258 28084 36260
rect 27916 36206 27918 36258
rect 27970 36206 28084 36258
rect 27916 36204 28084 36206
rect 27916 36194 27972 36204
rect 27692 35812 27748 35822
rect 27692 35718 27748 35756
rect 27468 35698 27524 35710
rect 27468 35646 27470 35698
rect 27522 35646 27524 35698
rect 27244 35586 27300 35598
rect 27244 35534 27246 35586
rect 27298 35534 27300 35586
rect 27244 35028 27300 35534
rect 27468 35588 27524 35646
rect 28028 35698 28084 36204
rect 28140 35922 28196 37100
rect 28140 35870 28142 35922
rect 28194 35870 28196 35922
rect 28140 35858 28196 35870
rect 28028 35646 28030 35698
rect 28082 35646 28084 35698
rect 28028 35634 28084 35646
rect 27468 35522 27524 35532
rect 28476 35138 28532 37660
rect 28588 36260 28644 36270
rect 28588 36166 28644 36204
rect 28588 35700 28644 35710
rect 28588 35606 28644 35644
rect 28476 35086 28478 35138
rect 28530 35086 28532 35138
rect 28476 35074 28532 35086
rect 27244 34962 27300 34972
rect 27356 34914 27412 34926
rect 27356 34862 27358 34914
rect 27410 34862 27412 34914
rect 27356 34804 27412 34862
rect 27580 34916 27636 34926
rect 27580 34822 27636 34860
rect 28252 34914 28308 34926
rect 28252 34862 28254 34914
rect 28306 34862 28308 34914
rect 27356 33458 27412 34748
rect 27468 34132 27524 34142
rect 27916 34132 27972 34142
rect 27468 34130 27972 34132
rect 27468 34078 27470 34130
rect 27522 34078 27918 34130
rect 27970 34078 27972 34130
rect 27468 34076 27972 34078
rect 27468 34066 27524 34076
rect 27356 33406 27358 33458
rect 27410 33406 27412 33458
rect 27356 33394 27412 33406
rect 27468 33572 27524 33582
rect 27132 32732 27412 32788
rect 26684 32722 26740 32732
rect 27020 32674 27076 32686
rect 27020 32622 27022 32674
rect 27074 32622 27076 32674
rect 26684 32340 26740 32350
rect 26460 31780 26516 31790
rect 26460 31686 26516 31724
rect 26012 30994 26068 31006
rect 26012 30942 26014 30994
rect 26066 30942 26068 30994
rect 26012 30772 26068 30942
rect 26684 30882 26740 32284
rect 27020 32340 27076 32622
rect 27244 32564 27300 32574
rect 27020 32274 27076 32284
rect 27132 32562 27300 32564
rect 27132 32510 27246 32562
rect 27298 32510 27300 32562
rect 27132 32508 27300 32510
rect 26796 31780 26852 31790
rect 26796 30994 26852 31724
rect 27132 31780 27188 32508
rect 27244 32498 27300 32508
rect 27132 31686 27188 31724
rect 26796 30942 26798 30994
rect 26850 30942 26852 30994
rect 26796 30930 26852 30942
rect 26684 30830 26686 30882
rect 26738 30830 26740 30882
rect 26684 30818 26740 30830
rect 26012 30706 26068 30716
rect 25900 30370 25956 30380
rect 25564 30212 25620 30222
rect 25788 30212 25844 30222
rect 26012 30212 26068 30222
rect 25564 30210 25732 30212
rect 25564 30158 25566 30210
rect 25618 30158 25732 30210
rect 25564 30156 25732 30158
rect 25564 30146 25620 30156
rect 25676 29652 25732 30156
rect 25788 30210 26068 30212
rect 25788 30158 25790 30210
rect 25842 30158 26014 30210
rect 26066 30158 26068 30210
rect 25788 30156 26068 30158
rect 25788 30146 25844 30156
rect 26012 30146 26068 30156
rect 27132 30210 27188 30222
rect 27132 30158 27134 30210
rect 27186 30158 27188 30210
rect 26348 30100 26404 30110
rect 26348 30098 26516 30100
rect 26348 30046 26350 30098
rect 26402 30046 26516 30098
rect 26348 30044 26516 30046
rect 26348 30034 26404 30044
rect 26236 29988 26292 29998
rect 25900 29986 26292 29988
rect 25900 29934 26238 29986
rect 26290 29934 26292 29986
rect 25900 29932 26292 29934
rect 25788 29652 25844 29662
rect 25676 29650 25844 29652
rect 25676 29598 25790 29650
rect 25842 29598 25844 29650
rect 25676 29596 25844 29598
rect 25788 29586 25844 29596
rect 25676 29426 25732 29438
rect 25676 29374 25678 29426
rect 25730 29374 25732 29426
rect 25676 29316 25732 29374
rect 25564 27748 25620 27758
rect 25676 27748 25732 29260
rect 25900 29426 25956 29932
rect 26236 29922 26292 29932
rect 25900 29374 25902 29426
rect 25954 29374 25956 29426
rect 25900 27860 25956 29374
rect 26236 29426 26292 29438
rect 26236 29374 26238 29426
rect 26290 29374 26292 29426
rect 26236 28980 26292 29374
rect 26460 29316 26516 30044
rect 27132 29650 27188 30158
rect 27132 29598 27134 29650
rect 27186 29598 27188 29650
rect 27132 29428 27188 29598
rect 27132 29362 27188 29372
rect 26572 29316 26628 29326
rect 26460 29260 26572 29316
rect 26572 29222 26628 29260
rect 27356 29204 27412 32732
rect 27468 32228 27524 33516
rect 27692 33458 27748 34076
rect 27916 34066 27972 34076
rect 28140 34130 28196 34142
rect 28140 34078 28142 34130
rect 28194 34078 28196 34130
rect 27692 33406 27694 33458
rect 27746 33406 27748 33458
rect 27692 33394 27748 33406
rect 27916 33348 27972 33358
rect 28140 33348 28196 34078
rect 28252 33570 28308 34862
rect 28700 34020 28756 43148
rect 28812 41860 28868 41870
rect 28812 41766 28868 41804
rect 29036 41748 29092 43486
rect 29372 43426 29428 43438
rect 29372 43374 29374 43426
rect 29426 43374 29428 43426
rect 29260 42868 29316 42878
rect 29260 42774 29316 42812
rect 29036 41682 29092 41692
rect 29148 42532 29204 42542
rect 29148 41076 29204 42476
rect 29372 42196 29428 43374
rect 29484 42866 29540 42878
rect 29484 42814 29486 42866
rect 29538 42814 29540 42866
rect 29484 42756 29540 42814
rect 29484 42690 29540 42700
rect 29484 42532 29540 42542
rect 29484 42438 29540 42476
rect 29260 42140 29428 42196
rect 29260 41972 29316 42140
rect 29484 41972 29540 41982
rect 29596 41972 29652 44268
rect 30492 44258 30548 44268
rect 30268 44212 30324 44222
rect 30268 44118 30324 44156
rect 30828 43988 30884 43998
rect 31164 43988 31220 45838
rect 31388 44996 31444 45006
rect 31388 44902 31444 44940
rect 31836 44548 31892 49200
rect 33404 46116 33460 49200
rect 33404 46050 33460 46060
rect 32172 45890 32228 45902
rect 32172 45838 32174 45890
rect 32226 45838 32228 45890
rect 31836 44482 31892 44492
rect 31948 44994 32004 45006
rect 31948 44942 31950 44994
rect 32002 44942 32004 44994
rect 30884 43932 31220 43988
rect 29708 43540 29764 43550
rect 29708 43446 29764 43484
rect 30156 43538 30212 43550
rect 30156 43486 30158 43538
rect 30210 43486 30212 43538
rect 30044 42868 30100 42878
rect 30044 42308 30100 42812
rect 30044 42242 30100 42252
rect 30044 41972 30100 41982
rect 29260 41412 29316 41916
rect 29260 41346 29316 41356
rect 29372 41970 30100 41972
rect 29372 41918 29486 41970
rect 29538 41918 30046 41970
rect 30098 41918 30100 41970
rect 29372 41916 30100 41918
rect 29148 40514 29204 41020
rect 29148 40462 29150 40514
rect 29202 40462 29204 40514
rect 29148 40450 29204 40462
rect 29036 40290 29092 40302
rect 29036 40238 29038 40290
rect 29090 40238 29092 40290
rect 29036 39844 29092 40238
rect 29036 39732 29092 39788
rect 29260 39732 29316 39742
rect 29036 39730 29316 39732
rect 29036 39678 29262 39730
rect 29314 39678 29316 39730
rect 29036 39676 29316 39678
rect 29260 39666 29316 39676
rect 29372 39732 29428 41916
rect 29484 41906 29540 41916
rect 30044 41906 30100 41916
rect 29932 41748 29988 41758
rect 30156 41748 30212 43486
rect 30828 43428 30884 43932
rect 31052 43764 31108 43774
rect 30940 43652 30996 43662
rect 30940 43558 30996 43596
rect 30828 43372 30996 43428
rect 30940 43204 30996 43372
rect 31052 43426 31108 43708
rect 31164 43540 31220 43550
rect 31612 43540 31668 43550
rect 31220 43538 31668 43540
rect 31220 43486 31614 43538
rect 31666 43486 31668 43538
rect 31220 43484 31668 43486
rect 31164 43446 31220 43484
rect 31612 43474 31668 43484
rect 31052 43374 31054 43426
rect 31106 43374 31108 43426
rect 31052 43362 31108 43374
rect 30940 43148 31108 43204
rect 30828 43092 30884 43102
rect 30268 42754 30324 42766
rect 30268 42702 30270 42754
rect 30322 42702 30324 42754
rect 30268 42532 30324 42702
rect 30268 42466 30324 42476
rect 30716 42084 30772 42094
rect 30716 41970 30772 42028
rect 30716 41918 30718 41970
rect 30770 41918 30772 41970
rect 30716 41906 30772 41918
rect 30604 41858 30660 41870
rect 30604 41806 30606 41858
rect 30658 41806 30660 41858
rect 30604 41748 30660 41806
rect 30156 41692 30548 41748
rect 29932 41298 29988 41692
rect 30156 41412 30212 41422
rect 30156 41318 30212 41356
rect 30492 41410 30548 41692
rect 30492 41358 30494 41410
rect 30546 41358 30548 41410
rect 30492 41346 30548 41358
rect 29932 41246 29934 41298
rect 29986 41246 29988 41298
rect 29932 41234 29988 41246
rect 29596 40962 29652 40974
rect 29596 40910 29598 40962
rect 29650 40910 29652 40962
rect 29596 40740 29652 40910
rect 29596 40674 29652 40684
rect 30156 40514 30212 40526
rect 30156 40462 30158 40514
rect 30210 40462 30212 40514
rect 30156 39956 30212 40462
rect 30268 40402 30324 40414
rect 30268 40350 30270 40402
rect 30322 40350 30324 40402
rect 30268 40292 30324 40350
rect 30268 40226 30324 40236
rect 30156 39890 30212 39900
rect 29372 39666 29428 39676
rect 29484 39618 29540 39630
rect 29484 39566 29486 39618
rect 29538 39566 29540 39618
rect 29036 39508 29092 39518
rect 29036 39058 29092 39452
rect 29484 39396 29540 39566
rect 30156 39620 30212 39630
rect 30156 39526 30212 39564
rect 29484 39330 29540 39340
rect 30604 39394 30660 41692
rect 30604 39342 30606 39394
rect 30658 39342 30660 39394
rect 30604 39330 30660 39342
rect 29036 39006 29038 39058
rect 29090 39006 29092 39058
rect 29036 38994 29092 39006
rect 29148 38948 29204 38958
rect 29148 38854 29204 38892
rect 30044 38948 30100 38958
rect 29708 38834 29764 38846
rect 29708 38782 29710 38834
rect 29762 38782 29764 38834
rect 28924 38722 28980 38734
rect 28924 38670 28926 38722
rect 28978 38670 28980 38722
rect 28924 38668 28980 38670
rect 29708 38668 29764 38782
rect 30044 38834 30100 38892
rect 30044 38782 30046 38834
rect 30098 38782 30100 38834
rect 30044 38770 30100 38782
rect 28924 38612 29764 38668
rect 28924 36596 28980 38612
rect 29596 38162 29652 38174
rect 29596 38110 29598 38162
rect 29650 38110 29652 38162
rect 29260 37938 29316 37950
rect 29260 37886 29262 37938
rect 29314 37886 29316 37938
rect 29260 37716 29316 37886
rect 29260 37650 29316 37660
rect 29484 37826 29540 37838
rect 29484 37774 29486 37826
rect 29538 37774 29540 37826
rect 29484 37604 29540 37774
rect 29596 37828 29652 38110
rect 29596 37762 29652 37772
rect 29708 38164 29764 38174
rect 29484 37538 29540 37548
rect 29260 37380 29316 37390
rect 29260 37286 29316 37324
rect 28924 36530 28980 36540
rect 29148 36372 29204 36382
rect 29148 36278 29204 36316
rect 29260 36258 29316 36270
rect 29260 36206 29262 36258
rect 29314 36206 29316 36258
rect 29148 35810 29204 35822
rect 29148 35758 29150 35810
rect 29202 35758 29204 35810
rect 29148 35700 29204 35758
rect 29260 35812 29316 36206
rect 29260 35746 29316 35756
rect 29372 36258 29428 36270
rect 29372 36206 29374 36258
rect 29426 36206 29428 36258
rect 29148 35634 29204 35644
rect 29372 35700 29428 36206
rect 29372 35634 29428 35644
rect 29596 36260 29652 36270
rect 29708 36260 29764 38108
rect 30044 38050 30100 38062
rect 30044 37998 30046 38050
rect 30098 37998 30100 38050
rect 30044 37604 30100 37998
rect 30268 38050 30324 38062
rect 30268 37998 30270 38050
rect 30322 37998 30324 38050
rect 30268 37716 30324 37998
rect 30828 38052 30884 43036
rect 30940 42980 30996 42990
rect 30940 42866 30996 42924
rect 30940 42814 30942 42866
rect 30994 42814 30996 42866
rect 30940 42802 30996 42814
rect 30828 37986 30884 37996
rect 30940 37938 30996 37950
rect 30940 37886 30942 37938
rect 30994 37886 30996 37938
rect 30268 37650 30324 37660
rect 30828 37828 30884 37838
rect 30044 37538 30100 37548
rect 30044 37268 30100 37278
rect 30044 37174 30100 37212
rect 30828 37266 30884 37772
rect 30828 37214 30830 37266
rect 30882 37214 30884 37266
rect 30828 37202 30884 37214
rect 30940 36820 30996 37886
rect 31052 37492 31108 43148
rect 31276 42756 31332 42766
rect 31836 42756 31892 42766
rect 31276 42662 31332 42700
rect 31500 42754 31892 42756
rect 31500 42702 31838 42754
rect 31890 42702 31892 42754
rect 31500 42700 31892 42702
rect 31500 42084 31556 42700
rect 31836 42690 31892 42700
rect 31164 41860 31220 41870
rect 31164 41766 31220 41804
rect 31500 41410 31556 42028
rect 31500 41358 31502 41410
rect 31554 41358 31556 41410
rect 31500 41346 31556 41358
rect 31836 42308 31892 42318
rect 31836 41186 31892 42252
rect 31948 41970 32004 44942
rect 32172 44996 32228 45838
rect 32956 45778 33012 45790
rect 32956 45726 32958 45778
rect 33010 45726 33012 45778
rect 32508 45108 32564 45118
rect 32508 45106 32900 45108
rect 32508 45054 32510 45106
rect 32562 45054 32900 45106
rect 32508 45052 32900 45054
rect 32508 45042 32564 45052
rect 32172 44930 32228 44940
rect 32396 44434 32452 44446
rect 32396 44382 32398 44434
rect 32450 44382 32452 44434
rect 32396 44324 32452 44382
rect 32732 44324 32788 44334
rect 32396 44322 32788 44324
rect 32396 44270 32734 44322
rect 32786 44270 32788 44322
rect 32396 44268 32788 44270
rect 32732 44258 32788 44268
rect 32284 44212 32340 44222
rect 32060 43652 32116 43662
rect 32060 43538 32116 43596
rect 32060 43486 32062 43538
rect 32114 43486 32116 43538
rect 32060 43092 32116 43486
rect 32060 43026 32116 43036
rect 31948 41918 31950 41970
rect 32002 41918 32004 41970
rect 31948 41906 32004 41918
rect 32172 42756 32228 42766
rect 31836 41134 31838 41186
rect 31890 41134 31892 41186
rect 31836 41122 31892 41134
rect 32172 41186 32228 42700
rect 32172 41134 32174 41186
rect 32226 41134 32228 41186
rect 32172 41122 32228 41134
rect 31164 41074 31220 41086
rect 31164 41022 31166 41074
rect 31218 41022 31220 41074
rect 31164 40402 31220 41022
rect 31948 41076 32004 41086
rect 31948 40982 32004 41020
rect 31164 40350 31166 40402
rect 31218 40350 31220 40402
rect 31164 39620 31220 40350
rect 31388 40962 31444 40974
rect 31388 40910 31390 40962
rect 31442 40910 31444 40962
rect 31388 40292 31444 40910
rect 31948 40852 32004 40862
rect 31388 40226 31444 40236
rect 31836 40292 31892 40302
rect 31164 39526 31220 39564
rect 31836 39618 31892 40236
rect 31836 39566 31838 39618
rect 31890 39566 31892 39618
rect 31836 39554 31892 39566
rect 31948 39620 32004 40796
rect 31276 38948 31332 38958
rect 31276 38854 31332 38892
rect 31836 38724 31892 38734
rect 31388 38276 31444 38286
rect 31388 38274 31668 38276
rect 31388 38222 31390 38274
rect 31442 38222 31668 38274
rect 31388 38220 31668 38222
rect 31388 38210 31444 38220
rect 31500 37938 31556 37950
rect 31500 37886 31502 37938
rect 31554 37886 31556 37938
rect 31388 37826 31444 37838
rect 31388 37774 31390 37826
rect 31442 37774 31444 37826
rect 31388 37716 31444 37774
rect 31388 37650 31444 37660
rect 31500 37604 31556 37886
rect 31500 37538 31556 37548
rect 31052 37426 31108 37436
rect 30828 36764 30996 36820
rect 31052 37266 31108 37278
rect 31052 37214 31054 37266
rect 31106 37214 31108 37266
rect 30380 36484 30436 36494
rect 29596 36258 29764 36260
rect 29596 36206 29598 36258
rect 29650 36206 29764 36258
rect 29596 36204 29764 36206
rect 29820 36482 30436 36484
rect 29820 36430 30382 36482
rect 30434 36430 30436 36482
rect 29820 36428 30436 36430
rect 29596 35588 29652 36204
rect 29708 35588 29764 35598
rect 29596 35586 29764 35588
rect 29596 35534 29710 35586
rect 29762 35534 29764 35586
rect 29596 35532 29764 35534
rect 29148 34914 29204 34926
rect 29148 34862 29150 34914
rect 29202 34862 29204 34914
rect 29148 34468 29204 34862
rect 29148 34402 29204 34412
rect 29372 34914 29428 34926
rect 29372 34862 29374 34914
rect 29426 34862 29428 34914
rect 28812 34244 28868 34254
rect 29372 34244 29428 34862
rect 29596 34356 29652 35532
rect 29708 35522 29764 35532
rect 29708 35140 29764 35150
rect 29820 35140 29876 36428
rect 30380 36418 30436 36428
rect 30044 35924 30100 35934
rect 30044 35810 30100 35868
rect 30044 35758 30046 35810
rect 30098 35758 30100 35810
rect 30044 35746 30100 35758
rect 30156 35810 30212 35822
rect 30156 35758 30158 35810
rect 30210 35758 30212 35810
rect 29708 35138 29876 35140
rect 29708 35086 29710 35138
rect 29762 35086 29876 35138
rect 29708 35084 29876 35086
rect 29708 35074 29764 35084
rect 30156 35028 30212 35758
rect 30156 34962 30212 34972
rect 30380 35698 30436 35710
rect 30380 35646 30382 35698
rect 30434 35646 30436 35698
rect 30380 34914 30436 35646
rect 30492 35700 30548 35710
rect 30492 35138 30548 35644
rect 30828 35586 30884 36764
rect 31052 36596 31108 37214
rect 31612 37268 31668 38220
rect 31724 37268 31780 37278
rect 31612 37266 31780 37268
rect 31612 37214 31726 37266
rect 31778 37214 31780 37266
rect 31612 37212 31780 37214
rect 31724 37202 31780 37212
rect 31836 37154 31892 38668
rect 31948 38500 32004 39564
rect 32060 39732 32116 39742
rect 32060 39058 32116 39676
rect 32172 39508 32228 39518
rect 32172 39414 32228 39452
rect 32060 39006 32062 39058
rect 32114 39006 32116 39058
rect 32060 38668 32116 39006
rect 32284 39060 32340 44156
rect 32844 43764 32900 45052
rect 32508 43428 32564 43438
rect 32508 43334 32564 43372
rect 32396 41970 32452 41982
rect 32396 41918 32398 41970
rect 32450 41918 32452 41970
rect 32396 41188 32452 41918
rect 32508 41972 32564 41982
rect 32508 41878 32564 41916
rect 32844 41410 32900 43708
rect 32844 41358 32846 41410
rect 32898 41358 32900 41410
rect 32844 41346 32900 41358
rect 32396 41122 32452 41132
rect 32508 40962 32564 40974
rect 32508 40910 32510 40962
rect 32562 40910 32564 40962
rect 32508 40740 32564 40910
rect 32508 40674 32564 40684
rect 32508 40516 32564 40526
rect 32508 40422 32564 40460
rect 32956 40180 33012 45726
rect 33180 45106 33236 45118
rect 33180 45054 33182 45106
rect 33234 45054 33236 45106
rect 33180 44996 33236 45054
rect 33180 44930 33236 44940
rect 33964 44994 34020 45006
rect 33964 44942 33966 44994
rect 34018 44942 34020 44994
rect 33740 44548 33796 44558
rect 33740 44454 33796 44492
rect 33964 44100 34020 44942
rect 33964 44034 34020 44044
rect 34860 44212 34916 44222
rect 34076 43762 34132 43774
rect 34076 43710 34078 43762
rect 34130 43710 34132 43762
rect 33404 43650 33460 43662
rect 33404 43598 33406 43650
rect 33458 43598 33460 43650
rect 33292 43538 33348 43550
rect 33292 43486 33294 43538
rect 33346 43486 33348 43538
rect 33180 42868 33236 42878
rect 33068 41970 33124 41982
rect 33068 41918 33070 41970
rect 33122 41918 33124 41970
rect 33068 41748 33124 41918
rect 33068 41682 33124 41692
rect 33180 41410 33236 42812
rect 33180 41358 33182 41410
rect 33234 41358 33236 41410
rect 33180 41346 33236 41358
rect 33068 41188 33124 41198
rect 33068 41074 33124 41132
rect 33068 41022 33070 41074
rect 33122 41022 33124 41074
rect 33068 40514 33124 41022
rect 33068 40462 33070 40514
rect 33122 40462 33124 40514
rect 33068 40450 33124 40462
rect 33292 40740 33348 43486
rect 33404 41636 33460 43598
rect 33964 43538 34020 43550
rect 33964 43486 33966 43538
rect 34018 43486 34020 43538
rect 33964 42868 34020 43486
rect 34076 43316 34132 43710
rect 34748 43652 34804 43662
rect 34076 43250 34132 43260
rect 34636 43596 34748 43652
rect 33964 42802 34020 42812
rect 34076 43092 34132 43102
rect 34076 42866 34132 43036
rect 34076 42814 34078 42866
rect 34130 42814 34132 42866
rect 34076 42802 34132 42814
rect 33740 42756 33796 42766
rect 33516 42754 33796 42756
rect 33516 42702 33742 42754
rect 33794 42702 33796 42754
rect 33516 42700 33796 42702
rect 33516 41858 33572 42700
rect 33740 42690 33796 42700
rect 34188 42756 34244 42766
rect 34188 42662 34244 42700
rect 33628 42420 33684 42430
rect 33628 41972 33684 42364
rect 34636 42082 34692 43596
rect 34748 43558 34804 43596
rect 34860 43650 34916 44156
rect 34860 43598 34862 43650
rect 34914 43598 34916 43650
rect 34860 43586 34916 43598
rect 34972 43428 35028 49200
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35084 46002 35140 46014
rect 35084 45950 35086 46002
rect 35138 45950 35140 46002
rect 35084 45892 35140 45950
rect 35084 45826 35140 45836
rect 35980 45892 36036 45902
rect 35980 45798 36036 45836
rect 36428 45106 36484 45118
rect 36428 45054 36430 45106
rect 36482 45054 36484 45106
rect 36092 44996 36148 45006
rect 35868 44994 36148 44996
rect 35868 44942 36094 44994
rect 36146 44942 36148 44994
rect 35868 44940 36148 44942
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35868 43652 35924 44940
rect 36092 44930 36148 44940
rect 36428 44996 36484 45054
rect 36428 44930 36484 44940
rect 36540 44548 36596 49200
rect 36988 46116 37044 46126
rect 36988 46022 37044 46060
rect 38108 46116 38164 49200
rect 39676 46340 39732 49200
rect 38108 46050 38164 46060
rect 39564 46284 39732 46340
rect 38892 45892 38948 45902
rect 38780 45890 38948 45892
rect 38780 45838 38894 45890
rect 38946 45838 38948 45890
rect 38780 45836 38948 45838
rect 37212 44996 37268 45006
rect 37212 44994 37828 44996
rect 37212 44942 37214 44994
rect 37266 44942 37828 44994
rect 37212 44940 37828 44942
rect 37212 44930 37268 44940
rect 36540 44482 36596 44492
rect 37212 44548 37268 44558
rect 37212 44454 37268 44492
rect 36316 44434 36372 44446
rect 36316 44382 36318 44434
rect 36370 44382 36372 44434
rect 35980 44324 36036 44334
rect 35980 44322 36260 44324
rect 35980 44270 35982 44322
rect 36034 44270 36260 44322
rect 35980 44268 36260 44270
rect 35980 44258 36036 44268
rect 35868 43586 35924 43596
rect 35420 43428 35476 43438
rect 34972 43426 35476 43428
rect 34972 43374 35422 43426
rect 35474 43374 35476 43426
rect 34972 43372 35476 43374
rect 35420 43362 35476 43372
rect 34748 43314 34804 43326
rect 34748 43262 34750 43314
rect 34802 43262 34804 43314
rect 34748 42644 34804 43262
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35308 42980 35364 42990
rect 35308 42866 35364 42924
rect 35308 42814 35310 42866
rect 35362 42814 35364 42866
rect 35308 42802 35364 42814
rect 35868 42980 35924 42990
rect 34748 42578 34804 42588
rect 35532 42754 35588 42766
rect 35532 42702 35534 42754
rect 35586 42702 35588 42754
rect 34636 42030 34638 42082
rect 34690 42030 34692 42082
rect 34636 42018 34692 42030
rect 33628 41906 33684 41916
rect 33516 41806 33518 41858
rect 33570 41806 33572 41858
rect 33516 41794 33572 41806
rect 34412 41860 34468 41870
rect 34412 41766 34468 41804
rect 35532 41860 35588 42702
rect 35868 41970 35924 42924
rect 36204 42866 36260 44268
rect 36316 44212 36372 44382
rect 36316 44146 36372 44156
rect 37548 43540 37604 43550
rect 37548 43446 37604 43484
rect 37548 43092 37604 43102
rect 37100 42980 37156 42990
rect 37100 42886 37156 42924
rect 36204 42814 36206 42866
rect 36258 42814 36260 42866
rect 36204 42802 36260 42814
rect 37100 42644 37156 42654
rect 37100 42550 37156 42588
rect 37212 42642 37268 42654
rect 37212 42590 37214 42642
rect 37266 42590 37268 42642
rect 37212 42196 37268 42590
rect 37212 42130 37268 42140
rect 36428 42084 36484 42094
rect 36428 41990 36484 42028
rect 36988 42082 37044 42094
rect 36988 42030 36990 42082
rect 37042 42030 37044 42082
rect 36764 41972 36820 41982
rect 35868 41918 35870 41970
rect 35922 41918 35924 41970
rect 35868 41906 35924 41918
rect 36540 41970 36820 41972
rect 36540 41918 36766 41970
rect 36818 41918 36820 41970
rect 36540 41916 36820 41918
rect 35532 41794 35588 41804
rect 33404 41570 33460 41580
rect 33740 41636 33796 41646
rect 33292 40402 33348 40684
rect 33292 40350 33294 40402
rect 33346 40350 33348 40402
rect 33292 40338 33348 40350
rect 33628 41186 33684 41198
rect 33628 41134 33630 41186
rect 33682 41134 33684 41186
rect 32956 40114 33012 40124
rect 33404 39956 33460 39966
rect 33404 39730 33460 39900
rect 33404 39678 33406 39730
rect 33458 39678 33460 39730
rect 33404 39666 33460 39678
rect 33516 39732 33572 39742
rect 33628 39732 33684 41134
rect 33740 40402 33796 41580
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 36540 41524 36596 41916
rect 36764 41906 36820 41916
rect 35196 41514 35460 41524
rect 35868 41468 36596 41524
rect 36876 41858 36932 41870
rect 36876 41806 36878 41858
rect 36930 41806 36932 41858
rect 35196 41188 35252 41198
rect 34300 41076 34356 41086
rect 34300 40982 34356 41020
rect 35196 40516 35252 41132
rect 33740 40350 33742 40402
rect 33794 40350 33796 40402
rect 33740 40338 33796 40350
rect 35084 40404 35140 40414
rect 35084 40310 35140 40348
rect 35196 40290 35252 40460
rect 35532 40516 35588 40526
rect 35868 40516 35924 41468
rect 36428 41300 36484 41310
rect 36428 41298 36596 41300
rect 36428 41246 36430 41298
rect 36482 41246 36596 41298
rect 36428 41244 36596 41246
rect 36428 41234 36484 41244
rect 35980 41076 36036 41086
rect 35980 40626 36036 41020
rect 36428 41076 36484 41086
rect 36316 40964 36372 40974
rect 35980 40574 35982 40626
rect 36034 40574 36036 40626
rect 35980 40562 36036 40574
rect 36204 40740 36260 40750
rect 35532 40514 35924 40516
rect 35532 40462 35534 40514
rect 35586 40462 35870 40514
rect 35922 40462 35924 40514
rect 35532 40460 35924 40462
rect 35532 40450 35588 40460
rect 35868 40450 35924 40460
rect 36204 40514 36260 40684
rect 36204 40462 36206 40514
rect 36258 40462 36260 40514
rect 36204 40450 36260 40462
rect 35196 40238 35198 40290
rect 35250 40238 35252 40290
rect 35196 40226 35252 40238
rect 36316 40404 36372 40908
rect 36428 40514 36484 41020
rect 36428 40462 36430 40514
rect 36482 40462 36484 40514
rect 36428 40450 36484 40462
rect 33572 39676 33684 39732
rect 33964 40180 34020 40190
rect 33516 39666 33572 39676
rect 32284 38724 32340 39004
rect 32508 39618 32564 39630
rect 32508 39566 32510 39618
rect 32562 39566 32564 39618
rect 32508 38948 32564 39566
rect 33180 39618 33236 39630
rect 33180 39566 33182 39618
rect 33234 39566 33236 39618
rect 32508 38882 32564 38892
rect 32732 39506 32788 39518
rect 32732 39454 32734 39506
rect 32786 39454 32788 39506
rect 32508 38724 32564 38734
rect 32284 38722 32564 38724
rect 32284 38670 32510 38722
rect 32562 38670 32564 38722
rect 32284 38668 32564 38670
rect 32060 38612 32228 38668
rect 32508 38658 32564 38668
rect 32732 38724 32788 39454
rect 32732 38658 32788 38668
rect 33180 38724 33236 39566
rect 33740 39618 33796 39630
rect 33740 39566 33742 39618
rect 33794 39566 33796 39618
rect 33628 39506 33684 39518
rect 33628 39454 33630 39506
rect 33682 39454 33684 39506
rect 33404 38948 33460 38958
rect 33628 38948 33684 39454
rect 33740 39508 33796 39566
rect 33740 39442 33796 39452
rect 33460 38892 33684 38948
rect 33404 38834 33460 38892
rect 33404 38782 33406 38834
rect 33458 38782 33460 38834
rect 33404 38770 33460 38782
rect 33180 38658 33236 38668
rect 31948 38434 32004 38444
rect 31948 38052 32004 38062
rect 32172 38052 32228 38612
rect 33852 38612 33908 38622
rect 32396 38500 32452 38510
rect 31948 38050 32228 38052
rect 31948 37998 31950 38050
rect 32002 37998 32228 38050
rect 31948 37996 32228 37998
rect 32284 38052 32340 38062
rect 31948 37268 32004 37996
rect 31948 37202 32004 37212
rect 31836 37102 31838 37154
rect 31890 37102 31892 37154
rect 31836 37090 31892 37102
rect 31052 36594 31220 36596
rect 31052 36542 31054 36594
rect 31106 36542 31220 36594
rect 31052 36540 31220 36542
rect 31052 36530 31108 36540
rect 30828 35534 30830 35586
rect 30882 35534 30884 35586
rect 30828 35522 30884 35534
rect 30940 36482 30996 36494
rect 30940 36430 30942 36482
rect 30994 36430 30996 36482
rect 30940 35700 30996 36430
rect 30940 35364 30996 35644
rect 30492 35086 30494 35138
rect 30546 35086 30548 35138
rect 30492 35074 30548 35086
rect 30828 35308 30996 35364
rect 31052 36372 31108 36382
rect 30380 34862 30382 34914
rect 30434 34862 30436 34914
rect 30380 34850 30436 34862
rect 29596 34290 29652 34300
rect 28812 34242 29428 34244
rect 28812 34190 28814 34242
rect 28866 34190 29428 34242
rect 28812 34188 29428 34190
rect 28812 34178 28868 34188
rect 29372 34132 29428 34188
rect 30828 34242 30884 35308
rect 30940 35026 30996 35038
rect 30940 34974 30942 35026
rect 30994 34974 30996 35026
rect 30940 34804 30996 34974
rect 30940 34738 30996 34748
rect 30828 34190 30830 34242
rect 30882 34190 30884 34242
rect 30828 34178 30884 34190
rect 29596 34132 29652 34142
rect 29372 34130 29652 34132
rect 29372 34078 29598 34130
rect 29650 34078 29652 34130
rect 29372 34076 29652 34078
rect 29596 34066 29652 34076
rect 29708 34132 29764 34142
rect 28700 33964 28980 34020
rect 28252 33518 28254 33570
rect 28306 33518 28308 33570
rect 28252 33506 28308 33518
rect 27916 33346 28196 33348
rect 27916 33294 27918 33346
rect 27970 33294 28196 33346
rect 27916 33292 28196 33294
rect 27916 32676 27972 33292
rect 27916 32610 27972 32620
rect 28700 32564 28756 32574
rect 28252 32508 28700 32564
rect 27804 32452 27860 32462
rect 27468 32162 27524 32172
rect 27692 32450 27860 32452
rect 27692 32398 27806 32450
rect 27858 32398 27860 32450
rect 27692 32396 27860 32398
rect 27468 30994 27524 31006
rect 27468 30942 27470 30994
rect 27522 30942 27524 30994
rect 27468 30884 27524 30942
rect 27580 30884 27636 30894
rect 27468 30828 27580 30884
rect 27580 30818 27636 30828
rect 27468 30210 27524 30222
rect 27468 30158 27470 30210
rect 27522 30158 27524 30210
rect 27468 29428 27524 30158
rect 27468 29362 27524 29372
rect 27580 29314 27636 29326
rect 27580 29262 27582 29314
rect 27634 29262 27636 29314
rect 27356 29148 27524 29204
rect 26236 28914 26292 28924
rect 26236 28754 26292 28766
rect 26236 28702 26238 28754
rect 26290 28702 26292 28754
rect 26236 27860 26292 28702
rect 26460 28644 26516 28654
rect 25900 27858 26292 27860
rect 25900 27806 25902 27858
rect 25954 27806 26292 27858
rect 25900 27804 26292 27806
rect 26348 28642 26516 28644
rect 26348 28590 26462 28642
rect 26514 28590 26516 28642
rect 26348 28588 26516 28590
rect 26348 27970 26404 28588
rect 26460 28578 26516 28588
rect 26684 28644 26740 28654
rect 26684 28550 26740 28588
rect 27020 28642 27076 28654
rect 27020 28590 27022 28642
rect 27074 28590 27076 28642
rect 26348 27918 26350 27970
rect 26402 27918 26404 27970
rect 25900 27794 25956 27804
rect 25564 27746 25732 27748
rect 25564 27694 25566 27746
rect 25618 27694 25732 27746
rect 25564 27692 25732 27694
rect 25564 27682 25620 27692
rect 26348 27074 26404 27918
rect 26908 28532 26964 28542
rect 26796 27860 26852 27870
rect 26460 27636 26516 27646
rect 26460 27186 26516 27580
rect 26460 27134 26462 27186
rect 26514 27134 26516 27186
rect 26460 27122 26516 27134
rect 26572 27634 26628 27646
rect 26572 27582 26574 27634
rect 26626 27582 26628 27634
rect 26348 27022 26350 27074
rect 26402 27022 26404 27074
rect 26348 27010 26404 27022
rect 26572 27074 26628 27582
rect 26572 27022 26574 27074
rect 26626 27022 26628 27074
rect 25452 26852 25620 26908
rect 25228 25106 25284 25116
rect 25452 26178 25508 26190
rect 25452 26126 25454 26178
rect 25506 26126 25508 26178
rect 25228 24724 25284 24734
rect 25452 24724 25508 26126
rect 25564 25956 25620 26852
rect 26572 26740 26628 27022
rect 26796 26964 26852 27804
rect 26908 27634 26964 28476
rect 26908 27582 26910 27634
rect 26962 27582 26964 27634
rect 26908 27570 26964 27582
rect 27020 27636 27076 28590
rect 27132 28644 27188 28654
rect 27132 27748 27188 28588
rect 27244 27972 27300 27982
rect 27244 27878 27300 27916
rect 27356 27858 27412 27870
rect 27356 27806 27358 27858
rect 27410 27806 27412 27858
rect 27244 27748 27300 27758
rect 27132 27746 27300 27748
rect 27132 27694 27246 27746
rect 27298 27694 27300 27746
rect 27132 27692 27300 27694
rect 27244 27682 27300 27692
rect 27020 27570 27076 27580
rect 27356 27188 27412 27806
rect 27356 27122 27412 27132
rect 27468 27186 27524 29148
rect 27580 28868 27636 29262
rect 27692 29204 27748 32396
rect 27804 32386 27860 32396
rect 27692 29138 27748 29148
rect 27804 32228 27860 32238
rect 27804 28980 27860 32172
rect 28028 31778 28084 31790
rect 28028 31726 28030 31778
rect 28082 31726 28084 31778
rect 28028 31106 28084 31726
rect 28252 31218 28308 32508
rect 28700 32470 28756 32508
rect 28588 31668 28644 31678
rect 28588 31574 28644 31612
rect 28924 31332 28980 33964
rect 29708 34018 29764 34076
rect 29708 33966 29710 34018
rect 29762 33966 29764 34018
rect 29708 33954 29764 33966
rect 31052 33570 31108 36316
rect 31164 35698 31220 36540
rect 31836 36372 31892 36382
rect 31164 35646 31166 35698
rect 31218 35646 31220 35698
rect 31164 35634 31220 35646
rect 31724 36370 31892 36372
rect 31724 36318 31838 36370
rect 31890 36318 31892 36370
rect 31724 36316 31892 36318
rect 31612 35588 31668 35598
rect 31612 35494 31668 35532
rect 31276 35028 31332 35038
rect 31052 33518 31054 33570
rect 31106 33518 31108 33570
rect 31052 33506 31108 33518
rect 31164 34972 31276 35028
rect 29708 33458 29764 33470
rect 30828 33460 30884 33470
rect 29708 33406 29710 33458
rect 29762 33406 29764 33458
rect 29372 33346 29428 33358
rect 29372 33294 29374 33346
rect 29426 33294 29428 33346
rect 29148 33234 29204 33246
rect 29148 33182 29150 33234
rect 29202 33182 29204 33234
rect 29148 32564 29204 33182
rect 29148 32498 29204 32508
rect 29260 33124 29316 33134
rect 29372 33124 29428 33294
rect 29708 33348 29764 33406
rect 30716 33458 30884 33460
rect 30716 33406 30830 33458
rect 30882 33406 30884 33458
rect 30716 33404 30884 33406
rect 30156 33348 30212 33358
rect 29708 33346 30212 33348
rect 29708 33294 30158 33346
rect 30210 33294 30212 33346
rect 29708 33292 30212 33294
rect 30156 33282 30212 33292
rect 29316 33068 29428 33124
rect 29260 32450 29316 33068
rect 29596 32676 29652 32686
rect 29596 32582 29652 32620
rect 30716 32676 30772 33404
rect 30828 33394 30884 33404
rect 29260 32398 29262 32450
rect 29314 32398 29316 32450
rect 29260 32386 29316 32398
rect 30604 32562 30660 32574
rect 30604 32510 30606 32562
rect 30658 32510 30660 32562
rect 30604 32228 30660 32510
rect 30716 32450 30772 32620
rect 30716 32398 30718 32450
rect 30770 32398 30772 32450
rect 30716 32386 30772 32398
rect 30940 33346 30996 33358
rect 30940 33294 30942 33346
rect 30994 33294 30996 33346
rect 30940 32340 30996 33294
rect 30828 32284 30996 32340
rect 30828 32228 30884 32284
rect 30604 32172 30884 32228
rect 30492 31778 30548 31790
rect 30492 31726 30494 31778
rect 30546 31726 30548 31778
rect 29148 31668 29204 31678
rect 29148 31574 29204 31612
rect 30380 31666 30436 31678
rect 30380 31614 30382 31666
rect 30434 31614 30436 31666
rect 29260 31556 29316 31566
rect 29260 31462 29316 31500
rect 29484 31556 29540 31566
rect 30380 31556 30436 31614
rect 29484 31554 29764 31556
rect 29484 31502 29486 31554
rect 29538 31502 29764 31554
rect 29484 31500 29764 31502
rect 29484 31490 29540 31500
rect 28924 31266 28980 31276
rect 28252 31166 28254 31218
rect 28306 31166 28308 31218
rect 28252 31154 28308 31166
rect 28028 31054 28030 31106
rect 28082 31054 28084 31106
rect 28028 30322 28084 31054
rect 28252 30994 28308 31006
rect 28252 30942 28254 30994
rect 28306 30942 28308 30994
rect 28252 30884 28308 30942
rect 28252 30818 28308 30828
rect 28476 30994 28532 31006
rect 28476 30942 28478 30994
rect 28530 30942 28532 30994
rect 28028 30270 28030 30322
rect 28082 30270 28084 30322
rect 28028 30258 28084 30270
rect 28476 29650 28532 30942
rect 28700 30996 28756 31006
rect 28700 30212 28756 30940
rect 29708 30994 29764 31500
rect 30156 31220 30212 31230
rect 30156 31106 30212 31164
rect 30156 31054 30158 31106
rect 30210 31054 30212 31106
rect 30156 31042 30212 31054
rect 29708 30942 29710 30994
rect 29762 30942 29764 30994
rect 29708 30930 29764 30942
rect 29484 30882 29540 30894
rect 29484 30830 29486 30882
rect 29538 30830 29540 30882
rect 29484 30212 29540 30830
rect 30380 30772 30436 31500
rect 30492 31668 30548 31726
rect 30492 31108 30548 31612
rect 30604 31218 30660 32172
rect 30604 31166 30606 31218
rect 30658 31166 30660 31218
rect 30604 31154 30660 31166
rect 30492 31042 30548 31052
rect 31164 31106 31220 34972
rect 31276 34962 31332 34972
rect 31388 34916 31444 34926
rect 31276 34804 31332 34814
rect 31276 34130 31332 34748
rect 31276 34078 31278 34130
rect 31330 34078 31332 34130
rect 31276 34066 31332 34078
rect 31388 34132 31444 34860
rect 31724 34804 31780 36316
rect 31836 36306 31892 36316
rect 31948 36258 32004 36270
rect 31948 36206 31950 36258
rect 32002 36206 32004 36258
rect 31948 35924 32004 36206
rect 31836 35868 32004 35924
rect 32172 36258 32228 36270
rect 32172 36206 32174 36258
rect 32226 36206 32228 36258
rect 32172 35924 32228 36206
rect 32284 36036 32340 37996
rect 32396 37044 32452 38444
rect 32732 37940 32788 37950
rect 32732 37846 32788 37884
rect 33740 37492 33796 37502
rect 32508 37268 32564 37278
rect 32508 37174 32564 37212
rect 33516 37268 33572 37278
rect 33516 37174 33572 37212
rect 32396 36988 32564 37044
rect 32396 36372 32452 36382
rect 32396 36278 32452 36316
rect 32284 35980 32452 36036
rect 31836 35476 31892 35868
rect 32172 35858 32228 35868
rect 32284 35812 32340 35822
rect 32284 35718 32340 35756
rect 31948 35700 32004 35710
rect 31948 35606 32004 35644
rect 31836 35420 32004 35476
rect 31948 34916 32004 35420
rect 31948 34850 32004 34860
rect 32396 34914 32452 35980
rect 32396 34862 32398 34914
rect 32450 34862 32452 34914
rect 31724 34738 31780 34748
rect 32396 34804 32452 34862
rect 32396 34738 32452 34748
rect 32508 34580 32564 36988
rect 32956 36484 33012 36494
rect 32956 36390 33012 36428
rect 33628 36484 33684 36494
rect 33628 36390 33684 36428
rect 33180 36372 33236 36382
rect 33180 35586 33236 36316
rect 33516 35924 33572 35934
rect 33516 35810 33572 35868
rect 33516 35758 33518 35810
rect 33570 35758 33572 35810
rect 33516 35746 33572 35758
rect 33180 35534 33182 35586
rect 33234 35534 33236 35586
rect 33180 35522 33236 35534
rect 32732 35028 32788 35038
rect 32732 34914 32788 34972
rect 32732 34862 32734 34914
rect 32786 34862 32788 34914
rect 32732 34850 32788 34862
rect 33292 35028 33348 35038
rect 32844 34692 32900 34702
rect 32844 34598 32900 34636
rect 32956 34690 33012 34702
rect 32956 34638 32958 34690
rect 33010 34638 33012 34690
rect 32060 34524 32564 34580
rect 31500 34132 31556 34142
rect 31388 34130 31556 34132
rect 31388 34078 31502 34130
rect 31554 34078 31556 34130
rect 31388 34076 31556 34078
rect 31500 34066 31556 34076
rect 32060 34020 32116 34524
rect 32172 34244 32228 34254
rect 32956 34244 33012 34638
rect 32172 34242 33012 34244
rect 32172 34190 32174 34242
rect 32226 34190 33012 34242
rect 32172 34188 33012 34190
rect 32172 34178 32228 34188
rect 32956 34130 33012 34188
rect 32956 34078 32958 34130
rect 33010 34078 33012 34130
rect 32956 34066 33012 34078
rect 33292 34130 33348 34972
rect 33404 34804 33460 34814
rect 33404 34710 33460 34748
rect 33292 34078 33294 34130
rect 33346 34078 33348 34130
rect 33292 34066 33348 34078
rect 33516 34692 33572 34702
rect 33516 34130 33572 34636
rect 33516 34078 33518 34130
rect 33570 34078 33572 34130
rect 33516 34066 33572 34078
rect 32060 33964 32228 34020
rect 32060 33348 32116 33358
rect 32060 33254 32116 33292
rect 31500 33236 31556 33246
rect 31500 32786 31556 33180
rect 31500 32734 31502 32786
rect 31554 32734 31556 32786
rect 31500 32722 31556 32734
rect 31164 31054 31166 31106
rect 31218 31054 31220 31106
rect 31164 31042 31220 31054
rect 31612 31778 31668 31790
rect 31612 31726 31614 31778
rect 31666 31726 31668 31778
rect 31612 31220 31668 31726
rect 31836 31220 31892 31230
rect 30828 30996 30884 31006
rect 30828 30902 30884 30940
rect 30380 30706 30436 30716
rect 31388 30772 31444 30782
rect 31388 30322 31444 30716
rect 31388 30270 31390 30322
rect 31442 30270 31444 30322
rect 31388 30258 31444 30270
rect 31612 30324 31668 31164
rect 31724 31164 31836 31220
rect 31724 30994 31780 31164
rect 31836 31154 31892 31164
rect 31724 30942 31726 30994
rect 31778 30942 31780 30994
rect 31724 30930 31780 30942
rect 31836 30884 31892 30894
rect 31836 30790 31892 30828
rect 31948 30324 32004 30334
rect 31612 30322 32004 30324
rect 31612 30270 31950 30322
rect 32002 30270 32004 30322
rect 31612 30268 32004 30270
rect 31948 30258 32004 30268
rect 30380 30212 30436 30222
rect 29484 30156 29764 30212
rect 28476 29598 28478 29650
rect 28530 29598 28532 29650
rect 28476 29586 28532 29598
rect 28588 29986 28644 29998
rect 28588 29934 28590 29986
rect 28642 29934 28644 29986
rect 28588 29652 28644 29934
rect 28588 29586 28644 29596
rect 27916 29540 27972 29550
rect 27916 29426 27972 29484
rect 27916 29374 27918 29426
rect 27970 29374 27972 29426
rect 27916 29362 27972 29374
rect 28588 29428 28644 29438
rect 28140 29316 28196 29326
rect 28140 29222 28196 29260
rect 27580 28802 27636 28812
rect 27692 28924 27860 28980
rect 27580 27860 27636 27870
rect 27580 27766 27636 27804
rect 27468 27134 27470 27186
rect 27522 27134 27524 27186
rect 27468 27122 27524 27134
rect 26796 26962 26964 26964
rect 26796 26910 26798 26962
rect 26850 26910 26964 26962
rect 26796 26908 26964 26910
rect 26796 26898 26852 26908
rect 26572 26674 26628 26684
rect 26908 26628 26964 26908
rect 27244 26962 27300 26974
rect 27244 26910 27246 26962
rect 27298 26910 27300 26962
rect 27244 26908 27300 26910
rect 27244 26852 27412 26908
rect 26908 26562 26964 26572
rect 26684 26516 26740 26526
rect 26684 26422 26740 26460
rect 26236 26404 26292 26414
rect 26236 26310 26292 26348
rect 26572 26290 26628 26302
rect 26572 26238 26574 26290
rect 26626 26238 26628 26290
rect 25788 26180 25844 26190
rect 25788 26086 25844 26124
rect 26572 26180 26628 26238
rect 26796 26292 26852 26302
rect 26796 26290 27076 26292
rect 26796 26238 26798 26290
rect 26850 26238 27076 26290
rect 26796 26236 27076 26238
rect 26796 26226 26852 26236
rect 25564 25900 26292 25956
rect 26236 25730 26292 25900
rect 26236 25678 26238 25730
rect 26290 25678 26292 25730
rect 26236 25666 26292 25678
rect 26012 25508 26068 25518
rect 26012 25414 26068 25452
rect 26236 25508 26292 25518
rect 25900 24948 25956 24958
rect 25284 24668 25508 24724
rect 25788 24892 25900 24948
rect 25228 24630 25284 24668
rect 24668 23214 24670 23266
rect 24722 23214 24724 23266
rect 24668 23202 24724 23214
rect 25004 23938 25060 23950
rect 25004 23886 25006 23938
rect 25058 23886 25060 23938
rect 24332 23102 24334 23154
rect 24386 23102 24388 23154
rect 24332 23090 24388 23102
rect 24556 22932 24612 22942
rect 24556 22838 24612 22876
rect 24444 22482 24500 22494
rect 24444 22430 24446 22482
rect 24498 22430 24500 22482
rect 24444 22148 24500 22430
rect 24892 22148 24948 22158
rect 24444 22082 24500 22092
rect 24780 22146 24948 22148
rect 24780 22094 24894 22146
rect 24946 22094 24948 22146
rect 24780 22092 24948 22094
rect 24332 21924 24388 21934
rect 24220 21868 24332 21924
rect 24332 21810 24388 21868
rect 24332 21758 24334 21810
rect 24386 21758 24388 21810
rect 24332 21746 24388 21758
rect 23996 21646 23998 21698
rect 24050 21646 24052 21698
rect 23996 21634 24052 21646
rect 23884 21586 23940 21598
rect 23884 21534 23886 21586
rect 23938 21534 23940 21586
rect 23884 21476 23940 21534
rect 23884 21410 23940 21420
rect 24556 21586 24612 21598
rect 24556 21534 24558 21586
rect 24610 21534 24612 21586
rect 24556 21364 24612 21534
rect 24556 21298 24612 21308
rect 24780 21140 24836 22092
rect 24892 22082 24948 22092
rect 23772 20710 23828 20748
rect 24332 21084 24836 21140
rect 24892 21924 24948 21934
rect 24108 20692 24164 20702
rect 23996 20690 24164 20692
rect 23996 20638 24110 20690
rect 24162 20638 24164 20690
rect 23996 20636 24164 20638
rect 23996 20188 24052 20636
rect 24108 20626 24164 20636
rect 24220 20692 24276 20702
rect 24220 20598 24276 20636
rect 23436 20132 23604 20188
rect 23548 19906 23604 20132
rect 23548 19854 23550 19906
rect 23602 19854 23604 19906
rect 23548 19796 23604 19854
rect 23548 19730 23604 19740
rect 23660 20132 24052 20188
rect 24108 20132 24164 20142
rect 23660 19460 23716 20132
rect 24108 20130 24276 20132
rect 24108 20078 24110 20130
rect 24162 20078 24276 20130
rect 24108 20076 24276 20078
rect 24108 20066 24164 20076
rect 23884 20020 23940 20030
rect 23884 20018 24052 20020
rect 23884 19966 23886 20018
rect 23938 19966 24052 20018
rect 23884 19964 24052 19966
rect 23884 19954 23940 19964
rect 23212 19394 23268 19404
rect 23548 19404 23716 19460
rect 23100 19070 23102 19122
rect 23154 19070 23156 19122
rect 23100 19058 23156 19070
rect 23324 19234 23380 19246
rect 23324 19182 23326 19234
rect 23378 19182 23380 19234
rect 23324 18452 23380 19182
rect 23436 18788 23492 18798
rect 23548 18788 23604 19404
rect 23492 18732 23604 18788
rect 23660 19236 23716 19246
rect 23436 18722 23492 18732
rect 23324 18358 23380 18396
rect 23548 18562 23604 18574
rect 23548 18510 23550 18562
rect 23602 18510 23604 18562
rect 23548 18228 23604 18510
rect 23548 18162 23604 18172
rect 23100 18116 23156 18126
rect 23156 18060 23268 18116
rect 23100 18050 23156 18060
rect 22988 16818 23044 16828
rect 23100 17666 23156 17678
rect 23100 17614 23102 17666
rect 23154 17614 23156 17666
rect 22764 16716 22932 16772
rect 22764 16212 22820 16716
rect 22988 16660 23044 16670
rect 21980 16156 22260 16212
rect 22316 16156 22484 16212
rect 21756 15988 21812 15998
rect 21756 15894 21812 15932
rect 21980 15874 22036 16156
rect 21980 15822 21982 15874
rect 22034 15822 22036 15874
rect 21980 15810 22036 15822
rect 22092 15986 22148 15998
rect 22092 15934 22094 15986
rect 22146 15934 22148 15986
rect 21644 15708 21812 15764
rect 21644 15202 21700 15214
rect 21644 15150 21646 15202
rect 21698 15150 21700 15202
rect 21644 14980 21700 15150
rect 21644 14914 21700 14924
rect 21756 14644 21812 15708
rect 21308 14530 21588 14532
rect 21308 14478 21310 14530
rect 21362 14478 21588 14530
rect 21308 14476 21588 14478
rect 21644 14588 21812 14644
rect 22092 14644 22148 15934
rect 21308 14466 21364 14476
rect 21420 14308 21476 14318
rect 21196 14306 21476 14308
rect 21196 14254 21422 14306
rect 21474 14254 21476 14306
rect 21196 14252 21476 14254
rect 21196 14084 21252 14094
rect 21196 12290 21252 14028
rect 21196 12238 21198 12290
rect 21250 12238 21252 12290
rect 21196 12226 21252 12238
rect 21308 12402 21364 14252
rect 21420 14242 21476 14252
rect 21308 12350 21310 12402
rect 21362 12350 21364 12402
rect 21308 11956 21364 12350
rect 21084 10994 21140 11004
rect 21196 11900 21364 11956
rect 21420 13746 21476 13758
rect 21420 13694 21422 13746
rect 21474 13694 21476 13746
rect 21420 13524 21476 13694
rect 21532 13748 21588 13758
rect 21532 13654 21588 13692
rect 21644 13524 21700 14588
rect 22092 14578 22148 14588
rect 22204 14642 22260 16156
rect 22204 14590 22206 14642
rect 22258 14590 22260 14642
rect 22204 14578 22260 14590
rect 22316 15986 22372 15998
rect 22316 15934 22318 15986
rect 22370 15934 22372 15986
rect 22316 14980 22372 15934
rect 22428 15764 22484 16156
rect 22764 16146 22820 16156
rect 22876 16658 23044 16660
rect 22876 16606 22990 16658
rect 23042 16606 23044 16658
rect 22876 16604 23044 16606
rect 22428 15698 22484 15708
rect 21756 14420 21812 14430
rect 21756 13972 21812 14364
rect 22092 14084 22148 14094
rect 21756 13916 21924 13972
rect 21196 10948 21252 11900
rect 21308 11732 21364 11742
rect 21308 11506 21364 11676
rect 21420 11620 21476 13468
rect 21532 13468 21700 13524
rect 21756 13746 21812 13758
rect 21756 13694 21758 13746
rect 21810 13694 21812 13746
rect 21532 12402 21588 13468
rect 21644 13076 21700 13086
rect 21756 13076 21812 13694
rect 21700 13020 21812 13076
rect 21644 13010 21700 13020
rect 21532 12350 21534 12402
rect 21586 12350 21588 12402
rect 21532 12338 21588 12350
rect 21644 12850 21700 12862
rect 21644 12798 21646 12850
rect 21698 12798 21700 12850
rect 21644 12740 21700 12798
rect 21756 12852 21812 12862
rect 21756 12758 21812 12796
rect 21532 11844 21588 11854
rect 21644 11844 21700 12684
rect 21868 12178 21924 13916
rect 21868 12126 21870 12178
rect 21922 12126 21924 12178
rect 21868 12114 21924 12126
rect 21980 13746 22036 13758
rect 21980 13694 21982 13746
rect 22034 13694 22036 13746
rect 21980 12850 22036 13694
rect 21980 12798 21982 12850
rect 22034 12798 22036 12850
rect 21588 11788 21700 11844
rect 21980 11844 22036 12798
rect 21532 11778 21588 11788
rect 21980 11778 22036 11788
rect 22092 13636 22148 14028
rect 22316 13860 22372 14924
rect 22876 14756 22932 16604
rect 22988 16594 23044 16604
rect 23100 16436 23156 17614
rect 23212 16772 23268 18060
rect 23660 17668 23716 19180
rect 23884 19234 23940 19246
rect 23884 19182 23886 19234
rect 23938 19182 23940 19234
rect 23772 19124 23828 19134
rect 23772 17890 23828 19068
rect 23884 18676 23940 19182
rect 23884 18610 23940 18620
rect 23996 18564 24052 19964
rect 23884 18452 23940 18462
rect 23996 18452 24052 18508
rect 23884 18450 24052 18452
rect 23884 18398 23886 18450
rect 23938 18398 24052 18450
rect 23884 18396 24052 18398
rect 24108 19348 24164 19358
rect 24108 18674 24164 19292
rect 24108 18622 24110 18674
rect 24162 18622 24164 18674
rect 23884 18386 23940 18396
rect 23884 18228 23940 18238
rect 23940 18172 24052 18228
rect 23884 18162 23940 18172
rect 23772 17838 23774 17890
rect 23826 17838 23828 17890
rect 23772 17826 23828 17838
rect 23884 17668 23940 17678
rect 23660 17666 23940 17668
rect 23660 17614 23886 17666
rect 23938 17614 23940 17666
rect 23660 17612 23940 17614
rect 23884 17602 23940 17612
rect 23324 17556 23380 17566
rect 23436 17556 23492 17566
rect 23324 17554 23436 17556
rect 23324 17502 23326 17554
rect 23378 17502 23436 17554
rect 23324 17500 23436 17502
rect 23492 17500 23716 17556
rect 23324 17490 23380 17500
rect 23436 17462 23492 17500
rect 23436 16882 23492 16894
rect 23436 16830 23438 16882
rect 23490 16830 23492 16882
rect 23212 16770 23380 16772
rect 23212 16718 23214 16770
rect 23266 16718 23380 16770
rect 23212 16716 23380 16718
rect 23212 16706 23268 16716
rect 23100 16098 23156 16380
rect 23324 16324 23380 16716
rect 23436 16660 23492 16830
rect 23548 16660 23604 16670
rect 23436 16604 23548 16660
rect 23548 16594 23604 16604
rect 23324 16258 23380 16268
rect 23100 16046 23102 16098
rect 23154 16046 23156 16098
rect 23100 16034 23156 16046
rect 23436 16210 23492 16222
rect 23436 16158 23438 16210
rect 23490 16158 23492 16210
rect 21476 11564 21588 11620
rect 21420 11554 21476 11564
rect 21308 11454 21310 11506
rect 21362 11454 21364 11506
rect 21308 11442 21364 11454
rect 21532 11506 21588 11564
rect 21532 11454 21534 11506
rect 21586 11454 21588 11506
rect 21532 11442 21588 11454
rect 21644 11508 21700 11518
rect 21700 11452 21812 11508
rect 21644 11442 21700 11452
rect 21196 10882 21252 10892
rect 20972 10610 21028 10622
rect 20972 10558 20974 10610
rect 21026 10558 21028 10610
rect 20972 10276 21028 10558
rect 21084 10612 21140 10622
rect 21084 10518 21140 10556
rect 21196 10610 21252 10622
rect 21196 10558 21198 10610
rect 21250 10558 21252 10610
rect 21196 10388 21252 10558
rect 21644 10388 21700 10398
rect 21196 10322 21252 10332
rect 21532 10386 21700 10388
rect 21532 10334 21646 10386
rect 21698 10334 21700 10386
rect 21532 10332 21700 10334
rect 20972 10210 21028 10220
rect 20860 8642 20916 8652
rect 21084 9940 21140 9950
rect 21084 8484 21140 9884
rect 21420 9044 21476 9054
rect 21420 8930 21476 8988
rect 21420 8878 21422 8930
rect 21474 8878 21476 8930
rect 21420 8866 21476 8878
rect 21084 8418 21140 8428
rect 21532 8372 21588 10332
rect 21644 10322 21700 10332
rect 21644 10164 21700 10174
rect 21644 9938 21700 10108
rect 21644 9886 21646 9938
rect 21698 9886 21700 9938
rect 21644 9874 21700 9886
rect 21756 9268 21812 11452
rect 21868 11172 21924 11182
rect 21868 11170 22036 11172
rect 21868 11118 21870 11170
rect 21922 11118 22036 11170
rect 21868 11116 22036 11118
rect 21868 11106 21924 11116
rect 21868 10724 21924 10734
rect 21868 10610 21924 10668
rect 21868 10558 21870 10610
rect 21922 10558 21924 10610
rect 21868 10386 21924 10558
rect 21868 10334 21870 10386
rect 21922 10334 21924 10386
rect 21868 10322 21924 10334
rect 21980 10498 22036 11116
rect 22092 10948 22148 13580
rect 22204 13804 22372 13860
rect 22428 14700 22932 14756
rect 22204 13412 22260 13804
rect 22316 13636 22372 13646
rect 22316 13542 22372 13580
rect 22204 13356 22372 13412
rect 22204 12850 22260 12862
rect 22204 12798 22206 12850
rect 22258 12798 22260 12850
rect 22204 11618 22260 12798
rect 22316 11732 22372 13356
rect 22428 13188 22484 14700
rect 22540 14530 22596 14542
rect 22540 14478 22542 14530
rect 22594 14478 22596 14530
rect 22540 13972 22596 14478
rect 22988 14420 23044 14430
rect 23324 14420 23380 14430
rect 22988 14418 23380 14420
rect 22988 14366 22990 14418
rect 23042 14366 23326 14418
rect 23378 14366 23380 14418
rect 22988 14364 23380 14366
rect 22988 14354 23044 14364
rect 23324 14354 23380 14364
rect 23436 14420 23492 16158
rect 23660 15148 23716 17500
rect 23772 17444 23828 17454
rect 23996 17444 24052 18172
rect 24108 17556 24164 18622
rect 24220 18004 24276 20076
rect 24332 20018 24388 21084
rect 24332 19966 24334 20018
rect 24386 19966 24388 20018
rect 24332 19954 24388 19966
rect 24444 20130 24500 20142
rect 24444 20078 24446 20130
rect 24498 20078 24500 20130
rect 24332 19796 24388 19806
rect 24332 18450 24388 19740
rect 24444 19684 24500 20078
rect 24444 19618 24500 19628
rect 24668 19906 24724 19918
rect 24668 19854 24670 19906
rect 24722 19854 24724 19906
rect 24556 19348 24612 19358
rect 24668 19348 24724 19854
rect 24556 19346 24724 19348
rect 24556 19294 24558 19346
rect 24610 19294 24724 19346
rect 24556 19292 24724 19294
rect 24780 19460 24836 19470
rect 24556 19282 24612 19292
rect 24444 18564 24500 18574
rect 24444 18470 24500 18508
rect 24332 18398 24334 18450
rect 24386 18398 24388 18450
rect 24332 18386 24388 18398
rect 24668 18340 24724 18350
rect 24668 18246 24724 18284
rect 24780 18228 24836 19404
rect 24892 18340 24948 21868
rect 25004 20580 25060 23886
rect 25340 23604 25396 23614
rect 25340 22484 25396 23548
rect 25340 22418 25396 22428
rect 25564 23154 25620 23166
rect 25564 23102 25566 23154
rect 25618 23102 25620 23154
rect 25116 22372 25172 22382
rect 25116 22146 25172 22316
rect 25452 22372 25508 22382
rect 25228 22260 25284 22270
rect 25228 22166 25284 22204
rect 25116 22094 25118 22146
rect 25170 22094 25172 22146
rect 25116 22082 25172 22094
rect 25228 21812 25284 21822
rect 25116 21700 25172 21710
rect 25228 21700 25284 21756
rect 25340 21812 25396 21822
rect 25452 21812 25508 22316
rect 25564 22148 25620 23102
rect 25564 22082 25620 22092
rect 25340 21810 25620 21812
rect 25340 21758 25342 21810
rect 25394 21758 25620 21810
rect 25340 21756 25620 21758
rect 25340 21746 25396 21756
rect 25116 21698 25284 21700
rect 25116 21646 25118 21698
rect 25170 21646 25284 21698
rect 25116 21644 25284 21646
rect 25564 21700 25620 21756
rect 25564 21644 25732 21700
rect 25116 21634 25172 21644
rect 25452 21586 25508 21598
rect 25452 21534 25454 21586
rect 25506 21534 25508 21586
rect 25452 21140 25508 21534
rect 25452 21074 25508 21084
rect 25564 20916 25620 20926
rect 25340 20804 25396 20814
rect 25396 20748 25508 20804
rect 25340 20710 25396 20748
rect 25004 20514 25060 20524
rect 25116 20244 25172 20254
rect 25452 20244 25508 20748
rect 25564 20802 25620 20860
rect 25564 20750 25566 20802
rect 25618 20750 25620 20802
rect 25564 20356 25620 20750
rect 25564 20290 25620 20300
rect 25172 20188 25284 20244
rect 25116 20178 25172 20188
rect 25228 20130 25284 20188
rect 25452 20178 25508 20188
rect 25228 20078 25230 20130
rect 25282 20078 25284 20130
rect 25228 20066 25284 20078
rect 25340 20132 25396 20142
rect 25340 20038 25396 20076
rect 25340 19796 25396 19806
rect 25340 19702 25396 19740
rect 25116 18676 25172 18686
rect 25116 18452 25172 18620
rect 25340 18452 25396 18462
rect 25116 18450 25396 18452
rect 25116 18398 25342 18450
rect 25394 18398 25396 18450
rect 25116 18396 25396 18398
rect 24892 18284 25172 18340
rect 24780 18172 25060 18228
rect 24220 17938 24276 17948
rect 24780 18004 24836 18014
rect 24836 17948 24948 18004
rect 24780 17938 24836 17948
rect 24668 17668 24724 17678
rect 24108 17490 24164 17500
rect 24444 17612 24668 17668
rect 24332 17444 24388 17454
rect 23772 17442 24052 17444
rect 23772 17390 23774 17442
rect 23826 17390 24052 17442
rect 23772 17388 24052 17390
rect 24220 17442 24388 17444
rect 24220 17390 24334 17442
rect 24386 17390 24388 17442
rect 24220 17388 24388 17390
rect 23772 17378 23828 17388
rect 23772 16884 23828 16894
rect 23772 16790 23828 16828
rect 23884 16436 23940 17388
rect 24220 16884 24276 17388
rect 24332 17378 24388 17388
rect 24332 17108 24388 17118
rect 24332 17014 24388 17052
rect 24220 16828 24388 16884
rect 23772 16380 23940 16436
rect 24108 16660 24164 16670
rect 23772 15764 23828 16380
rect 23884 16212 23940 16222
rect 23884 16118 23940 16156
rect 23772 15698 23828 15708
rect 23996 15986 24052 15998
rect 23996 15934 23998 15986
rect 24050 15934 24052 15986
rect 23996 15540 24052 15934
rect 23884 15484 24052 15540
rect 23548 15092 23716 15148
rect 23772 15202 23828 15214
rect 23772 15150 23774 15202
rect 23826 15150 23828 15202
rect 23548 14532 23604 15092
rect 23660 14756 23716 14766
rect 23772 14756 23828 15150
rect 23884 15148 23940 15484
rect 23884 15092 24052 15148
rect 23660 14754 23828 14756
rect 23660 14702 23662 14754
rect 23714 14702 23828 14754
rect 23660 14700 23828 14702
rect 23884 14756 23940 14766
rect 23660 14690 23716 14700
rect 23548 14476 23828 14532
rect 23436 14354 23492 14364
rect 23548 14306 23604 14318
rect 23548 14254 23550 14306
rect 23602 14254 23604 14306
rect 23548 14084 23604 14254
rect 23548 14018 23604 14028
rect 23324 13972 23380 13982
rect 22596 13916 22820 13972
rect 22540 13906 22596 13916
rect 22540 13524 22596 13534
rect 22540 13430 22596 13468
rect 22428 13132 22596 13188
rect 22428 12962 22484 12974
rect 22428 12910 22430 12962
rect 22482 12910 22484 12962
rect 22428 12852 22484 12910
rect 22428 12786 22484 12796
rect 22540 12628 22596 13132
rect 22764 12962 22820 13916
rect 22876 13748 22932 13758
rect 23212 13748 23268 13758
rect 22932 13692 23044 13748
rect 22876 13682 22932 13692
rect 22876 13522 22932 13534
rect 22876 13470 22878 13522
rect 22930 13470 22932 13522
rect 22876 13300 22932 13470
rect 22876 13234 22932 13244
rect 22764 12910 22766 12962
rect 22818 12910 22820 12962
rect 22764 12898 22820 12910
rect 22316 11666 22372 11676
rect 22428 12572 22596 12628
rect 22652 12738 22708 12750
rect 22988 12740 23044 13692
rect 23212 13654 23268 13692
rect 23324 13634 23380 13916
rect 23660 13860 23716 13870
rect 23660 13766 23716 13804
rect 23324 13582 23326 13634
rect 23378 13582 23380 13634
rect 23324 13570 23380 13582
rect 23436 13746 23492 13758
rect 23436 13694 23438 13746
rect 23490 13694 23492 13746
rect 23436 13300 23492 13694
rect 23212 13244 23492 13300
rect 23548 13748 23604 13758
rect 22652 12686 22654 12738
rect 22706 12686 22708 12738
rect 22204 11566 22206 11618
rect 22258 11566 22260 11618
rect 22204 11554 22260 11566
rect 22316 11394 22372 11406
rect 22316 11342 22318 11394
rect 22370 11342 22372 11394
rect 22316 11172 22372 11342
rect 22316 11106 22372 11116
rect 22092 10892 22372 10948
rect 21980 10446 21982 10498
rect 22034 10446 22036 10498
rect 21980 10388 22036 10446
rect 21980 10322 22036 10332
rect 22092 10610 22148 10622
rect 22092 10558 22094 10610
rect 22146 10558 22148 10610
rect 22092 10276 22148 10558
rect 22092 9492 22148 10220
rect 21196 8316 21476 8372
rect 21196 8260 21252 8316
rect 21196 8194 21252 8204
rect 20412 8054 20468 8092
rect 21420 8146 21476 8316
rect 21532 8258 21588 8316
rect 21532 8206 21534 8258
rect 21586 8206 21588 8258
rect 21532 8194 21588 8206
rect 21644 9212 21812 9268
rect 21980 9436 22148 9492
rect 21420 8094 21422 8146
rect 21474 8094 21476 8146
rect 21196 8036 21252 8046
rect 20524 8034 21252 8036
rect 20524 7982 21198 8034
rect 21250 7982 21252 8034
rect 20524 7980 21252 7982
rect 21420 8036 21476 8094
rect 21420 7980 21588 8036
rect 20524 7924 20580 7980
rect 21196 7970 21252 7980
rect 20300 7746 20356 7756
rect 20412 7868 20580 7924
rect 21532 7924 21588 7980
rect 20300 7476 20356 7486
rect 20412 7476 20468 7868
rect 21532 7858 21588 7868
rect 20860 7812 20916 7822
rect 20300 7474 20468 7476
rect 20300 7422 20302 7474
rect 20354 7422 20468 7474
rect 20300 7420 20468 7422
rect 20636 7586 20692 7598
rect 20636 7534 20638 7586
rect 20690 7534 20692 7586
rect 20300 7410 20356 7420
rect 20412 7252 20468 7262
rect 20412 7158 20468 7196
rect 20636 7028 20692 7534
rect 19852 6638 19854 6690
rect 19906 6638 19908 6690
rect 19852 6626 19908 6638
rect 20076 6692 20132 6702
rect 20188 6692 20244 6748
rect 20076 6690 20244 6692
rect 20076 6638 20078 6690
rect 20130 6638 20244 6690
rect 20076 6636 20244 6638
rect 20524 6972 20692 7028
rect 20076 6626 20132 6636
rect 19964 6468 20020 6478
rect 20412 6468 20468 6478
rect 20524 6468 20580 6972
rect 19964 6466 20244 6468
rect 19964 6414 19966 6466
rect 20018 6414 20244 6466
rect 19964 6412 20244 6414
rect 19964 6402 20020 6412
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19964 6132 20020 6142
rect 20188 6132 20244 6412
rect 20020 6076 20244 6132
rect 20412 6466 20580 6468
rect 20412 6414 20414 6466
rect 20466 6414 20580 6466
rect 20412 6412 20580 6414
rect 20636 6692 20692 6702
rect 19964 5906 20020 6076
rect 19964 5854 19966 5906
rect 20018 5854 20020 5906
rect 19964 5842 20020 5854
rect 20188 5906 20244 5918
rect 20188 5854 20190 5906
rect 20242 5854 20244 5906
rect 20076 5796 20132 5806
rect 20188 5796 20244 5854
rect 19628 5794 19796 5796
rect 19628 5742 19630 5794
rect 19682 5742 19796 5794
rect 19628 5740 19796 5742
rect 19628 5730 19684 5740
rect 19628 5348 19684 5358
rect 19628 5254 19684 5292
rect 19740 5346 19796 5740
rect 20132 5740 20244 5796
rect 20076 5730 20132 5740
rect 20412 5684 20468 6412
rect 19740 5294 19742 5346
rect 19794 5294 19796 5346
rect 19740 5282 19796 5294
rect 20188 5628 20468 5684
rect 19516 4498 19572 4508
rect 19628 5124 19684 5134
rect 19516 4228 19572 4238
rect 19516 3778 19572 4172
rect 19516 3726 19518 3778
rect 19570 3726 19572 3778
rect 19516 3714 19572 3726
rect 19292 3614 19294 3666
rect 19346 3614 19348 3666
rect 19292 3602 19348 3614
rect 19628 3666 19684 5068
rect 19964 5012 20020 5022
rect 20188 5012 20244 5628
rect 20412 5124 20468 5134
rect 20636 5124 20692 6636
rect 20748 6466 20804 6478
rect 20748 6414 20750 6466
rect 20802 6414 20804 6466
rect 20748 6132 20804 6414
rect 20748 5236 20804 6076
rect 20748 5170 20804 5180
rect 20412 5030 20468 5068
rect 20524 5122 20692 5124
rect 20524 5070 20638 5122
rect 20690 5070 20692 5122
rect 20524 5068 20692 5070
rect 19964 5010 20244 5012
rect 19964 4958 19966 5010
rect 20018 4958 20244 5010
rect 19964 4956 20244 4958
rect 20300 5012 20356 5022
rect 19964 4900 20020 4956
rect 20300 4918 20356 4956
rect 19964 4834 20020 4844
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19628 3614 19630 3666
rect 19682 3614 19684 3666
rect 19628 3602 19684 3614
rect 20076 4564 20132 4574
rect 20076 3666 20132 4508
rect 20412 4228 20468 4238
rect 20524 4228 20580 5068
rect 20636 5058 20692 5068
rect 20748 4340 20804 4350
rect 20748 4246 20804 4284
rect 20412 4226 20580 4228
rect 20412 4174 20414 4226
rect 20466 4174 20580 4226
rect 20412 4172 20580 4174
rect 20412 4162 20468 4172
rect 20076 3614 20078 3666
rect 20130 3614 20132 3666
rect 20076 3602 20132 3614
rect 20860 3668 20916 7756
rect 21420 7812 21476 7822
rect 21084 7588 21140 7598
rect 21084 7494 21140 7532
rect 20972 7474 21028 7486
rect 20972 7422 20974 7474
rect 21026 7422 21028 7474
rect 20972 7364 21028 7422
rect 21196 7474 21252 7486
rect 21420 7476 21476 7756
rect 21196 7422 21198 7474
rect 21250 7422 21252 7474
rect 20972 7308 21140 7364
rect 20972 7140 21028 7150
rect 20972 6130 21028 7084
rect 20972 6078 20974 6130
rect 21026 6078 21028 6130
rect 20972 6066 21028 6078
rect 21084 5012 21140 7308
rect 21196 7252 21252 7422
rect 21196 7186 21252 7196
rect 21308 7420 21476 7476
rect 21644 7700 21700 9212
rect 21756 9042 21812 9054
rect 21756 8990 21758 9042
rect 21810 8990 21812 9042
rect 21756 8148 21812 8990
rect 21868 8932 21924 8942
rect 21868 8838 21924 8876
rect 21980 8260 22036 9436
rect 22316 9380 22372 10892
rect 22428 9604 22484 12572
rect 22540 12292 22596 12302
rect 22652 12292 22708 12686
rect 22540 12290 22708 12292
rect 22540 12238 22542 12290
rect 22594 12238 22708 12290
rect 22540 12236 22708 12238
rect 22764 12684 23044 12740
rect 23100 13188 23156 13198
rect 23100 12850 23156 13132
rect 23100 12798 23102 12850
rect 23154 12798 23156 12850
rect 22540 12226 22596 12236
rect 22652 11620 22708 11630
rect 22540 11564 22652 11620
rect 22540 11506 22596 11564
rect 22652 11554 22708 11564
rect 22540 11454 22542 11506
rect 22594 11454 22596 11506
rect 22540 10386 22596 11454
rect 22764 11394 22820 12684
rect 23100 11844 23156 12798
rect 22764 11342 22766 11394
rect 22818 11342 22820 11394
rect 22764 11330 22820 11342
rect 22988 11788 23156 11844
rect 23212 11788 23268 13244
rect 23436 12964 23492 13002
rect 23436 12898 23492 12908
rect 23548 12850 23604 13692
rect 23772 13636 23828 14476
rect 23884 14530 23940 14700
rect 23884 14478 23886 14530
rect 23938 14478 23940 14530
rect 23884 14466 23940 14478
rect 23884 14308 23940 14318
rect 23884 13970 23940 14252
rect 23884 13918 23886 13970
rect 23938 13918 23940 13970
rect 23884 13906 23940 13918
rect 23996 13860 24052 15092
rect 24108 14418 24164 16604
rect 24220 16100 24276 16110
rect 24220 16006 24276 16044
rect 24332 15988 24388 16828
rect 24332 15922 24388 15932
rect 24444 15986 24500 17612
rect 24668 17574 24724 17612
rect 24556 17444 24612 17454
rect 24556 17106 24612 17388
rect 24556 17054 24558 17106
rect 24610 17054 24612 17106
rect 24556 17042 24612 17054
rect 24668 17220 24724 17230
rect 24668 16994 24724 17164
rect 24668 16942 24670 16994
rect 24722 16942 24724 16994
rect 24668 16930 24724 16942
rect 24780 17108 24836 17118
rect 24780 16884 24836 17052
rect 24780 16548 24836 16828
rect 24444 15934 24446 15986
rect 24498 15934 24500 15986
rect 24444 15922 24500 15934
rect 24556 16492 24836 16548
rect 24556 16098 24612 16492
rect 24892 16436 24948 17948
rect 25004 17666 25060 18172
rect 25004 17614 25006 17666
rect 25058 17614 25060 17666
rect 25004 17602 25060 17614
rect 25116 17444 25172 18284
rect 25116 17378 25172 17388
rect 25228 16772 25284 16782
rect 25228 16678 25284 16716
rect 24556 16046 24558 16098
rect 24610 16046 24612 16098
rect 24556 15764 24612 16046
rect 24780 16380 24948 16436
rect 24220 15708 24612 15764
rect 24668 15764 24724 15774
rect 24220 14530 24276 15708
rect 24220 14478 24222 14530
rect 24274 14478 24276 14530
rect 24220 14466 24276 14478
rect 24332 15540 24388 15550
rect 24108 14366 24110 14418
rect 24162 14366 24164 14418
rect 24108 14354 24164 14366
rect 24108 13860 24164 13870
rect 23996 13858 24164 13860
rect 23996 13806 24110 13858
rect 24162 13806 24164 13858
rect 23996 13804 24164 13806
rect 24108 13748 24164 13804
rect 24108 13682 24164 13692
rect 24220 13748 24276 13758
rect 24332 13748 24388 15484
rect 24444 15314 24500 15326
rect 24444 15262 24446 15314
rect 24498 15262 24500 15314
rect 24444 15204 24500 15262
rect 24668 15148 24724 15708
rect 24444 15138 24500 15148
rect 24220 13746 24388 13748
rect 24220 13694 24222 13746
rect 24274 13694 24388 13746
rect 24220 13692 24388 13694
rect 24556 15092 24724 15148
rect 23772 13580 23940 13636
rect 23772 13412 23828 13422
rect 23772 12962 23828 13356
rect 23772 12910 23774 12962
rect 23826 12910 23828 12962
rect 23772 12898 23828 12910
rect 23548 12798 23550 12850
rect 23602 12798 23604 12850
rect 23548 12786 23604 12798
rect 23660 11844 23716 11854
rect 22988 10836 23044 11788
rect 23212 11732 23380 11788
rect 23100 11620 23156 11630
rect 23324 11620 23380 11732
rect 23156 11564 23380 11620
rect 23436 11732 23492 11742
rect 23100 11526 23156 11564
rect 23324 11396 23380 11406
rect 23324 11282 23380 11340
rect 23324 11230 23326 11282
rect 23378 11230 23380 11282
rect 23324 11218 23380 11230
rect 23212 11170 23268 11182
rect 23212 11118 23214 11170
rect 23266 11118 23268 11170
rect 22988 10780 23156 10836
rect 22988 10612 23044 10622
rect 22988 10518 23044 10556
rect 22540 10334 22542 10386
rect 22594 10334 22596 10386
rect 22540 10322 22596 10334
rect 23100 9716 23156 10780
rect 23212 10724 23268 11118
rect 23324 10724 23380 10734
rect 23212 10722 23380 10724
rect 23212 10670 23326 10722
rect 23378 10670 23380 10722
rect 23212 10668 23380 10670
rect 23324 10658 23380 10668
rect 23100 9650 23156 9660
rect 23212 10276 23268 10286
rect 22428 9538 22484 9548
rect 22316 9324 22708 9380
rect 22092 9156 22148 9166
rect 22092 9062 22148 9100
rect 21756 8082 21812 8092
rect 21868 8204 22036 8260
rect 22204 9044 22260 9054
rect 21196 5796 21252 5806
rect 21196 5124 21252 5740
rect 21196 5058 21252 5068
rect 21084 4946 21140 4956
rect 20972 3668 21028 3678
rect 20860 3666 21028 3668
rect 20860 3614 20974 3666
rect 21026 3614 21028 3666
rect 20860 3612 21028 3614
rect 20972 3602 21028 3612
rect 21308 3388 21364 7420
rect 21532 6692 21588 6702
rect 21644 6692 21700 7644
rect 21532 6690 21700 6692
rect 21532 6638 21534 6690
rect 21586 6638 21700 6690
rect 21532 6636 21700 6638
rect 21756 7588 21812 7598
rect 21868 7588 21924 8204
rect 21980 8036 22036 8046
rect 21980 7942 22036 7980
rect 21980 7588 22036 7598
rect 21868 7586 22036 7588
rect 21868 7534 21982 7586
rect 22034 7534 22036 7586
rect 21868 7532 22036 7534
rect 21756 6804 21812 7532
rect 21980 7522 22036 7532
rect 22204 7474 22260 8988
rect 22652 8370 22708 9324
rect 23212 9154 23268 10220
rect 23324 10164 23380 10174
rect 23436 10164 23492 11676
rect 23548 11620 23604 11630
rect 23548 11172 23604 11564
rect 23548 11106 23604 11116
rect 23548 10388 23604 10398
rect 23548 10294 23604 10332
rect 23436 10108 23604 10164
rect 23324 9266 23380 10108
rect 23324 9214 23326 9266
rect 23378 9214 23380 9266
rect 23324 9202 23380 9214
rect 23436 9716 23492 9726
rect 23212 9102 23214 9154
rect 23266 9102 23268 9154
rect 23212 9090 23268 9102
rect 22764 8932 22820 8942
rect 23436 8932 23492 9660
rect 22764 8930 23044 8932
rect 22764 8878 22766 8930
rect 22818 8878 23044 8930
rect 22764 8876 23044 8878
rect 22764 8866 22820 8876
rect 22764 8708 22820 8718
rect 22820 8652 22932 8708
rect 22764 8642 22820 8652
rect 22652 8318 22654 8370
rect 22706 8318 22708 8370
rect 22652 8306 22708 8318
rect 22204 7422 22206 7474
rect 22258 7422 22260 7474
rect 22204 7252 22260 7422
rect 22764 7364 22820 7374
rect 22428 7252 22484 7262
rect 22204 7186 22260 7196
rect 22316 7250 22484 7252
rect 22316 7198 22430 7250
rect 22482 7198 22484 7250
rect 22316 7196 22484 7198
rect 21756 6692 21812 6748
rect 22092 6916 22148 6926
rect 21868 6692 21924 6702
rect 21756 6690 21924 6692
rect 21756 6638 21870 6690
rect 21922 6638 21924 6690
rect 21756 6636 21924 6638
rect 21532 6626 21588 6636
rect 21868 6626 21924 6636
rect 22092 6690 22148 6860
rect 22092 6638 22094 6690
rect 22146 6638 22148 6690
rect 22092 6626 22148 6638
rect 22316 6692 22372 7196
rect 22428 7186 22484 7196
rect 22652 7250 22708 7262
rect 22652 7198 22654 7250
rect 22706 7198 22708 7250
rect 22316 6626 22372 6636
rect 22428 6580 22484 6590
rect 22652 6580 22708 7198
rect 22428 6578 22708 6580
rect 22428 6526 22430 6578
rect 22482 6526 22708 6578
rect 22428 6524 22708 6526
rect 22092 6466 22148 6478
rect 22092 6414 22094 6466
rect 22146 6414 22148 6466
rect 22092 6132 22148 6414
rect 21532 6130 22148 6132
rect 21532 6078 22094 6130
rect 22146 6078 22148 6130
rect 21532 6076 22148 6078
rect 21532 5906 21588 6076
rect 22092 6066 22148 6076
rect 21532 5854 21534 5906
rect 21586 5854 21588 5906
rect 21532 5842 21588 5854
rect 22316 5906 22372 5918
rect 22316 5854 22318 5906
rect 22370 5854 22372 5906
rect 21756 5796 21812 5806
rect 21756 5702 21812 5740
rect 22204 5794 22260 5806
rect 22204 5742 22206 5794
rect 22258 5742 22260 5794
rect 22092 5348 22148 5358
rect 22204 5348 22260 5742
rect 22316 5796 22372 5854
rect 22316 5730 22372 5740
rect 22092 5346 22260 5348
rect 22092 5294 22094 5346
rect 22146 5294 22260 5346
rect 22092 5292 22260 5294
rect 22092 5282 22148 5292
rect 22204 5124 22260 5134
rect 22204 5030 22260 5068
rect 21420 4898 21476 4910
rect 21420 4846 21422 4898
rect 21474 4846 21476 4898
rect 21420 4340 21476 4846
rect 22428 4900 22484 6524
rect 22540 6020 22596 6030
rect 22540 5926 22596 5964
rect 22540 5460 22596 5470
rect 22540 5010 22596 5404
rect 22764 5236 22820 7308
rect 22876 6468 22932 8652
rect 22988 8484 23044 8876
rect 22988 8418 23044 8428
rect 23324 8820 23380 8830
rect 23100 8148 23156 8158
rect 22988 8034 23044 8046
rect 22988 7982 22990 8034
rect 23042 7982 23044 8034
rect 22988 6692 23044 7982
rect 23100 7698 23156 8092
rect 23324 8034 23380 8764
rect 23324 7982 23326 8034
rect 23378 7982 23380 8034
rect 23100 7646 23102 7698
rect 23154 7646 23156 7698
rect 23100 7634 23156 7646
rect 23212 7924 23268 7934
rect 22988 6636 23156 6692
rect 23100 6580 23156 6636
rect 23100 6514 23156 6524
rect 22988 6468 23044 6478
rect 22876 6466 23044 6468
rect 22876 6414 22990 6466
rect 23042 6414 23044 6466
rect 22876 6412 23044 6414
rect 22988 6402 23044 6412
rect 22988 6132 23044 6142
rect 22988 5684 23044 6076
rect 22988 5618 23044 5628
rect 22540 4958 22542 5010
rect 22594 4958 22596 5010
rect 22540 4946 22596 4958
rect 22652 5180 22820 5236
rect 22428 4834 22484 4844
rect 21420 3668 21476 4284
rect 21532 4228 21588 4238
rect 21532 4226 22148 4228
rect 21532 4174 21534 4226
rect 21586 4174 22148 4226
rect 21532 4172 22148 4174
rect 21532 4162 21588 4172
rect 22092 3778 22148 4172
rect 22428 3780 22484 3790
rect 22092 3726 22094 3778
rect 22146 3726 22148 3778
rect 22092 3714 22148 3726
rect 22204 3778 22484 3780
rect 22204 3726 22430 3778
rect 22482 3726 22484 3778
rect 22204 3724 22484 3726
rect 21420 3574 21476 3612
rect 21868 3668 21924 3678
rect 21868 3574 21924 3612
rect 22204 3666 22260 3724
rect 22428 3714 22484 3724
rect 22204 3614 22206 3666
rect 22258 3614 22260 3666
rect 22204 3602 22260 3614
rect 22652 3668 22708 5180
rect 23100 5122 23156 5134
rect 23100 5070 23102 5122
rect 23154 5070 23156 5122
rect 22764 5012 22820 5022
rect 22764 4918 22820 4956
rect 22876 4898 22932 4910
rect 22876 4846 22878 4898
rect 22930 4846 22932 4898
rect 22876 3778 22932 4846
rect 23100 4900 23156 5070
rect 23100 4228 23156 4844
rect 23100 4162 23156 4172
rect 22876 3726 22878 3778
rect 22930 3726 22932 3778
rect 22876 3714 22932 3726
rect 22764 3668 22820 3678
rect 22652 3666 22820 3668
rect 22652 3614 22766 3666
rect 22818 3614 22820 3666
rect 22652 3612 22820 3614
rect 22764 3602 22820 3612
rect 23212 3666 23268 7868
rect 23324 7364 23380 7982
rect 23436 7698 23492 8876
rect 23548 8036 23604 10108
rect 23660 8258 23716 11788
rect 23884 11506 23940 13580
rect 24108 12738 24164 12750
rect 24108 12686 24110 12738
rect 24162 12686 24164 12738
rect 24108 12292 24164 12686
rect 24108 12226 24164 12236
rect 24220 12068 24276 13692
rect 24220 12002 24276 12012
rect 24332 13300 24388 13310
rect 23996 11620 24052 11630
rect 24052 11564 24164 11620
rect 23996 11554 24052 11564
rect 23884 11454 23886 11506
rect 23938 11454 23940 11506
rect 23884 10836 23940 11454
rect 23884 10770 23940 10780
rect 23772 10724 23828 10734
rect 23772 10610 23828 10668
rect 23772 10558 23774 10610
rect 23826 10558 23828 10610
rect 23772 10546 23828 10558
rect 23996 10610 24052 10622
rect 23996 10558 23998 10610
rect 24050 10558 24052 10610
rect 23884 10498 23940 10510
rect 23884 10446 23886 10498
rect 23938 10446 23940 10498
rect 23772 9940 23828 9950
rect 23884 9940 23940 10446
rect 23996 10164 24052 10558
rect 23996 10098 24052 10108
rect 23772 9938 23940 9940
rect 23772 9886 23774 9938
rect 23826 9886 23940 9938
rect 23772 9884 23940 9886
rect 23772 9874 23828 9884
rect 23884 8930 23940 8942
rect 23884 8878 23886 8930
rect 23938 8878 23940 8930
rect 23884 8818 23940 8878
rect 23884 8766 23886 8818
rect 23938 8766 23940 8818
rect 23884 8754 23940 8766
rect 23660 8206 23662 8258
rect 23714 8206 23716 8258
rect 23660 8194 23716 8206
rect 23884 8260 23940 8270
rect 23772 8146 23828 8158
rect 23772 8094 23774 8146
rect 23826 8094 23828 8146
rect 23772 8036 23828 8094
rect 23548 7980 23828 8036
rect 23436 7646 23438 7698
rect 23490 7646 23492 7698
rect 23436 7634 23492 7646
rect 23884 7698 23940 8204
rect 23884 7646 23886 7698
rect 23938 7646 23940 7698
rect 23884 7634 23940 7646
rect 23324 7298 23380 7308
rect 24108 7140 24164 11564
rect 24332 10388 24388 13244
rect 24556 13188 24612 15092
rect 24668 13636 24724 13646
rect 24780 13636 24836 16380
rect 25228 16100 25284 16110
rect 25228 15986 25284 16044
rect 25228 15934 25230 15986
rect 25282 15934 25284 15986
rect 25228 15922 25284 15934
rect 24892 15876 24948 15886
rect 24892 14532 24948 15820
rect 25228 15316 25284 15326
rect 25340 15316 25396 18396
rect 25564 17780 25620 17790
rect 25676 17780 25732 21644
rect 25564 17778 25732 17780
rect 25564 17726 25566 17778
rect 25618 17726 25732 17778
rect 25564 17724 25732 17726
rect 25564 17714 25620 17724
rect 25788 17668 25844 24892
rect 25900 24882 25956 24892
rect 26012 23268 26068 23278
rect 26012 23174 26068 23212
rect 25900 23154 25956 23166
rect 25900 23102 25902 23154
rect 25954 23102 25956 23154
rect 25900 20692 25956 23102
rect 26012 21588 26068 21598
rect 26012 21494 26068 21532
rect 26124 20692 26180 20702
rect 25900 20690 26180 20692
rect 25900 20638 26126 20690
rect 26178 20638 26180 20690
rect 25900 20636 26180 20638
rect 26124 20468 26180 20636
rect 26124 20402 26180 20412
rect 26236 20242 26292 25452
rect 26572 25396 26628 26124
rect 26684 25508 26740 25518
rect 26684 25414 26740 25452
rect 26572 25330 26628 25340
rect 26908 25284 26964 25294
rect 27020 25284 27076 26236
rect 27244 26290 27300 26302
rect 27244 26238 27246 26290
rect 27298 26238 27300 26290
rect 27244 26180 27300 26238
rect 27244 26114 27300 26124
rect 26964 25228 27076 25284
rect 27244 25844 27300 25854
rect 26908 25218 26964 25228
rect 26796 23940 26852 23950
rect 26572 23938 26852 23940
rect 26572 23886 26798 23938
rect 26850 23886 26852 23938
rect 26572 23884 26852 23886
rect 26572 23268 26628 23884
rect 26796 23874 26852 23884
rect 27132 23938 27188 23950
rect 27132 23886 27134 23938
rect 27186 23886 27188 23938
rect 26572 23174 26628 23212
rect 27020 23714 27076 23726
rect 27020 23662 27022 23714
rect 27074 23662 27076 23714
rect 27020 22708 27076 23662
rect 27132 23154 27188 23886
rect 27132 23102 27134 23154
rect 27186 23102 27188 23154
rect 27132 22932 27188 23102
rect 27132 22866 27188 22876
rect 27132 22708 27188 22718
rect 27020 22652 27132 22708
rect 27132 22642 27188 22652
rect 26348 22370 26404 22382
rect 26348 22318 26350 22370
rect 26402 22318 26404 22370
rect 26348 21700 26404 22318
rect 26684 22146 26740 22158
rect 26684 22094 26686 22146
rect 26738 22094 26740 22146
rect 26684 22036 26740 22094
rect 27244 22036 27300 25788
rect 27356 25620 27412 26852
rect 27468 26852 27524 26862
rect 27468 26758 27524 26796
rect 27468 26404 27524 26414
rect 27468 26290 27524 26348
rect 27468 26238 27470 26290
rect 27522 26238 27524 26290
rect 27468 26226 27524 26238
rect 27580 26180 27636 26190
rect 27580 26086 27636 26124
rect 27692 25732 27748 28924
rect 28140 28868 28196 28878
rect 27804 28644 27860 28654
rect 28140 28644 28196 28812
rect 28476 28756 28532 28766
rect 28476 28662 28532 28700
rect 27804 28642 28196 28644
rect 27804 28590 27806 28642
rect 27858 28590 28142 28642
rect 28194 28590 28196 28642
rect 27804 28588 28196 28590
rect 27804 28084 27860 28588
rect 28140 28578 28196 28588
rect 28588 28532 28644 29372
rect 28700 29204 28756 30156
rect 29260 30100 29316 30110
rect 29148 29540 29204 29550
rect 29148 29446 29204 29484
rect 28812 29428 28868 29438
rect 28812 29334 28868 29372
rect 28700 29148 28868 29204
rect 28476 28476 28644 28532
rect 27804 28018 27860 28028
rect 28364 28420 28420 28430
rect 27804 27858 27860 27870
rect 28140 27860 28196 27870
rect 27804 27806 27806 27858
rect 27858 27806 27860 27858
rect 27804 27076 27860 27806
rect 27804 27010 27860 27020
rect 28028 27804 28140 27860
rect 28028 27186 28084 27804
rect 28140 27766 28196 27804
rect 28364 27412 28420 28364
rect 28364 27346 28420 27356
rect 28028 27134 28030 27186
rect 28082 27134 28084 27186
rect 28028 26180 28084 27134
rect 28252 27076 28308 27086
rect 28252 26982 28308 27020
rect 28028 26114 28084 26124
rect 27580 25620 27636 25658
rect 27356 25564 27580 25620
rect 27356 25396 27412 25564
rect 27580 25554 27636 25564
rect 27356 25330 27412 25340
rect 27580 25396 27636 25406
rect 26684 21980 27300 22036
rect 27356 25172 27412 25182
rect 27356 21810 27412 25116
rect 27580 23828 27636 25340
rect 27356 21758 27358 21810
rect 27410 21758 27412 21810
rect 27356 21746 27412 21758
rect 27468 23826 27636 23828
rect 27468 23774 27582 23826
rect 27634 23774 27636 23826
rect 27468 23772 27636 23774
rect 26684 21700 26740 21710
rect 26348 21698 26740 21700
rect 26348 21646 26686 21698
rect 26738 21646 26740 21698
rect 26348 21644 26740 21646
rect 26236 20190 26238 20242
rect 26290 20190 26292 20242
rect 26236 20178 26292 20190
rect 26460 20018 26516 21644
rect 26684 21364 26740 21644
rect 27468 21588 27524 23772
rect 27580 23762 27636 23772
rect 27692 23268 27748 25676
rect 27916 25394 27972 25406
rect 27916 25342 27918 25394
rect 27970 25342 27972 25394
rect 27916 24276 27972 25342
rect 28252 25284 28308 25294
rect 28252 25190 28308 25228
rect 27916 24220 28308 24276
rect 27916 23940 27972 23950
rect 27692 23212 27860 23268
rect 27580 22258 27636 22270
rect 27580 22206 27582 22258
rect 27634 22206 27636 22258
rect 27580 22148 27636 22206
rect 27580 22082 27636 22092
rect 26684 21298 26740 21308
rect 27356 21532 27524 21588
rect 27580 21586 27636 21598
rect 27580 21534 27582 21586
rect 27634 21534 27636 21586
rect 27020 20580 27076 20590
rect 27020 20486 27076 20524
rect 26460 19966 26462 20018
rect 26514 19966 26516 20018
rect 26460 19954 26516 19966
rect 26796 20020 26852 20030
rect 26796 19926 26852 19964
rect 27132 20020 27188 20030
rect 26908 19908 26964 19918
rect 26908 19906 27076 19908
rect 26908 19854 26910 19906
rect 26962 19854 27076 19906
rect 26908 19852 27076 19854
rect 26908 19842 26964 19852
rect 26684 19460 26740 19470
rect 26684 19346 26740 19404
rect 26684 19294 26686 19346
rect 26738 19294 26740 19346
rect 26684 19282 26740 19294
rect 27020 19348 27076 19852
rect 27020 19282 27076 19292
rect 26908 18900 26964 18910
rect 26012 18340 26068 18350
rect 26012 18246 26068 18284
rect 25676 17612 25844 17668
rect 25900 17668 25956 17678
rect 25228 15314 25396 15316
rect 25228 15262 25230 15314
rect 25282 15262 25396 15314
rect 25228 15260 25396 15262
rect 25564 16100 25620 16110
rect 25228 15204 25284 15260
rect 25228 15138 25284 15148
rect 24892 14438 24948 14476
rect 25452 14532 25508 14542
rect 25452 14438 25508 14476
rect 25116 14308 25172 14318
rect 25116 14214 25172 14252
rect 25116 13972 25172 13982
rect 25004 13748 25060 13758
rect 24668 13634 24948 13636
rect 24668 13582 24670 13634
rect 24722 13582 24948 13634
rect 24668 13580 24948 13582
rect 24668 13570 24724 13580
rect 24444 13132 24612 13188
rect 24444 11506 24500 13132
rect 24444 11454 24446 11506
rect 24498 11454 24500 11506
rect 24444 11442 24500 11454
rect 24556 12962 24612 12974
rect 24556 12910 24558 12962
rect 24610 12910 24612 12962
rect 24444 10498 24500 10510
rect 24444 10446 24446 10498
rect 24498 10446 24500 10498
rect 24444 10388 24500 10446
rect 24220 10332 24500 10388
rect 24220 7812 24276 10332
rect 24220 7746 24276 7756
rect 24332 9828 24388 9838
rect 24556 9828 24612 12910
rect 24668 12066 24724 12078
rect 24668 12014 24670 12066
rect 24722 12014 24724 12066
rect 24668 11844 24724 12014
rect 24668 11778 24724 11788
rect 24780 11508 24836 11518
rect 24780 11414 24836 11452
rect 24892 10500 24948 13580
rect 24892 10434 24948 10444
rect 24892 9828 24948 9838
rect 24388 9826 24892 9828
rect 24388 9774 24558 9826
rect 24610 9774 24892 9826
rect 24388 9772 24892 9774
rect 24220 7588 24276 7598
rect 24220 7494 24276 7532
rect 23884 7084 24164 7140
rect 23548 6690 23604 6702
rect 23548 6638 23550 6690
rect 23602 6638 23604 6690
rect 23324 6018 23380 6030
rect 23324 5966 23326 6018
rect 23378 5966 23380 6018
rect 23324 5460 23380 5966
rect 23324 5394 23380 5404
rect 23436 5796 23492 5806
rect 23436 5348 23492 5740
rect 23436 5254 23492 5292
rect 23212 3614 23214 3666
rect 23266 3614 23268 3666
rect 23212 3602 23268 3614
rect 23548 3556 23604 6638
rect 23772 6468 23828 6478
rect 23660 6466 23828 6468
rect 23660 6414 23774 6466
rect 23826 6414 23828 6466
rect 23660 6412 23828 6414
rect 23660 5012 23716 6412
rect 23772 6402 23828 6412
rect 23884 6130 23940 7084
rect 24220 6692 24276 6702
rect 24332 6692 24388 9772
rect 24556 9762 24612 9772
rect 24892 9734 24948 9772
rect 25004 9604 25060 13692
rect 25116 12180 25172 13916
rect 25564 13858 25620 16044
rect 25676 14084 25732 17612
rect 25900 17574 25956 17612
rect 26012 17554 26068 17566
rect 26012 17502 26014 17554
rect 26066 17502 26068 17554
rect 26012 17332 26068 17502
rect 26012 17266 26068 17276
rect 26348 17442 26404 17454
rect 26348 17390 26350 17442
rect 26402 17390 26404 17442
rect 26348 17108 26404 17390
rect 26348 17042 26404 17052
rect 26684 17442 26740 17454
rect 26684 17390 26686 17442
rect 26738 17390 26740 17442
rect 26236 16994 26292 17006
rect 26236 16942 26238 16994
rect 26290 16942 26292 16994
rect 25788 16884 25844 16894
rect 25788 16790 25844 16828
rect 26236 16212 26292 16942
rect 26572 16884 26628 16894
rect 26572 16790 26628 16828
rect 26684 16436 26740 17390
rect 26908 17108 26964 18844
rect 27132 17778 27188 19964
rect 27356 19458 27412 21532
rect 27580 20580 27636 21534
rect 27692 21588 27748 21598
rect 27692 20914 27748 21532
rect 27692 20862 27694 20914
rect 27746 20862 27748 20914
rect 27692 20850 27748 20862
rect 27580 20514 27636 20524
rect 27692 20356 27748 20366
rect 27468 20020 27524 20030
rect 27468 19926 27524 19964
rect 27692 20018 27748 20300
rect 27692 19966 27694 20018
rect 27746 19966 27748 20018
rect 27692 19954 27748 19966
rect 27356 19406 27358 19458
rect 27410 19406 27412 19458
rect 27356 19394 27412 19406
rect 27580 19236 27636 19246
rect 27580 19142 27636 19180
rect 27692 18900 27748 18910
rect 27804 18900 27860 23212
rect 27916 21700 27972 23884
rect 28140 23268 28196 23278
rect 27916 21634 27972 21644
rect 28028 22932 28084 22942
rect 28028 20802 28084 22876
rect 28140 22372 28196 23212
rect 28252 23154 28308 24220
rect 28476 23266 28532 28476
rect 28700 27970 28756 27982
rect 28700 27918 28702 27970
rect 28754 27918 28756 27970
rect 28700 27076 28756 27918
rect 28700 27010 28756 27020
rect 28588 26850 28644 26862
rect 28588 26798 28590 26850
rect 28642 26798 28644 26850
rect 28588 26516 28644 26798
rect 28588 26450 28644 26460
rect 28588 26290 28644 26302
rect 28588 26238 28590 26290
rect 28642 26238 28644 26290
rect 28588 25956 28644 26238
rect 28588 25890 28644 25900
rect 28588 25396 28644 25406
rect 28588 25302 28644 25340
rect 28812 24834 28868 29148
rect 29148 28530 29204 28542
rect 29148 28478 29150 28530
rect 29202 28478 29204 28530
rect 29148 28420 29204 28478
rect 29260 28532 29316 30044
rect 29372 29988 29428 29998
rect 29596 29988 29652 29998
rect 29372 29986 29540 29988
rect 29372 29934 29374 29986
rect 29426 29934 29540 29986
rect 29372 29932 29540 29934
rect 29372 29922 29428 29932
rect 29372 28866 29428 28878
rect 29372 28814 29374 28866
rect 29426 28814 29428 28866
rect 29372 28644 29428 28814
rect 29484 28868 29540 29932
rect 29596 29894 29652 29932
rect 29708 29764 29764 30156
rect 30268 30210 30436 30212
rect 30268 30158 30382 30210
rect 30434 30158 30436 30210
rect 30268 30156 30436 30158
rect 29932 30098 29988 30110
rect 29932 30046 29934 30098
rect 29986 30046 29988 30098
rect 29708 29314 29764 29708
rect 29708 29262 29710 29314
rect 29762 29262 29764 29314
rect 29708 29250 29764 29262
rect 29820 29986 29876 29998
rect 29820 29934 29822 29986
rect 29874 29934 29876 29986
rect 29484 28754 29540 28812
rect 29484 28702 29486 28754
rect 29538 28702 29540 28754
rect 29484 28690 29540 28702
rect 29372 28578 29428 28588
rect 29820 28644 29876 29934
rect 29932 28980 29988 30046
rect 30156 29540 30212 29550
rect 30156 29446 30212 29484
rect 29932 28914 29988 28924
rect 29820 28578 29876 28588
rect 29260 28466 29316 28476
rect 29148 28354 29204 28364
rect 28812 24782 28814 24834
rect 28866 24782 28868 24834
rect 28476 23214 28478 23266
rect 28530 23214 28532 23266
rect 28476 23202 28532 23214
rect 28588 24612 28644 24622
rect 28252 23102 28254 23154
rect 28306 23102 28308 23154
rect 28252 22708 28308 23102
rect 28252 22642 28308 22652
rect 28140 22278 28196 22316
rect 28476 20916 28532 20926
rect 28028 20750 28030 20802
rect 28082 20750 28084 20802
rect 27748 18844 27860 18900
rect 27916 20580 27972 20590
rect 27916 20132 27972 20524
rect 27916 19234 27972 20076
rect 28028 19794 28084 20750
rect 28028 19742 28030 19794
rect 28082 19742 28084 19794
rect 28028 19730 28084 19742
rect 28252 20804 28308 20814
rect 28140 19348 28196 19358
rect 28140 19254 28196 19292
rect 27916 19182 27918 19234
rect 27970 19182 27972 19234
rect 27692 18834 27748 18844
rect 27916 17892 27972 19182
rect 28140 18340 28196 18350
rect 28252 18340 28308 20748
rect 28476 20802 28532 20860
rect 28476 20750 28478 20802
rect 28530 20750 28532 20802
rect 28476 20738 28532 20750
rect 27132 17726 27134 17778
rect 27186 17726 27188 17778
rect 27132 17220 27188 17726
rect 27692 17836 27972 17892
rect 28028 18338 28308 18340
rect 28028 18286 28142 18338
rect 28194 18286 28308 18338
rect 28028 18284 28308 18286
rect 28364 20692 28420 20702
rect 27356 17554 27412 17566
rect 27356 17502 27358 17554
rect 27410 17502 27412 17554
rect 27356 17332 27412 17502
rect 27692 17554 27748 17836
rect 27692 17502 27694 17554
rect 27746 17502 27748 17554
rect 27692 17490 27748 17502
rect 28028 17666 28084 18284
rect 28140 18274 28196 18284
rect 28028 17614 28030 17666
rect 28082 17614 28084 17666
rect 28028 17332 28084 17614
rect 28364 17556 28420 20636
rect 28588 20244 28644 24556
rect 28476 20188 28644 20244
rect 28700 22148 28756 22158
rect 28476 18116 28532 20188
rect 28588 19906 28644 19918
rect 28588 19854 28590 19906
rect 28642 19854 28644 19906
rect 28588 18340 28644 19854
rect 28700 19348 28756 22092
rect 28700 19282 28756 19292
rect 28812 19236 28868 24782
rect 28924 28308 28980 28318
rect 28924 19906 28980 28252
rect 29708 27970 29764 27982
rect 29708 27918 29710 27970
rect 29762 27918 29764 27970
rect 29372 27860 29428 27870
rect 29372 27298 29428 27804
rect 29372 27246 29374 27298
rect 29426 27246 29428 27298
rect 29372 27234 29428 27246
rect 29148 27188 29204 27198
rect 29148 27094 29204 27132
rect 29708 27188 29764 27918
rect 29820 27860 29876 27870
rect 29820 27766 29876 27804
rect 29708 27122 29764 27132
rect 29484 27076 29540 27086
rect 29148 26404 29204 26414
rect 29148 25284 29204 26348
rect 29484 25730 29540 27020
rect 29708 26850 29764 26862
rect 29708 26798 29710 26850
rect 29762 26798 29764 26850
rect 29708 26292 29764 26798
rect 30268 26516 30324 30156
rect 30380 30146 30436 30156
rect 30940 30210 30996 30222
rect 30940 30158 30942 30210
rect 30994 30158 30996 30210
rect 30940 29764 30996 30158
rect 32060 30210 32116 30222
rect 32060 30158 32062 30210
rect 32114 30158 32116 30210
rect 30940 29698 30996 29708
rect 31052 30098 31108 30110
rect 31052 30046 31054 30098
rect 31106 30046 31108 30098
rect 30380 29540 30436 29550
rect 30380 28756 30436 29484
rect 31052 29540 31108 30046
rect 31948 30098 32004 30110
rect 31948 30046 31950 30098
rect 32002 30046 32004 30098
rect 31052 29474 31108 29484
rect 31500 29764 31556 29774
rect 30828 29428 30884 29438
rect 30828 28866 30884 29372
rect 31388 28980 31444 28990
rect 30828 28814 30830 28866
rect 30882 28814 30884 28866
rect 30828 28802 30884 28814
rect 31052 28868 31108 28878
rect 30380 27298 30436 28700
rect 31052 28642 31108 28812
rect 31052 28590 31054 28642
rect 31106 28590 31108 28642
rect 31052 27746 31108 28590
rect 31052 27694 31054 27746
rect 31106 27694 31108 27746
rect 31052 27682 31108 27694
rect 30380 27246 30382 27298
rect 30434 27246 30436 27298
rect 30380 27234 30436 27246
rect 30940 27186 30996 27198
rect 30940 27134 30942 27186
rect 30994 27134 30996 27186
rect 30604 27074 30660 27086
rect 30604 27022 30606 27074
rect 30658 27022 30660 27074
rect 30604 26964 30660 27022
rect 30604 26898 30660 26908
rect 29708 26226 29764 26236
rect 30156 26460 30324 26516
rect 30156 25844 30212 26460
rect 29932 25788 30212 25844
rect 30268 26290 30324 26302
rect 30268 26238 30270 26290
rect 30322 26238 30324 26290
rect 29484 25678 29486 25730
rect 29538 25678 29540 25730
rect 29484 25666 29540 25678
rect 29596 25732 29652 25742
rect 29596 25618 29652 25676
rect 29596 25566 29598 25618
rect 29650 25566 29652 25618
rect 29484 25508 29540 25518
rect 29484 25414 29540 25452
rect 29148 24052 29204 25228
rect 29148 24050 29540 24052
rect 29148 23998 29150 24050
rect 29202 23998 29540 24050
rect 29148 23996 29540 23998
rect 29148 23986 29204 23996
rect 29260 22370 29316 22382
rect 29260 22318 29262 22370
rect 29314 22318 29316 22370
rect 29036 21700 29092 21710
rect 29036 21606 29092 21644
rect 29260 21700 29316 22318
rect 29260 21140 29316 21644
rect 29484 21588 29540 23996
rect 29596 22594 29652 25566
rect 29932 24162 29988 25788
rect 30268 25732 30324 26238
rect 30156 25676 30324 25732
rect 30604 26290 30660 26302
rect 30604 26238 30606 26290
rect 30658 26238 30660 26290
rect 30604 25732 30660 26238
rect 30940 25956 30996 27134
rect 30940 25890 30996 25900
rect 31276 26852 31332 26862
rect 29932 24110 29934 24162
rect 29986 24110 29988 24162
rect 29932 24098 29988 24110
rect 30044 25620 30100 25630
rect 29932 23940 29988 23950
rect 29708 23716 29764 23726
rect 29708 23714 29876 23716
rect 29708 23662 29710 23714
rect 29762 23662 29876 23714
rect 29708 23660 29876 23662
rect 29708 23650 29764 23660
rect 29596 22542 29598 22594
rect 29650 22542 29652 22594
rect 29596 22530 29652 22542
rect 29708 22370 29764 22382
rect 29708 22318 29710 22370
rect 29762 22318 29764 22370
rect 29708 21924 29764 22318
rect 29708 21858 29764 21868
rect 29596 21588 29652 21598
rect 29484 21586 29652 21588
rect 29484 21534 29598 21586
rect 29650 21534 29652 21586
rect 29484 21532 29652 21534
rect 29596 21522 29652 21532
rect 29036 21084 29316 21140
rect 29036 20356 29092 21084
rect 29036 20290 29092 20300
rect 29148 20916 29204 20926
rect 28924 19854 28926 19906
rect 28978 19854 28980 19906
rect 28924 19842 28980 19854
rect 29148 19458 29204 20860
rect 29820 20916 29876 23660
rect 29932 22708 29988 23884
rect 30044 23266 30100 25564
rect 30044 23214 30046 23266
rect 30098 23214 30100 23266
rect 30044 23202 30100 23214
rect 30156 23828 30212 25676
rect 30604 25666 30660 25676
rect 31164 25618 31220 25630
rect 31164 25566 31166 25618
rect 31218 25566 31220 25618
rect 30492 25506 30548 25518
rect 30716 25508 30772 25518
rect 30492 25454 30494 25506
rect 30546 25454 30548 25506
rect 30492 25060 30548 25454
rect 30492 24994 30548 25004
rect 30604 25506 30772 25508
rect 30604 25454 30718 25506
rect 30770 25454 30772 25506
rect 30604 25452 30772 25454
rect 30156 23044 30212 23772
rect 30268 24724 30324 24734
rect 30268 23938 30324 24668
rect 30604 24612 30660 25452
rect 30716 25442 30772 25452
rect 31052 25284 31108 25294
rect 31052 25190 31108 25228
rect 31164 24834 31220 25566
rect 31276 25396 31332 26796
rect 31388 26402 31444 28924
rect 31500 28642 31556 29708
rect 31612 29538 31668 29550
rect 31612 29486 31614 29538
rect 31666 29486 31668 29538
rect 31612 29428 31668 29486
rect 31612 29362 31668 29372
rect 31836 29316 31892 29326
rect 31836 29222 31892 29260
rect 31948 28868 32004 30046
rect 32060 29988 32116 30158
rect 32060 29922 32116 29932
rect 31948 28802 32004 28812
rect 31612 28756 31668 28766
rect 31612 28662 31668 28700
rect 31500 28590 31502 28642
rect 31554 28590 31556 28642
rect 31500 28578 31556 28590
rect 32172 28420 32228 33964
rect 33180 34018 33236 34030
rect 33180 33966 33182 34018
rect 33234 33966 33236 34018
rect 32508 33572 32564 33582
rect 33180 33572 33236 33966
rect 33516 33908 33572 33918
rect 32508 32788 32564 33516
rect 32732 33516 33236 33572
rect 33404 33852 33516 33908
rect 32732 33458 32788 33516
rect 32732 33406 32734 33458
rect 32786 33406 32788 33458
rect 32732 33394 32788 33406
rect 32508 32694 32564 32732
rect 33180 32450 33236 32462
rect 33180 32398 33182 32450
rect 33234 32398 33236 32450
rect 32620 31892 32676 31902
rect 32620 31798 32676 31836
rect 33068 31780 33124 31790
rect 33068 31666 33124 31724
rect 33068 31614 33070 31666
rect 33122 31614 33124 31666
rect 33068 31602 33124 31614
rect 33180 31666 33236 32398
rect 33180 31614 33182 31666
rect 33234 31614 33236 31666
rect 32844 31556 32900 31566
rect 32620 31554 32900 31556
rect 32620 31502 32846 31554
rect 32898 31502 32900 31554
rect 32620 31500 32900 31502
rect 32620 30994 32676 31500
rect 32844 31490 32900 31500
rect 33180 31444 33236 31614
rect 33180 31378 33236 31388
rect 33068 31108 33124 31118
rect 33068 31014 33124 31052
rect 33292 31106 33348 31118
rect 33292 31054 33294 31106
rect 33346 31054 33348 31106
rect 32620 30942 32622 30994
rect 32674 30942 32676 30994
rect 32620 30930 32676 30942
rect 33180 30996 33236 31006
rect 33180 30902 33236 30940
rect 33292 30772 33348 31054
rect 33404 31108 33460 33852
rect 33516 33842 33572 33852
rect 33740 33012 33796 37436
rect 33852 35028 33908 38556
rect 33964 37154 34020 40124
rect 35532 40180 35588 40190
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35084 39732 35140 39742
rect 35084 39638 35140 39676
rect 34412 39620 34468 39630
rect 34412 39526 34468 39564
rect 35196 39620 35252 39630
rect 35532 39620 35588 40124
rect 36316 39842 36372 40348
rect 36316 39790 36318 39842
rect 36370 39790 36372 39842
rect 36316 39778 36372 39790
rect 35252 39618 35588 39620
rect 35252 39566 35534 39618
rect 35586 39566 35588 39618
rect 35252 39564 35588 39566
rect 34076 39396 34132 39406
rect 34076 38946 34132 39340
rect 35196 39058 35252 39564
rect 35532 39554 35588 39564
rect 35980 39732 36036 39742
rect 35196 39006 35198 39058
rect 35250 39006 35252 39058
rect 35196 38994 35252 39006
rect 34076 38894 34078 38946
rect 34130 38894 34132 38946
rect 34076 38882 34132 38894
rect 35644 38948 35700 38958
rect 34748 38834 34804 38846
rect 34748 38782 34750 38834
rect 34802 38782 34804 38834
rect 34748 38668 34804 38782
rect 34972 38834 35028 38846
rect 34972 38782 34974 38834
rect 35026 38782 35028 38834
rect 34300 38612 34804 38668
rect 34860 38722 34916 38734
rect 34860 38670 34862 38722
rect 34914 38670 34916 38722
rect 34188 38052 34244 38062
rect 33964 37102 33966 37154
rect 34018 37102 34020 37154
rect 33964 36036 34020 37102
rect 33964 35970 34020 35980
rect 34076 37996 34188 38052
rect 34076 35308 34132 37996
rect 34188 37986 34244 37996
rect 34300 37380 34356 38612
rect 34860 38388 34916 38670
rect 34972 38668 35028 38782
rect 35644 38724 35700 38892
rect 35756 38724 35812 38734
rect 35644 38722 35812 38724
rect 35644 38670 35758 38722
rect 35810 38670 35812 38722
rect 35644 38668 35812 38670
rect 34972 38612 35140 38668
rect 34860 38332 35028 38388
rect 34748 38164 34804 38174
rect 34412 37940 34468 37950
rect 34412 37490 34468 37884
rect 34412 37438 34414 37490
rect 34466 37438 34468 37490
rect 34412 37426 34468 37438
rect 34300 37286 34356 37324
rect 34636 37268 34692 37278
rect 34748 37268 34804 38108
rect 34860 38162 34916 38174
rect 34860 38110 34862 38162
rect 34914 38110 34916 38162
rect 34860 37940 34916 38110
rect 34860 37874 34916 37884
rect 34860 37380 34916 37390
rect 34972 37380 35028 38332
rect 35084 38164 35140 38612
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35084 38098 35140 38108
rect 35644 37940 35700 38668
rect 35756 38658 35812 38668
rect 35868 38164 35924 38174
rect 35868 38070 35924 38108
rect 35420 37884 35700 37940
rect 35308 37828 35364 37838
rect 34860 37378 35028 37380
rect 34860 37326 34862 37378
rect 34914 37326 35028 37378
rect 34860 37324 35028 37326
rect 35084 37772 35308 37828
rect 34860 37314 34916 37324
rect 34636 37266 34804 37268
rect 34636 37214 34638 37266
rect 34690 37214 34804 37266
rect 34636 37212 34804 37214
rect 34636 37202 34692 37212
rect 34188 36482 34244 36494
rect 34188 36430 34190 36482
rect 34242 36430 34244 36482
rect 34188 35812 34244 36430
rect 34748 36484 34804 37212
rect 35084 36594 35140 37772
rect 35308 37734 35364 37772
rect 35196 37380 35252 37390
rect 35196 37286 35252 37324
rect 35420 37266 35476 37884
rect 35980 37492 36036 39676
rect 36428 39620 36484 39630
rect 36540 39620 36596 41244
rect 36876 41076 36932 41806
rect 36876 41010 36932 41020
rect 36988 40740 37044 42030
rect 37324 41972 37380 41982
rect 36988 40674 37044 40684
rect 37212 41970 37380 41972
rect 37212 41918 37326 41970
rect 37378 41918 37380 41970
rect 37212 41916 37380 41918
rect 37212 41860 37268 41916
rect 37324 41906 37380 41916
rect 37100 40628 37156 40638
rect 37100 40534 37156 40572
rect 36876 40514 36932 40526
rect 36876 40462 36878 40514
rect 36930 40462 36932 40514
rect 36764 40404 36820 40414
rect 36764 40310 36820 40348
rect 36876 39844 36932 40462
rect 37212 40180 37268 41804
rect 37436 41636 37492 41646
rect 37436 41188 37492 41580
rect 37436 41094 37492 41132
rect 37548 41186 37604 43036
rect 37660 42980 37716 42990
rect 37660 42082 37716 42924
rect 37660 42030 37662 42082
rect 37714 42030 37716 42082
rect 37660 42018 37716 42030
rect 37772 41970 37828 44940
rect 38780 44772 38836 45836
rect 38892 45826 38948 45836
rect 39228 45778 39284 45790
rect 39228 45726 39230 45778
rect 39282 45726 39284 45778
rect 38220 44324 38276 44334
rect 38108 44212 38164 44222
rect 37996 43876 38052 43886
rect 37772 41918 37774 41970
rect 37826 41918 37828 41970
rect 37772 41906 37828 41918
rect 37884 43428 37940 43438
rect 37884 41524 37940 43372
rect 37996 42082 38052 43820
rect 38108 43764 38164 44156
rect 38108 43538 38164 43708
rect 38108 43486 38110 43538
rect 38162 43486 38164 43538
rect 38108 43474 38164 43486
rect 37996 42030 37998 42082
rect 38050 42030 38052 42082
rect 37996 42018 38052 42030
rect 38108 42754 38164 42766
rect 38108 42702 38110 42754
rect 38162 42702 38164 42754
rect 38108 41748 38164 42702
rect 38220 42082 38276 44268
rect 38332 44212 38388 44222
rect 38332 43876 38388 44156
rect 38332 43810 38388 43820
rect 38332 43652 38388 43662
rect 38332 43558 38388 43596
rect 38780 43650 38836 44716
rect 39116 45666 39172 45678
rect 39116 45614 39118 45666
rect 39170 45614 39172 45666
rect 39116 44548 39172 45614
rect 39228 44884 39284 45726
rect 39228 44818 39284 44828
rect 39340 44994 39396 45006
rect 39340 44942 39342 44994
rect 39394 44942 39396 44994
rect 39340 44772 39396 44942
rect 39564 44884 39620 46284
rect 40348 46116 40404 46126
rect 40348 46002 40404 46060
rect 41244 46116 41300 49200
rect 42812 46788 42868 49200
rect 42812 46732 43092 46788
rect 41244 46050 41300 46060
rect 40348 45950 40350 46002
rect 40402 45950 40404 46002
rect 40348 45938 40404 45950
rect 42364 45890 42420 45902
rect 42364 45838 42366 45890
rect 42418 45838 42420 45890
rect 39676 45332 39732 45342
rect 39676 45330 40180 45332
rect 39676 45278 39678 45330
rect 39730 45278 40180 45330
rect 39676 45276 40180 45278
rect 39676 45266 39732 45276
rect 39900 45106 39956 45118
rect 39900 45054 39902 45106
rect 39954 45054 39956 45106
rect 39788 44994 39844 45006
rect 39788 44942 39790 44994
rect 39842 44942 39844 44994
rect 39564 44828 39732 44884
rect 39340 44706 39396 44716
rect 39116 44492 39620 44548
rect 39116 44324 39172 44334
rect 38780 43598 38782 43650
rect 38834 43598 38836 43650
rect 38780 43586 38836 43598
rect 38892 44322 39172 44324
rect 38892 44270 39118 44322
rect 39170 44270 39172 44322
rect 38892 44268 39172 44270
rect 38556 43538 38612 43550
rect 38556 43486 38558 43538
rect 38610 43486 38612 43538
rect 38444 43426 38500 43438
rect 38444 43374 38446 43426
rect 38498 43374 38500 43426
rect 38220 42030 38222 42082
rect 38274 42030 38276 42082
rect 38220 42018 38276 42030
rect 38332 42754 38388 42766
rect 38332 42702 38334 42754
rect 38386 42702 38388 42754
rect 38332 42084 38388 42702
rect 38444 42420 38500 43374
rect 38556 43428 38612 43486
rect 38556 43362 38612 43372
rect 38892 42868 38948 44268
rect 39116 44258 39172 44268
rect 39340 44100 39396 44110
rect 39228 43652 39284 43662
rect 39116 43540 39172 43550
rect 39004 43538 39172 43540
rect 39004 43486 39118 43538
rect 39170 43486 39172 43538
rect 39004 43484 39172 43486
rect 39004 43092 39060 43484
rect 39116 43474 39172 43484
rect 39004 43026 39060 43036
rect 39116 43314 39172 43326
rect 39116 43262 39118 43314
rect 39170 43262 39172 43314
rect 38892 42802 38948 42812
rect 38556 42644 38612 42654
rect 39004 42644 39060 42654
rect 38556 42642 39060 42644
rect 38556 42590 38558 42642
rect 38610 42590 39006 42642
rect 39058 42590 39060 42642
rect 38556 42588 39060 42590
rect 38556 42578 38612 42588
rect 39004 42578 39060 42588
rect 38444 42364 38836 42420
rect 38332 42018 38388 42028
rect 38668 42084 38724 42094
rect 38668 41748 38724 42028
rect 38780 41970 38836 42364
rect 38892 42084 38948 42094
rect 38948 42028 39060 42084
rect 38892 41990 38948 42028
rect 38780 41918 38782 41970
rect 38834 41918 38836 41970
rect 38780 41906 38836 41918
rect 38108 41692 38500 41748
rect 38668 41692 38836 41748
rect 37884 41458 37940 41468
rect 37660 41300 37716 41310
rect 38332 41300 38388 41310
rect 37660 41298 38388 41300
rect 37660 41246 37662 41298
rect 37714 41246 38334 41298
rect 38386 41246 38388 41298
rect 37660 41244 38388 41246
rect 37660 41234 37716 41244
rect 37548 41134 37550 41186
rect 37602 41134 37604 41186
rect 37548 40964 37604 41134
rect 37996 41074 38052 41086
rect 37996 41022 37998 41074
rect 38050 41022 38052 41074
rect 37548 40898 37604 40908
rect 37772 40962 37828 40974
rect 37772 40910 37774 40962
rect 37826 40910 37828 40962
rect 37772 40628 37828 40910
rect 37772 40562 37828 40572
rect 37996 40516 38052 41022
rect 37212 40114 37268 40124
rect 37324 40402 37380 40414
rect 37324 40350 37326 40402
rect 37378 40350 37380 40402
rect 36876 39778 36932 39788
rect 36988 39620 37044 39630
rect 37212 39620 37268 39630
rect 36428 39618 36596 39620
rect 36428 39566 36430 39618
rect 36482 39566 36596 39618
rect 36428 39564 36596 39566
rect 36652 39618 37044 39620
rect 36652 39566 36990 39618
rect 37042 39566 37044 39618
rect 36652 39564 37044 39566
rect 36428 39554 36484 39564
rect 36540 38836 36596 38846
rect 36652 38836 36708 39564
rect 36988 39554 37044 39564
rect 37100 39618 37268 39620
rect 37100 39566 37214 39618
rect 37266 39566 37268 39618
rect 37100 39564 37268 39566
rect 36764 39060 36820 39070
rect 37100 39060 37156 39564
rect 37212 39554 37268 39564
rect 37324 39396 37380 40350
rect 37772 40404 37828 40414
rect 37772 40290 37828 40348
rect 37772 40238 37774 40290
rect 37826 40238 37828 40290
rect 37772 39956 37828 40238
rect 37772 39890 37828 39900
rect 37324 39330 37380 39340
rect 37436 39844 37492 39854
rect 37436 39618 37492 39788
rect 37548 39732 37604 39742
rect 37996 39732 38052 40460
rect 38108 40740 38164 40750
rect 38108 40404 38164 40684
rect 38332 40626 38388 41244
rect 38444 41298 38500 41692
rect 38444 41246 38446 41298
rect 38498 41246 38500 41298
rect 38444 41234 38500 41246
rect 38668 41412 38724 41422
rect 38668 41188 38724 41356
rect 38332 40574 38334 40626
rect 38386 40574 38388 40626
rect 38332 40562 38388 40574
rect 38556 41186 38724 41188
rect 38556 41134 38670 41186
rect 38722 41134 38724 41186
rect 38556 41132 38724 41134
rect 38556 40626 38612 41132
rect 38668 41094 38724 41132
rect 38556 40574 38558 40626
rect 38610 40574 38612 40626
rect 38556 40562 38612 40574
rect 38780 40626 38836 41692
rect 39004 41524 39060 42028
rect 38780 40574 38782 40626
rect 38834 40574 38836 40626
rect 38780 40562 38836 40574
rect 38892 41468 39060 41524
rect 38108 40338 38164 40348
rect 38444 40404 38500 40414
rect 38892 40404 38948 41468
rect 39116 41412 39172 43262
rect 39228 42756 39284 43596
rect 39340 42978 39396 44044
rect 39340 42926 39342 42978
rect 39394 42926 39396 42978
rect 39340 42914 39396 42926
rect 39452 43314 39508 43326
rect 39452 43262 39454 43314
rect 39506 43262 39508 43314
rect 39228 42700 39396 42756
rect 39228 42532 39284 42542
rect 39228 42438 39284 42476
rect 39116 41346 39172 41356
rect 38444 40402 38948 40404
rect 38444 40350 38446 40402
rect 38498 40350 38948 40402
rect 38444 40348 38948 40350
rect 39004 41188 39060 41198
rect 38444 40338 38500 40348
rect 37548 39730 38052 39732
rect 37548 39678 37550 39730
rect 37602 39678 38052 39730
rect 37548 39676 38052 39678
rect 38108 39956 38164 39966
rect 37548 39666 37604 39676
rect 37436 39566 37438 39618
rect 37490 39566 37492 39618
rect 36764 39058 37156 39060
rect 36764 39006 36766 39058
rect 36818 39006 37156 39058
rect 36764 39004 37156 39006
rect 36764 38994 36820 39004
rect 36540 38834 36708 38836
rect 36540 38782 36542 38834
rect 36594 38782 36708 38834
rect 36540 38780 36708 38782
rect 36092 38722 36148 38734
rect 36092 38670 36094 38722
rect 36146 38670 36148 38722
rect 36092 38276 36148 38670
rect 36540 38668 36596 38780
rect 36092 38210 36148 38220
rect 36428 38612 36596 38668
rect 36876 38724 36932 38762
rect 36876 38658 36932 38668
rect 35420 37214 35422 37266
rect 35474 37214 35476 37266
rect 35420 37202 35476 37214
rect 35532 37436 35980 37492
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35084 36542 35086 36594
rect 35138 36542 35140 36594
rect 35084 36530 35140 36542
rect 34748 36418 34804 36428
rect 34300 36372 34356 36382
rect 34636 36372 34692 36382
rect 34300 36370 34692 36372
rect 34300 36318 34302 36370
rect 34354 36318 34638 36370
rect 34690 36318 34692 36370
rect 34300 36316 34692 36318
rect 34300 36306 34356 36316
rect 34636 36306 34692 36316
rect 35084 36372 35140 36382
rect 34188 35700 34244 35756
rect 34972 35922 35028 35934
rect 34972 35870 34974 35922
rect 35026 35870 35028 35922
rect 34636 35700 34692 35710
rect 34188 35698 34692 35700
rect 34188 35646 34638 35698
rect 34690 35646 34692 35698
rect 34188 35644 34692 35646
rect 34636 35634 34692 35644
rect 34076 35242 34132 35252
rect 33852 34962 33908 34972
rect 34188 35028 34244 35038
rect 33852 34690 33908 34702
rect 33852 34638 33854 34690
rect 33906 34638 33908 34690
rect 33852 34132 33908 34638
rect 34188 34468 34244 34972
rect 34972 35028 35028 35870
rect 34300 34916 34356 34926
rect 34300 34822 34356 34860
rect 34412 34804 34468 34814
rect 34412 34802 34916 34804
rect 34412 34750 34414 34802
rect 34466 34750 34916 34802
rect 34412 34748 34916 34750
rect 34412 34738 34468 34748
rect 34188 34412 34580 34468
rect 34188 34132 34244 34142
rect 33852 34130 34244 34132
rect 33852 34078 34190 34130
rect 34242 34078 34244 34130
rect 33852 34076 34244 34078
rect 33852 33012 33908 33022
rect 33740 32956 33852 33012
rect 33852 32946 33908 32956
rect 33516 32674 33572 32686
rect 33516 32622 33518 32674
rect 33570 32622 33572 32674
rect 33516 31890 33572 32622
rect 33516 31838 33518 31890
rect 33570 31838 33572 31890
rect 33516 31780 33572 31838
rect 34188 32452 34244 34076
rect 33572 31724 33908 31780
rect 33516 31686 33572 31724
rect 33740 31444 33796 31454
rect 33404 31052 33572 31108
rect 33292 30706 33348 30716
rect 32732 30212 32788 30222
rect 33292 30212 33348 30222
rect 32620 30210 33348 30212
rect 32620 30158 32734 30210
rect 32786 30158 33294 30210
rect 33346 30158 33348 30210
rect 32620 30156 33348 30158
rect 33516 30212 33572 31052
rect 33740 30994 33796 31388
rect 33852 31220 33908 31724
rect 33964 31220 34020 31230
rect 33852 31218 34020 31220
rect 33852 31166 33966 31218
rect 34018 31166 34020 31218
rect 33852 31164 34020 31166
rect 33964 31154 34020 31164
rect 33740 30942 33742 30994
rect 33794 30942 33796 30994
rect 33740 30930 33796 30942
rect 33852 30884 33908 30894
rect 33852 30790 33908 30828
rect 34188 30212 34244 32396
rect 34524 31218 34580 34412
rect 34860 33458 34916 34748
rect 34972 34802 35028 34972
rect 34972 34750 34974 34802
rect 35026 34750 35028 34802
rect 34972 34738 35028 34750
rect 35084 34692 35140 36316
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35308 35140 35364 35150
rect 35196 34916 35252 34926
rect 35196 34822 35252 34860
rect 35308 34914 35364 35084
rect 35308 34862 35310 34914
rect 35362 34862 35364 34914
rect 35308 34850 35364 34862
rect 35252 34692 35308 34702
rect 35084 34636 35252 34692
rect 35252 34626 35308 34636
rect 35420 34690 35476 34702
rect 35420 34638 35422 34690
rect 35474 34638 35476 34690
rect 35420 34580 35476 34638
rect 35420 34514 35476 34524
rect 35532 34018 35588 37436
rect 35980 37398 36036 37436
rect 36092 37940 36148 37950
rect 35868 37268 35924 37278
rect 36092 37268 36148 37884
rect 36204 37938 36260 37950
rect 36204 37886 36206 37938
rect 36258 37886 36260 37938
rect 36204 37828 36260 37886
rect 36204 37762 36260 37772
rect 36316 37826 36372 37838
rect 36316 37774 36318 37826
rect 36370 37774 36372 37826
rect 35868 37266 36148 37268
rect 35868 37214 35870 37266
rect 35922 37214 36148 37266
rect 35868 37212 36148 37214
rect 36204 37268 36260 37278
rect 35868 37202 35924 37212
rect 35644 36820 35700 36830
rect 35644 35924 35700 36764
rect 36204 36482 36260 37212
rect 36316 36820 36372 37774
rect 36316 36754 36372 36764
rect 36316 36596 36372 36606
rect 36428 36596 36484 38612
rect 36652 38276 36708 38286
rect 36316 36594 36484 36596
rect 36316 36542 36318 36594
rect 36370 36542 36484 36594
rect 36316 36540 36484 36542
rect 36540 37826 36596 37838
rect 36540 37774 36542 37826
rect 36594 37774 36596 37826
rect 36316 36530 36372 36540
rect 36204 36430 36206 36482
rect 36258 36430 36260 36482
rect 36204 36418 36260 36430
rect 35756 36372 35812 36382
rect 35756 36278 35812 36316
rect 35980 36258 36036 36270
rect 35980 36206 35982 36258
rect 36034 36206 36036 36258
rect 35980 36148 36036 36206
rect 35980 36082 36036 36092
rect 36316 36258 36372 36270
rect 36316 36206 36318 36258
rect 36370 36206 36372 36258
rect 35644 35586 35700 35868
rect 35644 35534 35646 35586
rect 35698 35534 35700 35586
rect 35644 35522 35700 35534
rect 36316 35924 36372 36206
rect 36540 36148 36596 37774
rect 36540 36082 36596 36092
rect 36652 37604 36708 38220
rect 37100 38162 37156 39004
rect 37212 38948 37268 38958
rect 37436 38948 37492 39566
rect 37660 39396 37716 39406
rect 37660 39302 37716 39340
rect 37884 39060 37940 39070
rect 37548 38948 37604 38958
rect 37436 38946 37604 38948
rect 37436 38894 37550 38946
rect 37602 38894 37604 38946
rect 37436 38892 37604 38894
rect 37212 38724 37268 38892
rect 37548 38882 37604 38892
rect 37212 38658 37268 38668
rect 37100 38110 37102 38162
rect 37154 38110 37156 38162
rect 37100 38098 37156 38110
rect 36988 37938 37044 37950
rect 36988 37886 36990 37938
rect 37042 37886 37044 37938
rect 36988 37604 37044 37886
rect 37772 37940 37828 37950
rect 37772 37846 37828 37884
rect 36652 37548 37044 37604
rect 37212 37828 37268 37838
rect 37660 37828 37716 37838
rect 37212 37826 37716 37828
rect 37212 37774 37214 37826
rect 37266 37774 37662 37826
rect 37714 37774 37716 37826
rect 37212 37772 37716 37774
rect 36652 35924 36708 37548
rect 36988 37380 37044 37390
rect 36988 37286 37044 37324
rect 36764 37268 36820 37278
rect 36764 37266 36932 37268
rect 36764 37214 36766 37266
rect 36818 37214 36932 37266
rect 36764 37212 36932 37214
rect 36764 37202 36820 37212
rect 36316 35868 36708 35924
rect 36876 35924 36932 37212
rect 37100 37266 37156 37278
rect 37100 37214 37102 37266
rect 37154 37214 37156 37266
rect 37100 36708 37156 37214
rect 37212 37268 37268 37772
rect 37660 37762 37716 37772
rect 37212 37202 37268 37212
rect 37436 37492 37492 37502
rect 37436 37266 37492 37436
rect 37436 37214 37438 37266
rect 37490 37214 37492 37266
rect 37436 37202 37492 37214
rect 37100 36642 37156 36652
rect 36988 36372 37044 36382
rect 36988 36278 37044 36316
rect 37884 36372 37940 39004
rect 38108 38834 38164 39900
rect 38220 39844 38276 39854
rect 38220 39730 38276 39788
rect 38220 39678 38222 39730
rect 38274 39678 38276 39730
rect 38220 39666 38276 39678
rect 38108 38782 38110 38834
rect 38162 38782 38164 38834
rect 38108 38770 38164 38782
rect 38780 38836 38836 38846
rect 38780 38742 38836 38780
rect 39004 38724 39060 41132
rect 39116 41076 39172 41086
rect 39340 41076 39396 42700
rect 39452 41636 39508 43262
rect 39564 41972 39620 44492
rect 39676 43428 39732 44828
rect 39788 44324 39844 44942
rect 39788 44258 39844 44268
rect 39900 44212 39956 45054
rect 39900 44118 39956 44156
rect 40012 44884 40068 44894
rect 40012 44322 40068 44828
rect 40012 44270 40014 44322
rect 40066 44270 40068 44322
rect 40012 43652 40068 44270
rect 39676 43362 39732 43372
rect 39900 43596 40068 43652
rect 39900 42980 39956 43596
rect 40012 43426 40068 43438
rect 40012 43374 40014 43426
rect 40066 43374 40068 43426
rect 40012 43204 40068 43374
rect 40012 43138 40068 43148
rect 40124 42980 40180 45276
rect 40236 45108 40292 45118
rect 41020 45108 41076 45118
rect 40236 45106 40516 45108
rect 40236 45054 40238 45106
rect 40290 45054 40516 45106
rect 40236 45052 40516 45054
rect 40236 45042 40292 45052
rect 40348 44772 40404 44782
rect 40348 44322 40404 44716
rect 40348 44270 40350 44322
rect 40402 44270 40404 44322
rect 40348 44258 40404 44270
rect 40236 43540 40292 43550
rect 40236 43426 40292 43484
rect 40236 43374 40238 43426
rect 40290 43374 40292 43426
rect 40236 43362 40292 43374
rect 39900 42924 40068 42980
rect 39676 42868 39732 42878
rect 39676 42866 39956 42868
rect 39676 42814 39678 42866
rect 39730 42814 39956 42866
rect 39676 42812 39956 42814
rect 39676 42802 39732 42812
rect 39788 42194 39844 42206
rect 39788 42142 39790 42194
rect 39842 42142 39844 42194
rect 39788 42084 39844 42142
rect 39788 42018 39844 42028
rect 39676 41972 39732 41982
rect 39564 41970 39732 41972
rect 39564 41918 39678 41970
rect 39730 41918 39732 41970
rect 39564 41916 39732 41918
rect 39676 41906 39732 41916
rect 39900 41972 39956 42812
rect 39452 41570 39508 41580
rect 39676 41188 39732 41198
rect 39676 41094 39732 41132
rect 39900 41186 39956 41916
rect 39900 41134 39902 41186
rect 39954 41134 39956 41186
rect 39900 41122 39956 41134
rect 39116 41074 39396 41076
rect 39116 41022 39118 41074
rect 39170 41022 39396 41074
rect 39116 41020 39396 41022
rect 39116 41010 39172 41020
rect 40012 40964 40068 42924
rect 40124 42914 40180 42924
rect 40236 41860 40292 41870
rect 39788 40908 40012 40964
rect 39228 40852 39284 40862
rect 39228 40626 39284 40796
rect 39228 40574 39230 40626
rect 39282 40574 39284 40626
rect 39228 40562 39284 40574
rect 39788 40514 39844 40908
rect 40012 40870 40068 40908
rect 40124 41858 40292 41860
rect 40124 41806 40238 41858
rect 40290 41806 40292 41858
rect 40124 41804 40292 41806
rect 39788 40462 39790 40514
rect 39842 40462 39844 40514
rect 39788 40450 39844 40462
rect 40012 40404 40068 40414
rect 40012 40310 40068 40348
rect 40012 40180 40068 40190
rect 40124 40180 40180 41804
rect 40236 41794 40292 41804
rect 40460 41860 40516 45052
rect 41020 45106 41412 45108
rect 41020 45054 41022 45106
rect 41074 45054 41412 45106
rect 41020 45052 41412 45054
rect 41020 45042 41076 45052
rect 41356 44322 41412 45052
rect 41692 44996 41748 45006
rect 41692 44994 41972 44996
rect 41692 44942 41694 44994
rect 41746 44942 41972 44994
rect 41692 44940 41972 44942
rect 41692 44930 41748 44940
rect 41356 44270 41358 44322
rect 41410 44270 41412 44322
rect 41132 43428 41188 43438
rect 41132 43334 41188 43372
rect 41356 42868 41412 44270
rect 41020 42812 41356 42868
rect 40460 41794 40516 41804
rect 40572 42644 40628 42654
rect 40348 41748 40404 41758
rect 40348 41654 40404 41692
rect 40236 40628 40292 40638
rect 40236 40534 40292 40572
rect 40348 40516 40404 40526
rect 40348 40422 40404 40460
rect 40236 40180 40292 40190
rect 40124 40124 40236 40180
rect 40012 39060 40068 40124
rect 40236 40114 40292 40124
rect 40348 39508 40404 39518
rect 40012 38966 40068 39004
rect 40124 39506 40404 39508
rect 40124 39454 40350 39506
rect 40402 39454 40404 39506
rect 40124 39452 40404 39454
rect 39004 38658 39060 38668
rect 39452 38724 39508 38734
rect 39788 38724 39844 38734
rect 39452 38722 39844 38724
rect 39452 38670 39454 38722
rect 39506 38670 39790 38722
rect 39842 38670 39844 38722
rect 39452 38668 39844 38670
rect 39452 38658 39508 38668
rect 39788 38658 39844 38668
rect 40124 38722 40180 39452
rect 40348 39442 40404 39452
rect 40124 38670 40126 38722
rect 40178 38670 40180 38722
rect 40124 38658 40180 38670
rect 40348 39060 40404 39070
rect 38220 37828 38276 37838
rect 38220 37492 38276 37772
rect 38220 37426 38276 37436
rect 38780 37826 38836 37838
rect 38780 37774 38782 37826
rect 38834 37774 38836 37826
rect 38780 37380 38836 37774
rect 39116 37828 39172 37838
rect 39116 37734 39172 37772
rect 39900 37828 39956 37838
rect 38780 37314 38836 37324
rect 39116 37380 39172 37390
rect 38220 37156 38276 37166
rect 38220 37154 38612 37156
rect 38220 37102 38222 37154
rect 38274 37102 38612 37154
rect 38220 37100 38612 37102
rect 38220 37090 38276 37100
rect 37996 36708 38052 36718
rect 37996 36614 38052 36652
rect 38556 36596 38612 37100
rect 38668 36596 38724 36606
rect 38556 36594 38724 36596
rect 38556 36542 38670 36594
rect 38722 36542 38724 36594
rect 38556 36540 38724 36542
rect 38668 36530 38724 36540
rect 37884 36306 37940 36316
rect 38556 36372 38612 36382
rect 36876 35868 37044 35924
rect 36316 35588 36372 35868
rect 36316 35522 36372 35532
rect 36988 35138 37044 35868
rect 38556 35812 38612 36316
rect 38556 35746 38612 35756
rect 38780 36258 38836 36270
rect 38780 36206 38782 36258
rect 38834 36206 38836 36258
rect 38444 35698 38500 35710
rect 38444 35646 38446 35698
rect 38498 35646 38500 35698
rect 37772 35588 37828 35598
rect 36988 35086 36990 35138
rect 37042 35086 37044 35138
rect 36988 35074 37044 35086
rect 37324 35586 37828 35588
rect 37324 35534 37774 35586
rect 37826 35534 37828 35586
rect 37324 35532 37828 35534
rect 37324 35138 37380 35532
rect 37772 35522 37828 35532
rect 37324 35086 37326 35138
rect 37378 35086 37380 35138
rect 37324 35074 37380 35086
rect 37436 35364 37492 35374
rect 35980 35028 36036 35038
rect 35980 34934 36036 34972
rect 35532 33966 35534 34018
rect 35586 33966 35588 34018
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 34860 33406 34862 33458
rect 34914 33406 34916 33458
rect 34860 33394 34916 33406
rect 35420 33460 35476 33470
rect 35532 33460 35588 33966
rect 35476 33404 35588 33460
rect 35868 34914 35924 34926
rect 35868 34862 35870 34914
rect 35922 34862 35924 34914
rect 35868 34580 35924 34862
rect 35868 33460 35924 34524
rect 36204 34916 36260 34926
rect 36092 33572 36148 33582
rect 36204 33572 36260 34860
rect 36316 34802 36372 34814
rect 36316 34750 36318 34802
rect 36370 34750 36372 34802
rect 36316 34692 36372 34750
rect 36428 34804 36484 34814
rect 36484 34748 36596 34804
rect 36428 34738 36484 34748
rect 36316 34626 36372 34636
rect 36092 33570 36260 33572
rect 36092 33518 36094 33570
rect 36146 33518 36260 33570
rect 36092 33516 36260 33518
rect 36092 33506 36148 33516
rect 35420 33366 35476 33404
rect 35868 33394 35924 33404
rect 36092 33346 36148 33358
rect 36092 33294 36094 33346
rect 36146 33294 36148 33346
rect 35756 33236 35812 33246
rect 35756 33142 35812 33180
rect 36092 33236 36148 33294
rect 36428 33348 36484 33358
rect 36148 33180 36372 33236
rect 36092 33170 36148 33180
rect 34972 32788 35028 32798
rect 34748 32786 35028 32788
rect 34748 32734 34974 32786
rect 35026 32734 35028 32786
rect 34748 32732 35028 32734
rect 34524 31166 34526 31218
rect 34578 31166 34580 31218
rect 34524 31108 34580 31166
rect 34636 31668 34692 31678
rect 34636 31218 34692 31612
rect 34636 31166 34638 31218
rect 34690 31166 34692 31218
rect 34636 31154 34692 31166
rect 34524 31042 34580 31052
rect 34748 31106 34804 32732
rect 34972 32722 35028 32732
rect 36316 32786 36372 33180
rect 36316 32734 36318 32786
rect 36370 32734 36372 32786
rect 36316 32722 36372 32734
rect 35084 32676 35140 32686
rect 34748 31054 34750 31106
rect 34802 31054 34804 31106
rect 34748 31042 34804 31054
rect 34860 32562 34916 32574
rect 34860 32510 34862 32562
rect 34914 32510 34916 32562
rect 34860 31220 34916 32510
rect 34860 30996 34916 31164
rect 34860 30930 34916 30940
rect 35084 30882 35140 32620
rect 36428 32676 36484 33292
rect 36428 32582 36484 32620
rect 35980 32452 36036 32462
rect 35980 32358 36036 32396
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 36428 31778 36484 31790
rect 36428 31726 36430 31778
rect 36482 31726 36484 31778
rect 35644 31668 35700 31678
rect 35644 31574 35700 31612
rect 35084 30830 35086 30882
rect 35138 30830 35140 30882
rect 35084 30818 35140 30830
rect 35756 31108 35812 31118
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35756 30324 35812 31052
rect 33516 30156 34132 30212
rect 32284 29764 32340 29774
rect 32284 29650 32340 29708
rect 32284 29598 32286 29650
rect 32338 29598 32340 29650
rect 32284 29586 32340 29598
rect 32396 28644 32452 28654
rect 32620 28644 32676 30156
rect 32732 30146 32788 30156
rect 33292 30146 33348 30156
rect 33628 29986 33684 29998
rect 33628 29934 33630 29986
rect 33682 29934 33684 29986
rect 33180 29428 33236 29438
rect 33180 29334 33236 29372
rect 33628 29426 33684 29934
rect 34076 29538 34132 30156
rect 34188 30146 34244 30156
rect 34748 30210 34804 30222
rect 34748 30158 34750 30210
rect 34802 30158 34804 30210
rect 34748 29876 34804 30158
rect 34076 29486 34078 29538
rect 34130 29486 34132 29538
rect 34076 29474 34132 29486
rect 34188 29820 34804 29876
rect 33628 29374 33630 29426
rect 33682 29374 33684 29426
rect 33628 29362 33684 29374
rect 33740 29428 33796 29438
rect 32844 28980 32900 28990
rect 32844 28754 32900 28924
rect 32844 28702 32846 28754
rect 32898 28702 32900 28754
rect 32844 28690 32900 28702
rect 33740 28754 33796 29372
rect 33740 28702 33742 28754
rect 33794 28702 33796 28754
rect 33740 28690 33796 28702
rect 34188 28754 34244 29820
rect 34524 29652 34580 29662
rect 34524 29426 34580 29596
rect 34748 29428 34804 29820
rect 34972 30210 35028 30222
rect 34972 30158 34974 30210
rect 35026 30158 35028 30210
rect 34972 29652 35028 30158
rect 35756 30210 35812 30268
rect 35756 30158 35758 30210
rect 35810 30158 35812 30210
rect 35756 30146 35812 30158
rect 35868 30996 35924 31006
rect 35308 29988 35364 29998
rect 35308 29986 35700 29988
rect 35308 29934 35310 29986
rect 35362 29934 35700 29986
rect 35308 29932 35700 29934
rect 35308 29922 35364 29932
rect 34972 29586 35028 29596
rect 34524 29374 34526 29426
rect 34578 29374 34580 29426
rect 34188 28702 34190 28754
rect 34242 28702 34244 28754
rect 34188 28690 34244 28702
rect 34412 28756 34468 28766
rect 34524 28756 34580 29374
rect 34412 28754 34580 28756
rect 34412 28702 34414 28754
rect 34466 28702 34580 28754
rect 34412 28700 34580 28702
rect 34636 29426 34804 29428
rect 34636 29374 34750 29426
rect 34802 29374 34804 29426
rect 34636 29372 34804 29374
rect 35644 29428 35700 29932
rect 35868 29650 35924 30940
rect 36428 30436 36484 31726
rect 36428 30370 36484 30380
rect 35868 29598 35870 29650
rect 35922 29598 35924 29650
rect 35868 29586 35924 29598
rect 36092 30324 36148 30334
rect 35756 29428 35812 29438
rect 35644 29426 35812 29428
rect 35644 29374 35758 29426
rect 35810 29374 35812 29426
rect 35644 29372 35812 29374
rect 34412 28690 34468 28700
rect 32396 28642 32676 28644
rect 32396 28590 32398 28642
rect 32450 28590 32676 28642
rect 32396 28588 32676 28590
rect 33068 28644 33124 28654
rect 32396 28578 32452 28588
rect 33068 28550 33124 28588
rect 34412 28532 34468 28542
rect 32172 28364 32452 28420
rect 32060 27970 32116 27982
rect 32060 27918 32062 27970
rect 32114 27918 32116 27970
rect 31836 27858 31892 27870
rect 31836 27806 31838 27858
rect 31890 27806 31892 27858
rect 31836 27076 31892 27806
rect 31836 27010 31892 27020
rect 32060 26908 32116 27918
rect 32172 27188 32228 27198
rect 32172 27094 32228 27132
rect 31836 26852 31892 26862
rect 32060 26852 32340 26908
rect 31388 26350 31390 26402
rect 31442 26350 31444 26402
rect 31388 26338 31444 26350
rect 31612 26850 31892 26852
rect 31612 26798 31838 26850
rect 31890 26798 31892 26850
rect 31612 26796 31892 26798
rect 31276 25302 31332 25340
rect 31164 24782 31166 24834
rect 31218 24782 31220 24834
rect 30940 24724 30996 24734
rect 30940 24630 30996 24668
rect 30268 23886 30270 23938
rect 30322 23886 30324 23938
rect 30268 23604 30324 23886
rect 30268 23538 30324 23548
rect 30380 24556 30660 24612
rect 29932 22642 29988 22652
rect 30044 22988 30212 23044
rect 30268 23154 30324 23166
rect 30268 23102 30270 23154
rect 30322 23102 30324 23154
rect 30268 23044 30324 23102
rect 29820 20850 29876 20860
rect 29932 21028 29988 21038
rect 29372 20804 29428 20814
rect 29372 20710 29428 20748
rect 29148 19406 29150 19458
rect 29202 19406 29204 19458
rect 29148 19394 29204 19406
rect 29708 19572 29764 19582
rect 29708 19346 29764 19516
rect 29708 19294 29710 19346
rect 29762 19294 29764 19346
rect 29708 19282 29764 19294
rect 29484 19236 29540 19246
rect 28812 19180 29092 19236
rect 29036 18676 29092 19180
rect 29484 19142 29540 19180
rect 29932 18788 29988 20972
rect 30044 20916 30100 22988
rect 30268 22978 30324 22988
rect 30380 21810 30436 24556
rect 31164 24500 31220 24782
rect 30604 24444 31220 24500
rect 31276 25060 31332 25070
rect 30604 23938 30660 24444
rect 31276 24388 31332 25004
rect 31164 24332 31332 24388
rect 31500 24834 31556 24846
rect 31500 24782 31502 24834
rect 31554 24782 31556 24834
rect 30940 24276 30996 24286
rect 30828 24164 30884 24174
rect 30604 23886 30606 23938
rect 30658 23886 30660 23938
rect 30604 23874 30660 23886
rect 30716 24108 30828 24164
rect 30380 21758 30382 21810
rect 30434 21758 30436 21810
rect 30380 21746 30436 21758
rect 30604 22370 30660 22382
rect 30604 22318 30606 22370
rect 30658 22318 30660 22370
rect 30604 21812 30660 22318
rect 30716 22372 30772 24108
rect 30828 24098 30884 24108
rect 30940 24050 30996 24220
rect 30940 23998 30942 24050
rect 30994 23998 30996 24050
rect 30940 23986 30996 23998
rect 30828 23826 30884 23838
rect 30828 23774 30830 23826
rect 30882 23774 30884 23826
rect 30828 23380 30884 23774
rect 30828 23314 30884 23324
rect 30940 23154 30996 23166
rect 30940 23102 30942 23154
rect 30994 23102 30996 23154
rect 30828 23044 30884 23054
rect 30828 22950 30884 22988
rect 30828 22372 30884 22382
rect 30716 22370 30884 22372
rect 30716 22318 30830 22370
rect 30882 22318 30884 22370
rect 30716 22316 30884 22318
rect 30828 22306 30884 22316
rect 30940 21812 30996 23102
rect 31164 23044 31220 24332
rect 31388 24164 31444 24174
rect 31388 24050 31444 24108
rect 31388 23998 31390 24050
rect 31442 23998 31444 24050
rect 31388 23986 31444 23998
rect 31388 23492 31444 23502
rect 31164 22978 31220 22988
rect 31276 23266 31332 23278
rect 31276 23214 31278 23266
rect 31330 23214 31332 23266
rect 31276 21924 31332 23214
rect 31388 22482 31444 23436
rect 31500 23380 31556 24782
rect 31500 23314 31556 23324
rect 31388 22430 31390 22482
rect 31442 22430 31444 22482
rect 31388 22418 31444 22430
rect 31612 22260 31668 26796
rect 31836 26786 31892 26796
rect 32060 26516 32116 26526
rect 32116 26460 32228 26516
rect 32060 26450 32116 26460
rect 31836 26292 31892 26302
rect 31836 26198 31892 26236
rect 32172 26178 32228 26460
rect 32172 26126 32174 26178
rect 32226 26126 32228 26178
rect 32172 26114 32228 26126
rect 31836 25956 31892 25966
rect 31836 24946 31892 25900
rect 32284 25506 32340 26852
rect 32284 25454 32286 25506
rect 32338 25454 32340 25506
rect 31948 25396 32004 25406
rect 32172 25396 32228 25406
rect 32004 25340 32116 25396
rect 31948 25330 32004 25340
rect 31836 24894 31838 24946
rect 31890 24894 31892 24946
rect 31836 24882 31892 24894
rect 31724 24164 31780 24174
rect 31724 23940 31780 24108
rect 32060 24052 32116 25340
rect 32172 25302 32228 25340
rect 32284 24724 32340 25454
rect 32172 24276 32228 24286
rect 32284 24276 32340 24668
rect 32228 24220 32340 24276
rect 32172 24210 32228 24220
rect 32284 24052 32340 24062
rect 32396 24052 32452 28364
rect 33964 28140 34244 28196
rect 33964 28084 34020 28140
rect 33628 28028 34020 28084
rect 33404 27972 33460 27982
rect 33180 27858 33236 27870
rect 33180 27806 33182 27858
rect 33234 27806 33236 27858
rect 33180 26908 33236 27806
rect 33404 27858 33460 27916
rect 33404 27806 33406 27858
rect 33458 27806 33460 27858
rect 33404 27188 33460 27806
rect 33628 27858 33684 28028
rect 34076 27972 34132 27982
rect 34076 27878 34132 27916
rect 34188 27970 34244 28140
rect 34188 27918 34190 27970
rect 34242 27918 34244 27970
rect 34188 27906 34244 27918
rect 33628 27806 33630 27858
rect 33682 27806 33684 27858
rect 33516 27748 33572 27758
rect 33516 27654 33572 27692
rect 33180 26852 33348 26908
rect 32844 26628 32900 26638
rect 32844 26292 32900 26572
rect 32956 26292 33012 26302
rect 32844 26290 33012 26292
rect 32844 26238 32958 26290
rect 33010 26238 33012 26290
rect 32844 26236 33012 26238
rect 33292 26292 33348 26852
rect 33404 26514 33460 27132
rect 33404 26462 33406 26514
rect 33458 26462 33460 26514
rect 33404 26450 33460 26462
rect 33516 26292 33572 26302
rect 33292 26290 33572 26292
rect 33292 26238 33518 26290
rect 33570 26238 33572 26290
rect 33292 26236 33572 26238
rect 32844 26180 32900 26236
rect 32956 26226 33012 26236
rect 33516 26226 33572 26236
rect 33628 26292 33684 27806
rect 33628 26198 33684 26236
rect 33852 27858 33908 27870
rect 33852 27806 33854 27858
rect 33906 27806 33908 27858
rect 32060 23996 32228 24052
rect 31724 23938 31892 23940
rect 31724 23886 31726 23938
rect 31778 23886 31892 23938
rect 31724 23884 31892 23886
rect 31724 23874 31780 23884
rect 31724 23268 31780 23278
rect 31724 23174 31780 23212
rect 31724 22596 31780 22606
rect 31724 22482 31780 22540
rect 31724 22430 31726 22482
rect 31778 22430 31780 22482
rect 31724 22418 31780 22430
rect 31612 22204 31780 22260
rect 31276 21858 31332 21868
rect 31500 22148 31556 22158
rect 30604 21756 30996 21812
rect 30492 21700 30548 21710
rect 30492 21606 30548 21644
rect 30604 21588 30660 21598
rect 30156 20916 30212 20926
rect 30604 20916 30660 21532
rect 30044 20914 30212 20916
rect 30044 20862 30158 20914
rect 30210 20862 30212 20914
rect 30044 20860 30212 20862
rect 30156 20850 30212 20860
rect 30492 20860 30660 20916
rect 30716 21586 30772 21598
rect 30716 21534 30718 21586
rect 30770 21534 30772 21586
rect 30492 20244 30548 20860
rect 30716 20804 30772 21534
rect 30828 21140 30884 21756
rect 31052 21588 31108 21598
rect 31052 21494 31108 21532
rect 31500 21474 31556 22092
rect 31500 21422 31502 21474
rect 31554 21422 31556 21474
rect 31500 21410 31556 21422
rect 30828 21084 31108 21140
rect 30716 20738 30772 20748
rect 30604 20690 30660 20702
rect 30604 20638 30606 20690
rect 30658 20638 30660 20690
rect 30604 20468 30660 20638
rect 30604 20402 30660 20412
rect 30268 20242 30548 20244
rect 30268 20190 30494 20242
rect 30546 20190 30548 20242
rect 30268 20188 30548 20190
rect 30156 20020 30212 20030
rect 30268 20020 30324 20188
rect 30156 20018 30324 20020
rect 30156 19966 30158 20018
rect 30210 19966 30324 20018
rect 30156 19964 30324 19966
rect 30156 19954 30212 19964
rect 30156 19348 30212 19358
rect 30156 19254 30212 19292
rect 30268 18900 30324 18910
rect 29932 18732 30100 18788
rect 28812 18620 29092 18676
rect 28588 18338 28756 18340
rect 28588 18286 28590 18338
rect 28642 18286 28756 18338
rect 28588 18284 28756 18286
rect 28588 18274 28644 18284
rect 28476 18060 28644 18116
rect 28588 17666 28644 18060
rect 28588 17614 28590 17666
rect 28642 17614 28644 17666
rect 28588 17602 28644 17614
rect 28476 17556 28532 17566
rect 28420 17554 28532 17556
rect 28420 17502 28478 17554
rect 28530 17502 28532 17554
rect 28420 17500 28532 17502
rect 28364 17462 28420 17500
rect 28476 17490 28532 17500
rect 27356 17276 28084 17332
rect 28252 17442 28308 17454
rect 28252 17390 28254 17442
rect 28306 17390 28308 17442
rect 27132 17154 27188 17164
rect 26796 17052 26964 17108
rect 27692 17108 27748 17118
rect 26796 16660 26852 17052
rect 27020 16996 27076 17006
rect 27020 16994 27188 16996
rect 27020 16942 27022 16994
rect 27074 16942 27188 16994
rect 27020 16940 27188 16942
rect 27020 16930 27076 16940
rect 26908 16884 26964 16894
rect 26908 16790 26964 16828
rect 27132 16660 27188 16940
rect 27356 16940 27636 16996
rect 26796 16604 26964 16660
rect 26684 16370 26740 16380
rect 26796 16324 26852 16334
rect 26012 16156 26292 16212
rect 26684 16210 26740 16222
rect 26684 16158 26686 16210
rect 26738 16158 26740 16210
rect 25900 15988 25956 15998
rect 25900 15894 25956 15932
rect 25788 15874 25844 15886
rect 25788 15822 25790 15874
rect 25842 15822 25844 15874
rect 25788 15428 25844 15822
rect 26012 15652 26068 16156
rect 26124 15986 26180 15998
rect 26124 15934 26126 15986
rect 26178 15934 26180 15986
rect 26124 15764 26180 15934
rect 26124 15708 26628 15764
rect 26012 15596 26180 15652
rect 26012 15428 26068 15438
rect 25788 15426 26068 15428
rect 25788 15374 26014 15426
rect 26066 15374 26068 15426
rect 25788 15372 26068 15374
rect 26012 15362 26068 15372
rect 26124 15204 26180 15596
rect 26012 15148 26180 15204
rect 26012 14868 26068 15148
rect 25788 14532 25844 14542
rect 25788 14418 25844 14476
rect 25788 14366 25790 14418
rect 25842 14366 25844 14418
rect 25788 14354 25844 14366
rect 26012 14196 26068 14812
rect 26460 14868 26516 14878
rect 25676 14018 25732 14028
rect 25788 14140 26068 14196
rect 26124 14530 26180 14542
rect 26124 14478 26126 14530
rect 26178 14478 26180 14530
rect 25564 13806 25566 13858
rect 25618 13806 25620 13858
rect 25564 13636 25620 13806
rect 25788 13748 25844 14140
rect 26124 13972 26180 14478
rect 26460 14530 26516 14812
rect 26572 14642 26628 15708
rect 26684 15148 26740 16158
rect 26796 15986 26852 16268
rect 26796 15934 26798 15986
rect 26850 15934 26852 15986
rect 26796 15922 26852 15934
rect 26908 15148 26964 16604
rect 27132 16594 27188 16604
rect 27244 16882 27300 16894
rect 27244 16830 27246 16882
rect 27298 16830 27300 16882
rect 27020 16324 27076 16334
rect 27244 16324 27300 16830
rect 27020 16322 27300 16324
rect 27020 16270 27022 16322
rect 27074 16270 27300 16322
rect 27020 16268 27300 16270
rect 27020 16258 27076 16268
rect 27244 15540 27300 16268
rect 27244 15474 27300 15484
rect 27356 15428 27412 16940
rect 26684 15092 26852 15148
rect 26908 15092 27300 15148
rect 26572 14590 26574 14642
rect 26626 14590 26628 14642
rect 26572 14578 26628 14590
rect 26460 14478 26462 14530
rect 26514 14478 26516 14530
rect 26460 14466 26516 14478
rect 26684 14308 26740 14318
rect 26684 14214 26740 14252
rect 26124 13906 26180 13916
rect 26572 14196 26628 14206
rect 26572 13970 26628 14140
rect 26796 14084 26852 15092
rect 27132 14980 27188 14990
rect 27132 14642 27188 14924
rect 27132 14590 27134 14642
rect 27186 14590 27188 14642
rect 27132 14578 27188 14590
rect 26572 13918 26574 13970
rect 26626 13918 26628 13970
rect 26572 13906 26628 13918
rect 26684 14028 26852 14084
rect 25900 13748 25956 13758
rect 25788 13746 25956 13748
rect 25788 13694 25902 13746
rect 25954 13694 25956 13746
rect 25788 13692 25956 13694
rect 25564 13570 25620 13580
rect 25676 13634 25732 13646
rect 25676 13582 25678 13634
rect 25730 13582 25732 13634
rect 25676 13524 25732 13582
rect 25900 13524 25956 13692
rect 26124 13748 26180 13758
rect 26124 13746 26516 13748
rect 26124 13694 26126 13746
rect 26178 13694 26516 13746
rect 26124 13692 26516 13694
rect 26124 13682 26180 13692
rect 26236 13524 26292 13534
rect 25900 13522 26292 13524
rect 25900 13470 26238 13522
rect 26290 13470 26292 13522
rect 25900 13468 26292 13470
rect 25676 13458 25732 13468
rect 26236 13458 26292 13468
rect 26348 13524 26404 13534
rect 25676 13300 25732 13310
rect 25732 13244 25956 13300
rect 25676 13234 25732 13244
rect 25228 12964 25284 12974
rect 25228 12870 25284 12908
rect 25340 12404 25396 12414
rect 25340 12310 25396 12348
rect 25116 11282 25172 12124
rect 25676 12178 25732 12190
rect 25676 12126 25678 12178
rect 25730 12126 25732 12178
rect 25116 11230 25118 11282
rect 25170 11230 25172 11282
rect 25116 11218 25172 11230
rect 25340 11396 25396 11406
rect 25676 11396 25732 12126
rect 25900 11506 25956 13244
rect 26348 12404 26404 13468
rect 26348 12310 26404 12348
rect 26460 12402 26516 13692
rect 26460 12350 26462 12402
rect 26514 12350 26516 12402
rect 26460 12338 26516 12350
rect 26572 13300 26628 13310
rect 26572 12402 26628 13244
rect 26572 12350 26574 12402
rect 26626 12350 26628 12402
rect 26572 12338 26628 12350
rect 26012 12292 26068 12302
rect 26012 12198 26068 12236
rect 25900 11454 25902 11506
rect 25954 11454 25956 11506
rect 25900 11442 25956 11454
rect 26124 12180 26180 12190
rect 26684 12180 26740 14028
rect 27020 13636 27076 13646
rect 27020 13542 27076 13580
rect 25340 11394 25732 11396
rect 25340 11342 25342 11394
rect 25394 11342 25732 11394
rect 25340 11340 25732 11342
rect 25340 11284 25396 11340
rect 25340 11218 25396 11228
rect 26124 10722 26180 12124
rect 26572 12124 26740 12180
rect 26796 12628 26852 12638
rect 26348 12068 26404 12078
rect 26348 11506 26404 12012
rect 26348 11454 26350 11506
rect 26402 11454 26404 11506
rect 26348 11442 26404 11454
rect 26460 11956 26516 11966
rect 26124 10670 26126 10722
rect 26178 10670 26180 10722
rect 26124 10658 26180 10670
rect 26348 10724 26404 10734
rect 25676 10612 25732 10622
rect 25564 10610 25732 10612
rect 25564 10558 25678 10610
rect 25730 10558 25732 10610
rect 25564 10556 25732 10558
rect 25228 10500 25284 10510
rect 25228 10406 25284 10444
rect 25564 9716 25620 10556
rect 25676 10546 25732 10556
rect 26236 10498 26292 10510
rect 26236 10446 26238 10498
rect 26290 10446 26292 10498
rect 26236 10052 26292 10446
rect 25676 9996 26292 10052
rect 25676 9938 25732 9996
rect 25676 9886 25678 9938
rect 25730 9886 25732 9938
rect 25676 9874 25732 9886
rect 26348 9828 26404 10668
rect 26124 9772 26404 9828
rect 26460 10722 26516 11900
rect 26460 10670 26462 10722
rect 26514 10670 26516 10722
rect 25564 9660 25732 9716
rect 24556 9548 25508 9604
rect 24556 9266 24612 9548
rect 24556 9214 24558 9266
rect 24610 9214 24612 9266
rect 24556 9202 24612 9214
rect 25452 9266 25508 9548
rect 25452 9214 25454 9266
rect 25506 9214 25508 9266
rect 25452 9202 25508 9214
rect 25564 9380 25620 9390
rect 24668 8818 24724 8830
rect 24668 8766 24670 8818
rect 24722 8766 24724 8818
rect 24668 8484 24724 8766
rect 24556 7476 24612 7486
rect 24556 7382 24612 7420
rect 24556 7028 24612 7038
rect 23884 6078 23886 6130
rect 23938 6078 23940 6130
rect 23884 6066 23940 6078
rect 23996 6690 24388 6692
rect 23996 6638 24222 6690
rect 24274 6638 24388 6690
rect 23996 6636 24388 6638
rect 24444 6972 24556 7028
rect 23772 5908 23828 5918
rect 23772 5346 23828 5852
rect 23772 5294 23774 5346
rect 23826 5294 23828 5346
rect 23772 5282 23828 5294
rect 23884 5572 23940 5582
rect 23884 5124 23940 5516
rect 23996 5348 24052 6636
rect 24220 6626 24276 6636
rect 24332 6132 24388 6142
rect 24444 6132 24500 6972
rect 24556 6962 24612 6972
rect 24332 6130 24500 6132
rect 24332 6078 24334 6130
rect 24386 6078 24500 6130
rect 24332 6076 24500 6078
rect 24108 5908 24164 5918
rect 24108 5814 24164 5852
rect 24220 5794 24276 5806
rect 24220 5742 24222 5794
rect 24274 5742 24276 5794
rect 24220 5348 24276 5742
rect 24332 5572 24388 6076
rect 24556 6020 24612 6030
rect 24556 5926 24612 5964
rect 24332 5506 24388 5516
rect 24556 5684 24612 5694
rect 24332 5348 24388 5358
rect 23996 5292 24164 5348
rect 24220 5346 24388 5348
rect 24220 5294 24334 5346
rect 24386 5294 24388 5346
rect 24220 5292 24388 5294
rect 23996 5124 24052 5134
rect 23884 5122 24052 5124
rect 23884 5070 23998 5122
rect 24050 5070 24052 5122
rect 23884 5068 24052 5070
rect 23996 5058 24052 5068
rect 23660 4946 23716 4956
rect 24108 4564 24164 5292
rect 24332 5282 24388 5292
rect 24444 5348 24500 5358
rect 24444 5254 24500 5292
rect 23660 4228 23716 4238
rect 23660 4134 23716 4172
rect 24108 3668 24164 4508
rect 24556 4562 24612 5628
rect 24556 4510 24558 4562
rect 24610 4510 24612 4562
rect 24556 4498 24612 4510
rect 24164 3612 24612 3668
rect 24108 3574 24164 3612
rect 23660 3556 23716 3566
rect 23548 3554 23716 3556
rect 23548 3502 23662 3554
rect 23714 3502 23716 3554
rect 23548 3500 23716 3502
rect 21084 3332 21364 3388
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 21084 2884 21140 3332
rect 21084 2818 21140 2828
rect 23660 3220 23716 3500
rect 24556 3554 24612 3612
rect 24556 3502 24558 3554
rect 24610 3502 24612 3554
rect 24556 3490 24612 3502
rect 24668 3388 24724 8428
rect 25116 7588 25172 7598
rect 25004 7364 25060 7374
rect 24892 6692 24948 6702
rect 24892 6598 24948 6636
rect 25004 6468 25060 7308
rect 24892 6412 25060 6468
rect 24780 5460 24836 5470
rect 24780 5010 24836 5404
rect 24780 4958 24782 5010
rect 24834 4958 24836 5010
rect 24780 4946 24836 4958
rect 18508 2482 18564 2492
rect 23660 2548 23716 3164
rect 23660 2482 23716 2492
rect 24556 3332 24724 3388
rect 24556 1428 24612 3332
rect 24892 1652 24948 6412
rect 25116 5906 25172 7532
rect 25564 7476 25620 9324
rect 25676 9268 25732 9660
rect 25676 9202 25732 9212
rect 26012 9268 26068 9278
rect 26012 9174 26068 9212
rect 25900 8260 25956 8270
rect 25900 8166 25956 8204
rect 25788 7588 25844 7598
rect 25788 7494 25844 7532
rect 25564 7474 25732 7476
rect 25564 7422 25566 7474
rect 25618 7422 25732 7474
rect 25564 7420 25732 7422
rect 25564 7410 25620 7420
rect 25676 6132 25732 7420
rect 26124 7364 26180 9772
rect 26460 9268 26516 10670
rect 26572 10052 26628 12124
rect 26796 11394 26852 12572
rect 27020 12292 27076 12302
rect 27020 12178 27076 12236
rect 27020 12126 27022 12178
rect 27074 12126 27076 12178
rect 27020 12114 27076 12126
rect 26796 11342 26798 11394
rect 26850 11342 26852 11394
rect 26796 11330 26852 11342
rect 26908 11170 26964 11182
rect 26908 11118 26910 11170
rect 26962 11118 26964 11170
rect 26684 10724 26740 10734
rect 26908 10724 26964 11118
rect 27020 11172 27076 11182
rect 27020 11170 27188 11172
rect 27020 11118 27022 11170
rect 27074 11118 27188 11170
rect 27020 11116 27188 11118
rect 27020 11106 27076 11116
rect 26684 10722 26964 10724
rect 26684 10670 26686 10722
rect 26738 10670 26964 10722
rect 26684 10668 26964 10670
rect 26684 10658 26740 10668
rect 27132 10052 27188 11116
rect 27244 10388 27300 15092
rect 27356 13412 27412 15372
rect 27468 16772 27524 16782
rect 27468 15316 27524 16716
rect 27580 16770 27636 16940
rect 27580 16718 27582 16770
rect 27634 16718 27636 16770
rect 27580 16706 27636 16718
rect 27692 16770 27748 17052
rect 27692 16718 27694 16770
rect 27746 16718 27748 16770
rect 27692 16706 27748 16718
rect 27916 16660 27972 16670
rect 27916 16566 27972 16604
rect 28028 16658 28084 16670
rect 28028 16606 28030 16658
rect 28082 16606 28084 16658
rect 27468 15250 27524 15260
rect 27580 16436 27636 16446
rect 27580 14756 27636 16380
rect 28028 16212 28084 16606
rect 28252 16324 28308 17390
rect 28700 17108 28756 18284
rect 28588 17052 28756 17108
rect 28364 16994 28420 17006
rect 28364 16942 28366 16994
rect 28418 16942 28420 16994
rect 28364 16660 28420 16942
rect 28364 16594 28420 16604
rect 28476 16884 28532 16894
rect 28252 16268 28420 16324
rect 27692 16156 28084 16212
rect 27692 16098 27748 16156
rect 27692 16046 27694 16098
rect 27746 16046 27748 16098
rect 27692 16034 27748 16046
rect 28028 16100 28084 16156
rect 28252 16100 28308 16110
rect 28028 16098 28308 16100
rect 28028 16046 28254 16098
rect 28306 16046 28308 16098
rect 28028 16044 28308 16046
rect 28252 16034 28308 16044
rect 27916 15876 27972 15886
rect 27916 15782 27972 15820
rect 28364 15540 28420 16268
rect 28252 15484 28420 15540
rect 27580 14642 27636 14700
rect 28140 15202 28196 15214
rect 28140 15150 28142 15202
rect 28194 15150 28196 15202
rect 28140 14868 28196 15150
rect 27580 14590 27582 14642
rect 27634 14590 27636 14642
rect 27580 14578 27636 14590
rect 28028 14644 28084 14654
rect 28028 14550 28084 14588
rect 27692 14532 27748 14542
rect 27468 13748 27524 13758
rect 27468 13654 27524 13692
rect 27356 13346 27412 13356
rect 27356 13188 27412 13198
rect 27356 13074 27412 13132
rect 27356 13022 27358 13074
rect 27410 13022 27412 13074
rect 27356 13010 27412 13022
rect 27692 12964 27748 14476
rect 28140 14532 28196 14812
rect 28140 14466 28196 14476
rect 27916 13636 27972 13646
rect 27804 13634 27972 13636
rect 27804 13582 27918 13634
rect 27970 13582 27972 13634
rect 27804 13580 27972 13582
rect 27804 13522 27860 13580
rect 27916 13570 27972 13580
rect 27804 13470 27806 13522
rect 27858 13470 27860 13522
rect 27804 13458 27860 13470
rect 28028 13522 28084 13534
rect 28028 13470 28030 13522
rect 28082 13470 28084 13522
rect 28028 12964 28084 13470
rect 28140 13076 28196 13086
rect 28140 12982 28196 13020
rect 27580 12962 28084 12964
rect 27580 12910 28030 12962
rect 28082 12910 28084 12962
rect 27580 12908 28084 12910
rect 27468 12292 27524 12302
rect 27468 11394 27524 12236
rect 27580 12290 27636 12908
rect 28028 12898 28084 12908
rect 28252 12740 28308 15484
rect 27580 12238 27582 12290
rect 27634 12238 27636 12290
rect 27580 12180 27636 12238
rect 27580 12114 27636 12124
rect 27692 12684 28308 12740
rect 28364 15316 28420 15326
rect 28364 12962 28420 15260
rect 28476 14754 28532 16828
rect 28588 16772 28644 17052
rect 28812 16996 28868 18620
rect 29932 18564 29988 18574
rect 29036 18452 29092 18462
rect 29596 18452 29652 18462
rect 29036 18450 29428 18452
rect 29036 18398 29038 18450
rect 29090 18398 29428 18450
rect 29036 18396 29428 18398
rect 29036 18386 29092 18396
rect 29260 18228 29316 18238
rect 29148 17892 29204 17902
rect 29148 17668 29204 17836
rect 29036 17666 29204 17668
rect 29036 17614 29150 17666
rect 29202 17614 29204 17666
rect 29036 17612 29204 17614
rect 28812 16930 28868 16940
rect 28924 17332 28980 17342
rect 28588 16706 28644 16716
rect 28700 16884 28756 16894
rect 28588 15874 28644 15886
rect 28588 15822 28590 15874
rect 28642 15822 28644 15874
rect 28588 15764 28644 15822
rect 28588 15698 28644 15708
rect 28588 15314 28644 15326
rect 28588 15262 28590 15314
rect 28642 15262 28644 15314
rect 28588 14868 28644 15262
rect 28588 14802 28644 14812
rect 28700 14980 28756 16828
rect 28924 16884 28980 17276
rect 28924 16818 28980 16828
rect 29036 16660 29092 17612
rect 29148 17602 29204 17612
rect 29148 17108 29204 17118
rect 29260 17108 29316 18172
rect 29372 17556 29428 18396
rect 29596 18358 29652 18396
rect 29932 18338 29988 18508
rect 29932 18286 29934 18338
rect 29986 18286 29988 18338
rect 29484 17556 29540 17566
rect 29372 17554 29540 17556
rect 29372 17502 29486 17554
rect 29538 17502 29540 17554
rect 29372 17500 29540 17502
rect 29148 17106 29316 17108
rect 29148 17054 29150 17106
rect 29202 17054 29316 17106
rect 29148 17052 29316 17054
rect 29484 17108 29540 17500
rect 29820 17108 29876 17118
rect 29484 17106 29876 17108
rect 29484 17054 29486 17106
rect 29538 17054 29822 17106
rect 29874 17054 29876 17106
rect 29484 17052 29876 17054
rect 29148 17042 29204 17052
rect 29484 17042 29540 17052
rect 28476 14702 28478 14754
rect 28530 14702 28532 14754
rect 28476 14690 28532 14702
rect 28588 14644 28644 14654
rect 28476 13972 28532 13982
rect 28588 13972 28644 14588
rect 28476 13970 28644 13972
rect 28476 13918 28478 13970
rect 28530 13918 28644 13970
rect 28476 13916 28644 13918
rect 28700 13972 28756 14924
rect 28476 13906 28532 13916
rect 28700 13906 28756 13916
rect 28812 16604 29092 16660
rect 29148 16772 29204 16782
rect 28812 13970 28868 16604
rect 29148 16324 29204 16716
rect 28812 13918 28814 13970
rect 28866 13918 28868 13970
rect 28812 13906 28868 13918
rect 28924 16268 29204 16324
rect 28364 12910 28366 12962
rect 28418 12910 28420 12962
rect 27468 11342 27470 11394
rect 27522 11342 27524 11394
rect 27468 11330 27524 11342
rect 27356 10836 27412 10846
rect 27356 10610 27412 10780
rect 27356 10558 27358 10610
rect 27410 10558 27412 10610
rect 27356 10546 27412 10558
rect 27244 10322 27300 10332
rect 26572 9996 27076 10052
rect 26460 9174 26516 9212
rect 26796 9156 26852 9166
rect 26348 8148 26404 8158
rect 26348 8054 26404 8092
rect 26460 8034 26516 8046
rect 26460 7982 26462 8034
rect 26514 7982 26516 8034
rect 26348 7588 26404 7598
rect 26124 7298 26180 7308
rect 26236 7532 26348 7588
rect 26124 6132 26180 6142
rect 25676 6076 25956 6132
rect 25564 6020 25620 6030
rect 25564 5926 25620 5964
rect 25116 5854 25118 5906
rect 25170 5854 25172 5906
rect 25116 5842 25172 5854
rect 25340 5908 25396 5918
rect 25788 5908 25844 5918
rect 25340 5814 25396 5852
rect 25676 5852 25788 5908
rect 25340 5124 25396 5134
rect 25676 5124 25732 5852
rect 25788 5814 25844 5852
rect 25340 5122 25732 5124
rect 25340 5070 25342 5122
rect 25394 5070 25732 5122
rect 25340 5068 25732 5070
rect 25788 5124 25844 5134
rect 25340 5058 25396 5068
rect 25788 5030 25844 5068
rect 25004 5012 25060 5022
rect 25004 4918 25060 4956
rect 25116 4898 25172 4910
rect 25116 4846 25118 4898
rect 25170 4846 25172 4898
rect 25116 4452 25172 4846
rect 25788 4564 25844 4574
rect 25900 4564 25956 6076
rect 26124 6038 26180 6076
rect 26236 5908 26292 7532
rect 26348 7522 26404 7532
rect 26460 7476 26516 7982
rect 26572 8036 26628 8046
rect 26572 7586 26628 7980
rect 26572 7534 26574 7586
rect 26626 7534 26628 7586
rect 26572 7522 26628 7534
rect 26460 7410 26516 7420
rect 26348 7364 26404 7374
rect 26348 7270 26404 7308
rect 26684 7362 26740 7374
rect 26684 7310 26686 7362
rect 26738 7310 26740 7362
rect 26684 6692 26740 7310
rect 26684 6626 26740 6636
rect 26796 6132 26852 9100
rect 27020 9042 27076 9996
rect 27132 9986 27188 9996
rect 27244 9156 27300 9166
rect 27244 9154 27524 9156
rect 27244 9102 27246 9154
rect 27298 9102 27524 9154
rect 27244 9100 27524 9102
rect 27244 9090 27300 9100
rect 27020 8990 27022 9042
rect 27074 8990 27076 9042
rect 27020 8708 27076 8990
rect 27020 8642 27076 8652
rect 27132 8036 27188 8046
rect 27020 7980 27132 8036
rect 26908 7474 26964 7486
rect 26908 7422 26910 7474
rect 26962 7422 26964 7474
rect 26908 6916 26964 7422
rect 27020 7140 27076 7980
rect 27132 7970 27188 7980
rect 27468 7586 27524 9100
rect 27580 8372 27636 8382
rect 27580 7698 27636 8316
rect 27580 7646 27582 7698
rect 27634 7646 27636 7698
rect 27580 7634 27636 7646
rect 27468 7534 27470 7586
rect 27522 7534 27524 7586
rect 27132 7476 27188 7486
rect 27132 7474 27300 7476
rect 27132 7422 27134 7474
rect 27186 7422 27300 7474
rect 27132 7420 27300 7422
rect 27132 7410 27188 7420
rect 27020 7084 27188 7140
rect 26908 6850 26964 6860
rect 26348 5908 26404 5918
rect 26236 5906 26404 5908
rect 26236 5854 26350 5906
rect 26402 5854 26404 5906
rect 26236 5852 26404 5854
rect 26348 5842 26404 5852
rect 26460 5236 26516 5246
rect 26460 5142 26516 5180
rect 25788 4562 25956 4564
rect 25788 4510 25790 4562
rect 25842 4510 25956 4562
rect 25788 4508 25956 4510
rect 26236 4564 26292 4574
rect 25228 4452 25284 4462
rect 25116 4450 25284 4452
rect 25116 4398 25230 4450
rect 25282 4398 25284 4450
rect 25116 4396 25284 4398
rect 25228 4386 25284 4396
rect 25340 4114 25396 4126
rect 25340 4062 25342 4114
rect 25394 4062 25396 4114
rect 25340 3666 25396 4062
rect 25340 3614 25342 3666
rect 25394 3614 25396 3666
rect 25340 3602 25396 3614
rect 24892 1586 24948 1596
rect 24556 1362 24612 1372
rect 15036 1250 15092 1260
rect 25788 1316 25844 4508
rect 26236 3668 26292 4508
rect 26796 4562 26852 6076
rect 27020 6802 27076 6814
rect 27020 6750 27022 6802
rect 27074 6750 27076 6802
rect 27020 6356 27076 6750
rect 27020 6020 27076 6300
rect 27020 5954 27076 5964
rect 27132 6804 27188 7084
rect 27244 6916 27300 7420
rect 27468 7364 27524 7534
rect 27468 7298 27524 7308
rect 27244 6860 27524 6916
rect 27132 6018 27188 6748
rect 27468 6802 27524 6860
rect 27468 6750 27470 6802
rect 27522 6750 27524 6802
rect 27468 6738 27524 6750
rect 27356 6692 27412 6702
rect 27356 6598 27412 6636
rect 27580 6578 27636 6590
rect 27580 6526 27582 6578
rect 27634 6526 27636 6578
rect 27580 6468 27636 6526
rect 27356 6412 27636 6468
rect 27356 6356 27412 6412
rect 27356 6290 27412 6300
rect 27692 6244 27748 12684
rect 27804 12404 27860 12414
rect 27804 12402 28084 12404
rect 27804 12350 27806 12402
rect 27858 12350 28084 12402
rect 27804 12348 28084 12350
rect 27804 12338 27860 12348
rect 27916 12178 27972 12190
rect 27916 12126 27918 12178
rect 27970 12126 27972 12178
rect 27916 11844 27972 12126
rect 27916 11778 27972 11788
rect 27804 11172 27860 11182
rect 27804 11078 27860 11116
rect 28028 10722 28084 12348
rect 28140 12180 28196 12190
rect 28140 12086 28196 12124
rect 28364 11788 28420 12910
rect 28588 12850 28644 12862
rect 28588 12798 28590 12850
rect 28642 12798 28644 12850
rect 28476 12404 28532 12414
rect 28476 12310 28532 12348
rect 28588 12402 28644 12798
rect 28588 12350 28590 12402
rect 28642 12350 28644 12402
rect 28588 12338 28644 12350
rect 28700 12516 28756 12526
rect 28700 12402 28756 12460
rect 28700 12350 28702 12402
rect 28754 12350 28756 12402
rect 28700 12338 28756 12350
rect 28140 11732 28420 11788
rect 28140 11172 28196 11732
rect 28140 11106 28196 11116
rect 28252 11170 28308 11182
rect 28252 11118 28254 11170
rect 28306 11118 28308 11170
rect 28252 11060 28308 11118
rect 28252 11004 28532 11060
rect 28028 10670 28030 10722
rect 28082 10670 28084 10722
rect 28028 10658 28084 10670
rect 28140 10836 28196 10846
rect 27804 10388 27860 10398
rect 27860 10332 27972 10388
rect 27804 10322 27860 10332
rect 27804 10052 27860 10062
rect 27804 9938 27860 9996
rect 27804 9886 27806 9938
rect 27858 9886 27860 9938
rect 27804 9874 27860 9886
rect 27804 9268 27860 9278
rect 27916 9268 27972 10332
rect 28140 10052 28196 10780
rect 27804 9266 27972 9268
rect 27804 9214 27806 9266
rect 27858 9214 27972 9266
rect 27804 9212 27972 9214
rect 28028 9996 28196 10052
rect 27804 9202 27860 9212
rect 27916 8818 27972 8830
rect 27916 8766 27918 8818
rect 27970 8766 27972 8818
rect 27804 8708 27860 8718
rect 27804 8258 27860 8652
rect 27804 8206 27806 8258
rect 27858 8206 27860 8258
rect 27804 8194 27860 8206
rect 27804 7700 27860 7710
rect 27804 7606 27860 7644
rect 27916 7476 27972 8766
rect 27804 7420 27972 7476
rect 28028 7474 28084 9996
rect 28476 9940 28532 11004
rect 28476 9884 28644 9940
rect 28252 9826 28308 9838
rect 28252 9774 28254 9826
rect 28306 9774 28308 9826
rect 28252 9716 28308 9774
rect 28140 9660 28252 9716
rect 28140 9266 28196 9660
rect 28252 9650 28308 9660
rect 28588 9828 28644 9884
rect 28140 9214 28142 9266
rect 28194 9214 28196 9266
rect 28140 8820 28196 9214
rect 28140 8754 28196 8764
rect 28476 9604 28532 9614
rect 28476 8818 28532 9548
rect 28588 9266 28644 9772
rect 28588 9214 28590 9266
rect 28642 9214 28644 9266
rect 28588 9202 28644 9214
rect 28476 8766 28478 8818
rect 28530 8766 28532 8818
rect 28476 8754 28532 8766
rect 28588 8372 28644 8382
rect 28588 8278 28644 8316
rect 28140 8036 28196 8046
rect 28140 7942 28196 7980
rect 28924 7812 28980 16268
rect 29596 16098 29652 17052
rect 29820 17042 29876 17052
rect 29596 16046 29598 16098
rect 29650 16046 29652 16098
rect 29596 16034 29652 16046
rect 29372 15988 29428 15998
rect 29372 15894 29428 15932
rect 29260 15202 29316 15214
rect 29260 15150 29262 15202
rect 29314 15150 29316 15202
rect 29260 14642 29316 15150
rect 29932 15148 29988 18286
rect 30044 16884 30100 18732
rect 30044 16818 30100 16828
rect 30156 17666 30212 17678
rect 30156 17614 30158 17666
rect 30210 17614 30212 17666
rect 29932 15092 30100 15148
rect 29260 14590 29262 14642
rect 29314 14590 29316 14642
rect 29260 14578 29316 14590
rect 29708 14756 29764 14766
rect 29036 14530 29092 14542
rect 29036 14478 29038 14530
rect 29090 14478 29092 14530
rect 29036 13522 29092 14478
rect 29372 14530 29428 14542
rect 29372 14478 29374 14530
rect 29426 14478 29428 14530
rect 29372 14196 29428 14478
rect 29708 14530 29764 14700
rect 29708 14478 29710 14530
rect 29762 14478 29764 14530
rect 29708 14466 29764 14478
rect 29372 14130 29428 14140
rect 29372 13972 29428 13982
rect 29372 13878 29428 13916
rect 30044 13972 30100 15092
rect 30156 14868 30212 17614
rect 30268 16548 30324 18844
rect 30380 18450 30436 20188
rect 30492 20178 30548 20188
rect 30940 20356 30996 20366
rect 30828 19684 30884 19694
rect 30492 19236 30548 19246
rect 30492 19142 30548 19180
rect 30380 18398 30382 18450
rect 30434 18398 30436 18450
rect 30380 18386 30436 18398
rect 30828 18450 30884 19628
rect 30940 19346 30996 20300
rect 31052 19906 31108 21084
rect 31612 20802 31668 20814
rect 31612 20750 31614 20802
rect 31666 20750 31668 20802
rect 31164 20690 31220 20702
rect 31164 20638 31166 20690
rect 31218 20638 31220 20690
rect 31164 20468 31220 20638
rect 31164 20402 31220 20412
rect 31052 19854 31054 19906
rect 31106 19854 31108 19906
rect 31052 19572 31108 19854
rect 31052 19506 31108 19516
rect 31388 20018 31444 20030
rect 31388 19966 31390 20018
rect 31442 19966 31444 20018
rect 30940 19294 30942 19346
rect 30994 19294 30996 19346
rect 30940 19282 30996 19294
rect 31276 19348 31332 19358
rect 30828 18398 30830 18450
rect 30882 18398 30884 18450
rect 30828 18386 30884 18398
rect 31164 18450 31220 18462
rect 31164 18398 31166 18450
rect 31218 18398 31220 18450
rect 31164 17780 31220 18398
rect 31276 18228 31332 19292
rect 31388 18452 31444 19966
rect 31612 19236 31668 20750
rect 31724 19460 31780 22204
rect 31836 21586 31892 23884
rect 31836 21534 31838 21586
rect 31890 21534 31892 21586
rect 31836 20580 31892 21534
rect 32060 23380 32116 23390
rect 32060 20914 32116 23324
rect 32172 21810 32228 23996
rect 32284 24050 32452 24052
rect 32284 23998 32286 24050
rect 32338 23998 32452 24050
rect 32284 23996 32452 23998
rect 32284 23986 32340 23996
rect 32172 21758 32174 21810
rect 32226 21758 32228 21810
rect 32172 21746 32228 21758
rect 32284 21924 32340 21934
rect 32396 21924 32452 23996
rect 32508 24610 32564 24622
rect 32508 24558 32510 24610
rect 32562 24558 32564 24610
rect 32508 24052 32564 24558
rect 32508 23986 32564 23996
rect 32732 24164 32788 24174
rect 32732 24050 32788 24108
rect 32732 23998 32734 24050
rect 32786 23998 32788 24050
rect 32732 23986 32788 23998
rect 32508 23156 32564 23166
rect 32508 23062 32564 23100
rect 32396 21868 32676 21924
rect 32284 21700 32340 21868
rect 32396 21700 32452 21710
rect 32284 21698 32452 21700
rect 32284 21646 32398 21698
rect 32450 21646 32452 21698
rect 32284 21644 32452 21646
rect 32284 21252 32340 21644
rect 32396 21634 32452 21644
rect 32508 21588 32564 21598
rect 32508 21494 32564 21532
rect 32060 20862 32062 20914
rect 32114 20862 32116 20914
rect 32060 20850 32116 20862
rect 32172 21196 32340 21252
rect 31836 20514 31892 20524
rect 32060 20578 32116 20590
rect 32060 20526 32062 20578
rect 32114 20526 32116 20578
rect 31836 20356 31892 20366
rect 32060 20356 32116 20526
rect 32172 20356 32228 21196
rect 32620 21028 32676 21868
rect 32844 21812 32900 26124
rect 33068 25396 33124 25406
rect 33068 24836 33124 25340
rect 33628 25396 33684 25406
rect 33852 25396 33908 27806
rect 34300 27748 34356 27758
rect 34300 27186 34356 27692
rect 34300 27134 34302 27186
rect 34354 27134 34356 27186
rect 34300 27122 34356 27134
rect 33628 25394 33908 25396
rect 33628 25342 33630 25394
rect 33682 25342 33908 25394
rect 33628 25340 33908 25342
rect 33964 26740 34020 26750
rect 33516 25282 33572 25294
rect 33516 25230 33518 25282
rect 33570 25230 33572 25282
rect 33516 25172 33572 25230
rect 33516 25106 33572 25116
rect 33068 24050 33124 24780
rect 33628 24722 33684 25340
rect 33740 24836 33796 24846
rect 33964 24836 34020 26684
rect 34076 26180 34132 26190
rect 34076 26086 34132 26124
rect 34412 25732 34468 28476
rect 34636 27746 34692 29372
rect 34748 29362 34804 29372
rect 35756 29362 35812 29372
rect 35420 29316 35476 29326
rect 35420 29314 35588 29316
rect 35420 29262 35422 29314
rect 35474 29262 35588 29314
rect 35420 29260 35588 29262
rect 35420 29250 35476 29260
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 34748 28868 34804 28878
rect 34748 28774 34804 28812
rect 35308 28644 35364 28654
rect 35532 28644 35588 29260
rect 35308 28642 35588 28644
rect 35308 28590 35310 28642
rect 35362 28590 35588 28642
rect 35308 28588 35588 28590
rect 35644 28644 35700 28654
rect 35868 28644 35924 28654
rect 35644 28642 35812 28644
rect 35644 28590 35646 28642
rect 35698 28590 35812 28642
rect 35644 28588 35812 28590
rect 35308 28532 35364 28588
rect 35644 28578 35700 28588
rect 35308 28466 35364 28476
rect 35532 28418 35588 28430
rect 35532 28366 35534 28418
rect 35586 28366 35588 28418
rect 35532 28196 35588 28366
rect 35532 28130 35588 28140
rect 35756 28420 35812 28588
rect 35868 28550 35924 28588
rect 34636 27694 34638 27746
rect 34690 27694 34692 27746
rect 34636 27682 34692 27694
rect 34636 27524 34692 27534
rect 34524 26178 34580 26190
rect 34524 26126 34526 26178
rect 34578 26126 34580 26178
rect 34524 25956 34580 26126
rect 34524 25890 34580 25900
rect 34524 25732 34580 25742
rect 34412 25676 34524 25732
rect 34524 25506 34580 25676
rect 34524 25454 34526 25506
rect 34578 25454 34580 25506
rect 34524 25442 34580 25454
rect 33740 24834 34020 24836
rect 33740 24782 33742 24834
rect 33794 24782 34020 24834
rect 33740 24780 34020 24782
rect 34300 25284 34356 25294
rect 33740 24770 33796 24780
rect 33628 24670 33630 24722
rect 33682 24670 33684 24722
rect 33628 24658 33684 24670
rect 34300 24722 34356 25228
rect 34300 24670 34302 24722
rect 34354 24670 34356 24722
rect 34300 24658 34356 24670
rect 33852 24612 33908 24622
rect 33852 24518 33908 24556
rect 33068 23998 33070 24050
rect 33122 23998 33124 24050
rect 33068 23986 33124 23998
rect 34524 23604 34580 23614
rect 32956 23154 33012 23166
rect 33404 23156 33460 23166
rect 32956 23102 32958 23154
rect 33010 23102 33012 23154
rect 32956 22708 33012 23102
rect 32956 22036 33012 22652
rect 32956 21970 33012 21980
rect 33068 23154 33460 23156
rect 33068 23102 33406 23154
rect 33458 23102 33460 23154
rect 33068 23100 33460 23102
rect 32844 21756 33012 21812
rect 32508 20972 32676 21028
rect 32284 20804 32340 20814
rect 32284 20710 32340 20748
rect 32508 20468 32564 20972
rect 32620 20804 32676 20814
rect 32620 20802 32900 20804
rect 32620 20750 32622 20802
rect 32674 20750 32900 20802
rect 32620 20748 32900 20750
rect 32620 20738 32676 20748
rect 32508 20412 32788 20468
rect 32060 20300 32676 20356
rect 31836 20130 31892 20300
rect 31836 20078 31838 20130
rect 31890 20078 31892 20130
rect 31836 20066 31892 20078
rect 32060 20020 32116 20030
rect 32060 20018 32228 20020
rect 32060 19966 32062 20018
rect 32114 19966 32228 20018
rect 32060 19964 32228 19966
rect 32060 19954 32116 19964
rect 31948 19906 32004 19918
rect 31948 19854 31950 19906
rect 32002 19854 32004 19906
rect 31948 19796 32004 19854
rect 31724 19394 31780 19404
rect 31836 19740 32004 19796
rect 32060 19796 32116 19806
rect 31612 19170 31668 19180
rect 31500 19124 31556 19134
rect 31500 18674 31556 19068
rect 31500 18622 31502 18674
rect 31554 18622 31556 18674
rect 31500 18610 31556 18622
rect 31836 18562 31892 19740
rect 31836 18510 31838 18562
rect 31890 18510 31892 18562
rect 31836 18498 31892 18510
rect 31948 18564 32004 18574
rect 31388 18386 31444 18396
rect 31500 18450 31556 18462
rect 31500 18398 31502 18450
rect 31554 18398 31556 18450
rect 31276 18172 31444 18228
rect 30716 17724 31164 17780
rect 30716 16994 30772 17724
rect 31164 17686 31220 17724
rect 30828 17554 30884 17566
rect 30828 17502 30830 17554
rect 30882 17502 30884 17554
rect 30828 17106 30884 17502
rect 30828 17054 30830 17106
rect 30882 17054 30884 17106
rect 30828 17042 30884 17054
rect 30716 16942 30718 16994
rect 30770 16942 30772 16994
rect 30716 16930 30772 16942
rect 30940 16882 30996 16894
rect 30940 16830 30942 16882
rect 30994 16830 30996 16882
rect 30380 16772 30436 16782
rect 30380 16678 30436 16716
rect 30268 16492 30660 16548
rect 30268 16100 30324 16110
rect 30268 16006 30324 16044
rect 30156 14802 30212 14812
rect 30380 15874 30436 15886
rect 30380 15822 30382 15874
rect 30434 15822 30436 15874
rect 30380 14756 30436 15822
rect 30380 14690 30436 14700
rect 30492 15874 30548 15886
rect 30492 15822 30494 15874
rect 30546 15822 30548 15874
rect 30492 15092 30548 15822
rect 30492 14532 30548 15036
rect 29820 13636 29876 13646
rect 29036 13470 29038 13522
rect 29090 13470 29092 13522
rect 29036 13458 29092 13470
rect 29708 13634 29876 13636
rect 29708 13582 29822 13634
rect 29874 13582 29876 13634
rect 29708 13580 29876 13582
rect 29148 12962 29204 12974
rect 29148 12910 29150 12962
rect 29202 12910 29204 12962
rect 29036 12292 29092 12302
rect 29036 12178 29092 12236
rect 29036 12126 29038 12178
rect 29090 12126 29092 12178
rect 29036 12114 29092 12126
rect 29148 10836 29204 12910
rect 29372 12404 29428 12414
rect 29372 12310 29428 12348
rect 29484 12180 29540 12190
rect 29484 12086 29540 12124
rect 29596 12178 29652 12190
rect 29596 12126 29598 12178
rect 29650 12126 29652 12178
rect 29260 11844 29316 11854
rect 29260 11172 29316 11788
rect 29260 11170 29540 11172
rect 29260 11118 29262 11170
rect 29314 11118 29540 11170
rect 29260 11116 29540 11118
rect 29260 11106 29316 11116
rect 29260 10836 29316 10846
rect 29148 10780 29260 10836
rect 29260 9826 29316 10780
rect 29260 9774 29262 9826
rect 29314 9774 29316 9826
rect 29260 9762 29316 9774
rect 29372 10276 29428 10286
rect 29372 9380 29428 10220
rect 29484 10164 29540 11116
rect 29596 10388 29652 12126
rect 29708 11844 29764 13580
rect 29820 13570 29876 13580
rect 29932 13076 29988 13086
rect 29932 12982 29988 13020
rect 29820 12292 29876 12302
rect 29820 12198 29876 12236
rect 29708 11778 29764 11788
rect 30044 11844 30100 13916
rect 30268 14476 30548 14532
rect 30044 11778 30100 11788
rect 30156 12180 30212 12190
rect 29708 11396 29764 11406
rect 29708 11302 29764 11340
rect 30156 10724 30212 12124
rect 30156 10658 30212 10668
rect 29596 10322 29652 10332
rect 30044 10500 30100 10510
rect 29484 10108 29652 10164
rect 29372 9314 29428 9324
rect 29484 9268 29540 9278
rect 29148 9156 29204 9166
rect 29148 9062 29204 9100
rect 29484 9154 29540 9212
rect 29484 9102 29486 9154
rect 29538 9102 29540 9154
rect 29484 9090 29540 9102
rect 29596 9044 29652 10108
rect 29932 9716 29988 9726
rect 29708 9714 29988 9716
rect 29708 9662 29934 9714
rect 29986 9662 29988 9714
rect 29708 9660 29988 9662
rect 29708 9266 29764 9660
rect 29932 9650 29988 9660
rect 29708 9214 29710 9266
rect 29762 9214 29764 9266
rect 29708 9202 29764 9214
rect 29820 9156 29876 9166
rect 29820 9062 29876 9100
rect 30044 9154 30100 10444
rect 30156 10498 30212 10510
rect 30156 10446 30158 10498
rect 30210 10446 30212 10498
rect 30156 10388 30212 10446
rect 30156 10322 30212 10332
rect 30268 9492 30324 14476
rect 30380 14306 30436 14318
rect 30380 14254 30382 14306
rect 30434 14254 30436 14306
rect 30380 14196 30436 14254
rect 30380 14130 30436 14140
rect 30380 13748 30436 13758
rect 30604 13748 30660 16492
rect 30828 16100 30884 16110
rect 30828 16006 30884 16044
rect 30940 15148 30996 16830
rect 31276 16884 31332 16894
rect 31276 16790 31332 16828
rect 31388 16210 31444 18172
rect 31500 18004 31556 18398
rect 31500 17938 31556 17948
rect 31948 17106 32004 18508
rect 32060 18452 32116 19740
rect 32172 19012 32228 19964
rect 32508 19908 32564 19918
rect 32508 19814 32564 19852
rect 32396 19794 32452 19806
rect 32396 19742 32398 19794
rect 32450 19742 32452 19794
rect 32396 19236 32452 19742
rect 32620 19684 32676 20300
rect 32396 19170 32452 19180
rect 32508 19628 32676 19684
rect 32228 18956 32340 19012
rect 32172 18946 32228 18956
rect 32172 18452 32228 18462
rect 32060 18450 32228 18452
rect 32060 18398 32174 18450
rect 32226 18398 32228 18450
rect 32060 18396 32228 18398
rect 32172 18386 32228 18396
rect 31948 17054 31950 17106
rect 32002 17054 32004 17106
rect 31948 17042 32004 17054
rect 32172 17108 32228 17118
rect 32284 17108 32340 18956
rect 32508 18562 32564 19628
rect 32508 18510 32510 18562
rect 32562 18510 32564 18562
rect 32508 18498 32564 18510
rect 32172 17106 32340 17108
rect 32172 17054 32174 17106
rect 32226 17054 32340 17106
rect 32172 17052 32340 17054
rect 32172 17042 32228 17052
rect 31388 16158 31390 16210
rect 31442 16158 31444 16210
rect 31388 16146 31444 16158
rect 31500 16882 31556 16894
rect 31500 16830 31502 16882
rect 31554 16830 31556 16882
rect 31500 16772 31556 16830
rect 32060 16884 32116 16894
rect 32060 16790 32116 16828
rect 31388 15202 31444 15214
rect 31388 15150 31390 15202
rect 31442 15150 31444 15202
rect 31388 15148 31444 15150
rect 30716 15092 30996 15148
rect 31164 15092 31444 15148
rect 30716 14196 30772 15092
rect 31164 15026 31220 15036
rect 31500 14980 31556 16716
rect 32732 16100 32788 20412
rect 32844 19796 32900 20748
rect 32844 19730 32900 19740
rect 32956 19572 33012 21756
rect 33068 21476 33124 23100
rect 33404 23090 33460 23100
rect 33628 23154 33684 23166
rect 34412 23156 34468 23166
rect 33628 23102 33630 23154
rect 33682 23102 33684 23154
rect 33516 23042 33572 23054
rect 33516 22990 33518 23042
rect 33570 22990 33572 23042
rect 33516 22372 33572 22990
rect 33628 22484 33684 23102
rect 34076 23154 34468 23156
rect 34076 23102 34414 23154
rect 34466 23102 34468 23154
rect 34076 23100 34468 23102
rect 33964 23044 34020 23054
rect 33964 22950 34020 22988
rect 33628 22428 34020 22484
rect 33180 22316 33572 22372
rect 33180 21586 33236 22316
rect 33852 22260 33908 22270
rect 33516 22258 33908 22260
rect 33516 22206 33854 22258
rect 33906 22206 33908 22258
rect 33516 22204 33908 22206
rect 33516 21810 33572 22204
rect 33852 22194 33908 22204
rect 33516 21758 33518 21810
rect 33570 21758 33572 21810
rect 33516 21746 33572 21758
rect 33628 22036 33684 22046
rect 33180 21534 33182 21586
rect 33234 21534 33236 21586
rect 33180 21522 33236 21534
rect 33292 21586 33348 21598
rect 33292 21534 33294 21586
rect 33346 21534 33348 21586
rect 33068 21410 33124 21420
rect 33292 21476 33348 21534
rect 33292 21410 33348 21420
rect 33628 21028 33684 21980
rect 33516 20972 33684 21028
rect 33740 21588 33796 21598
rect 33964 21588 34020 22428
rect 33740 21586 34020 21588
rect 33740 21534 33742 21586
rect 33794 21534 34020 21586
rect 33740 21532 34020 21534
rect 33180 20916 33236 20926
rect 33180 20822 33236 20860
rect 33516 20018 33572 20972
rect 33516 19966 33518 20018
rect 33570 19966 33572 20018
rect 33516 19954 33572 19966
rect 33628 20802 33684 20814
rect 33628 20750 33630 20802
rect 33682 20750 33684 20802
rect 32620 15988 32676 15998
rect 31276 14924 31556 14980
rect 31612 15876 31668 15886
rect 31612 15314 31668 15820
rect 31724 15874 31780 15886
rect 31724 15822 31726 15874
rect 31778 15822 31780 15874
rect 31724 15652 31780 15822
rect 31948 15876 32004 15886
rect 31948 15782 32004 15820
rect 32060 15874 32116 15886
rect 32060 15822 32062 15874
rect 32114 15822 32116 15874
rect 31724 15596 32004 15652
rect 31612 15262 31614 15314
rect 31666 15262 31668 15314
rect 30828 14868 30884 14878
rect 30828 14532 30884 14812
rect 30828 14530 30996 14532
rect 30828 14478 30830 14530
rect 30882 14478 30996 14530
rect 30828 14476 30996 14478
rect 30828 14466 30884 14476
rect 30828 14196 30884 14206
rect 30716 14140 30828 14196
rect 30828 13970 30884 14140
rect 30828 13918 30830 13970
rect 30882 13918 30884 13970
rect 30828 13906 30884 13918
rect 30380 13746 30660 13748
rect 30380 13694 30382 13746
rect 30434 13694 30660 13746
rect 30380 13692 30660 13694
rect 30380 12068 30436 13692
rect 30828 12178 30884 12190
rect 30828 12126 30830 12178
rect 30882 12126 30884 12178
rect 30492 12068 30548 12078
rect 30380 12066 30660 12068
rect 30380 12014 30494 12066
rect 30546 12014 30660 12066
rect 30380 12012 30660 12014
rect 30492 12002 30548 12012
rect 30604 11956 30660 12012
rect 30604 11900 30772 11956
rect 30492 11844 30548 11854
rect 30492 11172 30548 11788
rect 30268 9426 30324 9436
rect 30380 11170 30548 11172
rect 30380 11118 30494 11170
rect 30546 11118 30548 11170
rect 30380 11116 30548 11118
rect 30044 9102 30046 9154
rect 30098 9102 30100 9154
rect 30044 9090 30100 9102
rect 29596 8978 29652 8988
rect 30380 8820 30436 11116
rect 30492 11106 30548 11116
rect 30716 10948 30772 11900
rect 30828 11844 30884 12126
rect 30828 11778 30884 11788
rect 30492 10892 30772 10948
rect 30828 11396 30884 11406
rect 30492 8932 30548 10892
rect 30828 10836 30884 11340
rect 30604 10780 30884 10836
rect 30940 11394 30996 14476
rect 31276 13746 31332 14924
rect 31612 14868 31668 15262
rect 31836 15202 31892 15214
rect 31836 15150 31838 15202
rect 31890 15150 31892 15202
rect 31836 15148 31892 15150
rect 31276 13694 31278 13746
rect 31330 13694 31332 13746
rect 31164 13636 31220 13646
rect 31276 13636 31332 13694
rect 31388 14812 31668 14868
rect 31724 15092 31892 15148
rect 31948 15204 32004 15596
rect 32060 15540 32116 15822
rect 32172 15874 32228 15886
rect 32172 15822 32174 15874
rect 32226 15822 32228 15874
rect 32172 15764 32228 15822
rect 32228 15708 32340 15764
rect 32172 15698 32228 15708
rect 32060 15484 32228 15540
rect 32060 15316 32116 15326
rect 32060 15222 32116 15260
rect 32172 15314 32228 15484
rect 32172 15262 32174 15314
rect 32226 15262 32228 15314
rect 32172 15250 32228 15262
rect 31948 15138 32004 15148
rect 31388 13748 31444 14812
rect 31724 14756 31780 15092
rect 31500 14700 31780 14756
rect 31500 14642 31556 14700
rect 31500 14590 31502 14642
rect 31554 14590 31556 14642
rect 31500 14578 31556 14590
rect 31612 14084 31668 14094
rect 31612 13970 31668 14028
rect 31612 13918 31614 13970
rect 31666 13918 31668 13970
rect 31612 13906 31668 13918
rect 31388 13692 31668 13748
rect 31220 13580 31332 13636
rect 31164 13570 31220 13580
rect 31164 12404 31220 12414
rect 30940 11342 30942 11394
rect 30994 11342 30996 11394
rect 30940 10836 30996 11342
rect 30604 10722 30660 10780
rect 30604 10670 30606 10722
rect 30658 10670 30660 10722
rect 30604 10658 30660 10670
rect 30828 10612 30884 10622
rect 30828 10518 30884 10556
rect 30716 10500 30772 10510
rect 30716 10406 30772 10444
rect 30940 10500 30996 10780
rect 30940 10434 30996 10444
rect 31052 12068 31108 12078
rect 31052 10276 31108 12012
rect 31164 10948 31220 12348
rect 31612 12402 31668 13692
rect 32060 13634 32116 13646
rect 32060 13582 32062 13634
rect 32114 13582 32116 13634
rect 32060 13524 32116 13582
rect 32060 13458 32116 13468
rect 32060 13074 32116 13086
rect 32060 13022 32062 13074
rect 32114 13022 32116 13074
rect 32060 12516 32116 13022
rect 32060 12450 32116 12460
rect 31612 12350 31614 12402
rect 31666 12350 31668 12402
rect 31276 12292 31332 12302
rect 31276 12198 31332 12236
rect 31388 12290 31444 12302
rect 31388 12238 31390 12290
rect 31442 12238 31444 12290
rect 31388 11620 31444 12238
rect 31388 11554 31444 11564
rect 31500 12066 31556 12078
rect 31500 12014 31502 12066
rect 31554 12014 31556 12066
rect 31500 11508 31556 12014
rect 31612 12068 31668 12350
rect 31836 12292 31892 12302
rect 31836 12198 31892 12236
rect 32060 12290 32116 12302
rect 32060 12238 32062 12290
rect 32114 12238 32116 12290
rect 31612 12002 31668 12012
rect 31612 11508 31668 11518
rect 31500 11506 31668 11508
rect 31500 11454 31614 11506
rect 31666 11454 31668 11506
rect 31500 11452 31668 11454
rect 31612 11442 31668 11452
rect 31948 11396 32004 11406
rect 31836 11340 31948 11396
rect 31164 10892 31556 10948
rect 30604 10220 31108 10276
rect 31164 10610 31220 10622
rect 31164 10558 31166 10610
rect 31218 10558 31220 10610
rect 30604 9268 30660 10220
rect 30604 9154 30660 9212
rect 30828 9716 30884 9726
rect 30828 9266 30884 9660
rect 31164 9604 31220 10558
rect 31164 9380 31220 9548
rect 30828 9214 30830 9266
rect 30882 9214 30884 9266
rect 30828 9202 30884 9214
rect 31052 9324 31220 9380
rect 30604 9102 30606 9154
rect 30658 9102 30660 9154
rect 30604 9090 30660 9102
rect 30828 9044 30884 9054
rect 30492 8876 30772 8932
rect 30380 8764 30548 8820
rect 29708 8260 29764 8270
rect 29764 8204 29876 8260
rect 29708 8194 29764 8204
rect 29484 8146 29540 8158
rect 29484 8094 29486 8146
rect 29538 8094 29540 8146
rect 29148 8036 29204 8046
rect 29148 7942 29204 7980
rect 29260 8034 29316 8046
rect 29260 7982 29262 8034
rect 29314 7982 29316 8034
rect 28028 7422 28030 7474
rect 28082 7422 28084 7474
rect 27804 6578 27860 7420
rect 28028 6692 28084 7422
rect 28700 7756 28980 7812
rect 28364 6916 28420 6926
rect 28364 6802 28420 6860
rect 28364 6750 28366 6802
rect 28418 6750 28420 6802
rect 28364 6738 28420 6750
rect 27804 6526 27806 6578
rect 27858 6526 27860 6578
rect 27804 6468 27860 6526
rect 27804 6402 27860 6412
rect 27916 6580 27972 6590
rect 27580 6188 27748 6244
rect 27132 5966 27134 6018
rect 27186 5966 27188 6018
rect 27132 5954 27188 5966
rect 27356 6132 27412 6142
rect 27356 5906 27412 6076
rect 27356 5854 27358 5906
rect 27410 5854 27412 5906
rect 27356 5842 27412 5854
rect 27244 5794 27300 5806
rect 27244 5742 27246 5794
rect 27298 5742 27300 5794
rect 27244 5236 27300 5742
rect 27468 5796 27524 5806
rect 27468 5348 27524 5740
rect 27244 5170 27300 5180
rect 27356 5292 27524 5348
rect 26796 4510 26798 4562
rect 26850 4510 26852 4562
rect 26796 4498 26852 4510
rect 27356 3668 27412 5292
rect 27468 5124 27524 5134
rect 27468 4338 27524 5068
rect 27468 4286 27470 4338
rect 27522 4286 27524 4338
rect 27468 4274 27524 4286
rect 27468 3668 27524 3678
rect 27356 3666 27524 3668
rect 27356 3614 27470 3666
rect 27522 3614 27524 3666
rect 27356 3612 27524 3614
rect 26236 3602 26292 3612
rect 27468 3602 27524 3612
rect 27580 2772 27636 6188
rect 27692 6018 27748 6030
rect 27692 5966 27694 6018
rect 27746 5966 27748 6018
rect 27692 5908 27748 5966
rect 27804 5908 27860 5918
rect 27692 5852 27804 5908
rect 27804 5842 27860 5852
rect 27916 5906 27972 6524
rect 27916 5854 27918 5906
rect 27970 5854 27972 5906
rect 27916 5842 27972 5854
rect 28028 5124 28084 6636
rect 28364 6132 28420 6142
rect 28028 5058 28084 5068
rect 28140 5796 28196 5806
rect 28140 4450 28196 5740
rect 28364 5684 28420 6076
rect 28588 6020 28644 6030
rect 28588 5926 28644 5964
rect 28476 5908 28532 5918
rect 28476 5814 28532 5852
rect 28364 5628 28644 5684
rect 28588 5234 28644 5628
rect 28588 5182 28590 5234
rect 28642 5182 28644 5234
rect 28588 5170 28644 5182
rect 28140 4398 28142 4450
rect 28194 4398 28196 4450
rect 28140 4386 28196 4398
rect 28588 3668 28644 3678
rect 28588 3574 28644 3612
rect 28700 3388 28756 7756
rect 29260 7700 29316 7982
rect 29372 8036 29428 8046
rect 29372 7942 29428 7980
rect 28812 7644 29316 7700
rect 29484 7700 29540 8094
rect 28812 7586 28868 7644
rect 29484 7634 29540 7644
rect 29596 8148 29652 8158
rect 28812 7534 28814 7586
rect 28866 7534 28868 7586
rect 28812 7522 28868 7534
rect 29596 7252 29652 8092
rect 29596 7186 29652 7196
rect 28812 6804 28868 6814
rect 28812 5906 28868 6748
rect 29484 6466 29540 6478
rect 29484 6414 29486 6466
rect 29538 6414 29540 6466
rect 29484 6244 29540 6414
rect 29260 6188 29484 6244
rect 28812 5854 28814 5906
rect 28866 5854 28868 5906
rect 28812 5842 28868 5854
rect 29148 6020 29204 6030
rect 29036 5796 29092 5806
rect 29036 5702 29092 5740
rect 29148 5122 29204 5964
rect 29260 6018 29316 6188
rect 29484 6178 29540 6188
rect 29596 6468 29652 6478
rect 29260 5966 29262 6018
rect 29314 5966 29316 6018
rect 29260 5954 29316 5966
rect 29372 5906 29428 5918
rect 29372 5854 29374 5906
rect 29426 5854 29428 5906
rect 29260 5236 29316 5246
rect 29372 5236 29428 5854
rect 29260 5234 29428 5236
rect 29260 5182 29262 5234
rect 29314 5182 29428 5234
rect 29260 5180 29428 5182
rect 29260 5170 29316 5180
rect 29148 5070 29150 5122
rect 29202 5070 29204 5122
rect 29148 5058 29204 5070
rect 29596 5124 29652 6412
rect 29820 6132 29876 8204
rect 30380 8146 30436 8158
rect 30380 8094 30382 8146
rect 30434 8094 30436 8146
rect 30268 8036 30324 8046
rect 30268 7942 30324 7980
rect 30380 7700 30436 8094
rect 30492 8148 30548 8764
rect 30492 8082 30548 8092
rect 30380 7634 30436 7644
rect 30268 7476 30324 7486
rect 29932 6692 29988 6702
rect 29988 6636 30212 6692
rect 29932 6598 29988 6636
rect 29932 6132 29988 6142
rect 29820 6130 29988 6132
rect 29820 6078 29934 6130
rect 29986 6078 29988 6130
rect 29820 6076 29988 6078
rect 29932 6066 29988 6076
rect 30156 5236 30212 6636
rect 30268 6690 30324 7420
rect 30268 6638 30270 6690
rect 30322 6638 30324 6690
rect 30268 6244 30324 6638
rect 30268 6178 30324 6188
rect 30380 7364 30436 7374
rect 30380 5906 30436 7308
rect 30492 6692 30548 6702
rect 30492 6466 30548 6636
rect 30492 6414 30494 6466
rect 30546 6414 30548 6466
rect 30492 6402 30548 6414
rect 30604 6578 30660 6590
rect 30604 6526 30606 6578
rect 30658 6526 30660 6578
rect 30604 6132 30660 6526
rect 30604 6066 30660 6076
rect 30380 5854 30382 5906
rect 30434 5854 30436 5906
rect 30380 5842 30436 5854
rect 30604 5908 30660 5918
rect 30604 5814 30660 5852
rect 30716 5572 30772 8876
rect 30828 8034 30884 8988
rect 31052 8932 31108 9324
rect 31164 9156 31220 9166
rect 31164 9062 31220 9100
rect 31388 9042 31444 9054
rect 31388 8990 31390 9042
rect 31442 8990 31444 9042
rect 31388 8932 31444 8990
rect 31052 8876 31444 8932
rect 31276 8148 31332 8158
rect 31276 8054 31332 8092
rect 30828 7982 30830 8034
rect 30882 7982 30884 8034
rect 30828 7140 30884 7982
rect 30940 7700 30996 7710
rect 30996 7644 31444 7700
rect 30940 7362 30996 7644
rect 31388 7586 31444 7644
rect 31388 7534 31390 7586
rect 31442 7534 31444 7586
rect 31388 7522 31444 7534
rect 31276 7476 31332 7486
rect 31276 7382 31332 7420
rect 30940 7310 30942 7362
rect 30994 7310 30996 7362
rect 30940 7298 30996 7310
rect 31500 7252 31556 10892
rect 31836 10164 31892 11340
rect 31948 11330 32004 11340
rect 32060 10836 32116 12238
rect 32172 12292 32228 12302
rect 32284 12292 32340 15708
rect 32620 15148 32676 15932
rect 32508 15092 32676 15148
rect 32508 14196 32564 15092
rect 32172 12290 32340 12292
rect 32172 12238 32174 12290
rect 32226 12238 32340 12290
rect 32172 12236 32340 12238
rect 32396 14084 32452 14094
rect 32172 11396 32228 12236
rect 32172 11330 32228 11340
rect 32060 10780 32340 10836
rect 32060 10612 32116 10622
rect 31948 10500 32004 10510
rect 31948 10406 32004 10444
rect 31836 10108 32004 10164
rect 31948 9716 32004 10108
rect 32060 9938 32116 10556
rect 32060 9886 32062 9938
rect 32114 9886 32116 9938
rect 32060 9874 32116 9886
rect 32172 10500 32228 10510
rect 31948 9660 32116 9716
rect 32060 9266 32116 9660
rect 32060 9214 32062 9266
rect 32114 9214 32116 9266
rect 32060 9202 32116 9214
rect 31948 9156 32004 9166
rect 31948 9062 32004 9100
rect 31836 9044 31892 9054
rect 31836 8950 31892 8988
rect 32060 8372 32116 8382
rect 32172 8372 32228 10444
rect 32284 8932 32340 10780
rect 32396 10834 32452 14028
rect 32508 12852 32564 14140
rect 32620 13076 32676 13086
rect 32732 13076 32788 16044
rect 32844 19516 33012 19572
rect 33180 19906 33236 19918
rect 33180 19854 33182 19906
rect 33234 19854 33236 19906
rect 32844 15204 32900 19516
rect 33180 19236 33236 19854
rect 33180 19170 33236 19180
rect 33068 19124 33124 19134
rect 33068 19030 33124 19068
rect 32956 19012 33012 19022
rect 32956 18788 33012 18956
rect 33516 19012 33572 19022
rect 32956 18732 33124 18788
rect 33068 18676 33124 18732
rect 33068 18674 33236 18676
rect 33068 18622 33070 18674
rect 33122 18622 33236 18674
rect 33068 18620 33236 18622
rect 33068 18610 33124 18620
rect 32956 18564 33012 18574
rect 32956 17778 33012 18508
rect 32956 17726 32958 17778
rect 33010 17726 33012 17778
rect 32956 17714 33012 17726
rect 33180 17444 33236 18620
rect 33404 18562 33460 18574
rect 33404 18510 33406 18562
rect 33458 18510 33460 18562
rect 33292 17780 33348 17790
rect 33404 17780 33460 18510
rect 33348 17724 33460 17780
rect 33292 17666 33348 17724
rect 33292 17614 33294 17666
rect 33346 17614 33348 17666
rect 33292 17602 33348 17614
rect 33404 17556 33460 17566
rect 33516 17556 33572 18956
rect 33628 18564 33684 20750
rect 33740 20020 33796 21532
rect 33964 21364 34020 21374
rect 33964 20802 34020 21308
rect 34076 21140 34132 23100
rect 34412 23090 34468 23100
rect 34524 22372 34580 23548
rect 34076 21074 34132 21084
rect 34188 22370 34580 22372
rect 34188 22318 34526 22370
rect 34578 22318 34580 22370
rect 34188 22316 34580 22318
rect 34188 21586 34244 22316
rect 34524 22306 34580 22316
rect 34188 21534 34190 21586
rect 34242 21534 34244 21586
rect 34188 20916 34244 21534
rect 34636 21252 34692 27468
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35084 27076 35140 27086
rect 35084 26982 35140 27020
rect 35756 26402 35812 28364
rect 35756 26350 35758 26402
rect 35810 26350 35812 26402
rect 35756 26338 35812 26350
rect 34972 26290 35028 26302
rect 34972 26238 34974 26290
rect 35026 26238 35028 26290
rect 34972 26180 35028 26238
rect 35420 26292 35476 26302
rect 35420 26198 35476 26236
rect 35868 26290 35924 26302
rect 35868 26238 35870 26290
rect 35922 26238 35924 26290
rect 34972 26114 35028 26124
rect 35868 26068 35924 26238
rect 35868 26002 35924 26012
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35980 25732 36036 25742
rect 35980 25618 36036 25676
rect 35980 25566 35982 25618
rect 36034 25566 36036 25618
rect 35980 25554 36036 25566
rect 34972 25508 35028 25518
rect 34972 25414 35028 25452
rect 36092 25508 36148 30268
rect 36540 30212 36596 34748
rect 37212 34692 37268 34702
rect 37212 34598 37268 34636
rect 37324 34244 37380 34254
rect 37436 34244 37492 35308
rect 37212 34242 37492 34244
rect 37212 34190 37326 34242
rect 37378 34190 37492 34242
rect 37212 34188 37492 34190
rect 37996 34916 38052 34926
rect 38444 34916 38500 35646
rect 38780 35364 38836 36206
rect 39116 35924 39172 37324
rect 39900 37044 39956 37772
rect 40348 37828 40404 39004
rect 40348 37826 40516 37828
rect 40348 37774 40350 37826
rect 40402 37774 40516 37826
rect 40348 37772 40516 37774
rect 40348 37762 40404 37772
rect 40348 37156 40404 37166
rect 40348 37062 40404 37100
rect 39900 36988 40292 37044
rect 40236 36932 40292 36988
rect 40236 36876 40404 36932
rect 39228 36482 39284 36494
rect 39228 36430 39230 36482
rect 39282 36430 39284 36482
rect 39228 36372 39284 36430
rect 39340 36484 39396 36494
rect 39340 36390 39396 36428
rect 39676 36484 39732 36494
rect 39676 36390 39732 36428
rect 39228 36306 39284 36316
rect 39564 36258 39620 36270
rect 39564 36206 39566 36258
rect 39618 36206 39620 36258
rect 39564 36148 39620 36206
rect 39564 36082 39620 36092
rect 40124 36258 40180 36270
rect 40124 36206 40126 36258
rect 40178 36206 40180 36258
rect 39340 35924 39396 35934
rect 39116 35868 39284 35924
rect 38892 35812 38948 35822
rect 38892 35718 38948 35756
rect 39116 35698 39172 35710
rect 39116 35646 39118 35698
rect 39170 35646 39172 35698
rect 38780 35298 38836 35308
rect 39004 35586 39060 35598
rect 39004 35534 39006 35586
rect 39058 35534 39060 35586
rect 39004 35140 39060 35534
rect 38668 35084 39060 35140
rect 38668 35026 38724 35084
rect 38668 34974 38670 35026
rect 38722 34974 38724 35026
rect 38668 34962 38724 34974
rect 37996 34914 38500 34916
rect 37996 34862 37998 34914
rect 38050 34862 38500 34914
rect 37996 34860 38500 34862
rect 37100 34018 37156 34030
rect 37100 33966 37102 34018
rect 37154 33966 37156 34018
rect 36988 33236 37044 33246
rect 36988 33142 37044 33180
rect 37100 32788 37156 33966
rect 37212 33124 37268 34188
rect 37324 34178 37380 34188
rect 37996 33572 38052 34860
rect 38668 34242 38724 34254
rect 38668 34190 38670 34242
rect 38722 34190 38724 34242
rect 38444 34132 38500 34142
rect 37996 33506 38052 33516
rect 38332 34130 38500 34132
rect 38332 34078 38446 34130
rect 38498 34078 38500 34130
rect 38332 34076 38500 34078
rect 37324 33460 37380 33470
rect 37324 33366 37380 33404
rect 37660 33346 37716 33358
rect 37660 33294 37662 33346
rect 37714 33294 37716 33346
rect 37660 33236 37716 33294
rect 38332 33346 38388 34076
rect 38444 34066 38500 34076
rect 38332 33294 38334 33346
rect 38386 33294 38388 33346
rect 38332 33282 38388 33294
rect 38668 33348 38724 34190
rect 39004 34132 39060 34142
rect 38668 33282 38724 33292
rect 38780 33796 38836 33806
rect 38780 33346 38836 33740
rect 38780 33294 38782 33346
rect 38834 33294 38836 33346
rect 37996 33236 38052 33246
rect 37660 33234 38052 33236
rect 37660 33182 37998 33234
rect 38050 33182 38052 33234
rect 37660 33180 38052 33182
rect 37212 33030 37268 33068
rect 37436 33124 37492 33134
rect 37436 33030 37492 33068
rect 37100 32732 37380 32788
rect 37100 32562 37156 32574
rect 37100 32510 37102 32562
rect 37154 32510 37156 32562
rect 37100 32452 37156 32510
rect 36428 30156 36596 30212
rect 36988 32396 37100 32452
rect 36988 30212 37044 32396
rect 37100 32386 37156 32396
rect 37324 31890 37380 32732
rect 37772 32676 37828 33180
rect 37996 33170 38052 33180
rect 38108 33124 38164 33134
rect 38444 33124 38500 33134
rect 38164 33122 38500 33124
rect 38164 33070 38446 33122
rect 38498 33070 38500 33122
rect 38164 33068 38500 33070
rect 38108 33030 38164 33068
rect 38444 33058 38500 33068
rect 38668 33122 38724 33134
rect 38668 33070 38670 33122
rect 38722 33070 38724 33122
rect 38332 32900 38388 32910
rect 37772 32620 38164 32676
rect 37324 31838 37326 31890
rect 37378 31838 37380 31890
rect 37324 31826 37380 31838
rect 37884 32452 37940 32462
rect 37436 31554 37492 31566
rect 37436 31502 37438 31554
rect 37490 31502 37492 31554
rect 37436 31220 37492 31502
rect 37212 31164 37492 31220
rect 37548 31554 37604 31566
rect 37548 31502 37550 31554
rect 37602 31502 37604 31554
rect 37212 31106 37268 31164
rect 37212 31054 37214 31106
rect 37266 31054 37268 31106
rect 37212 31042 37268 31054
rect 37548 30548 37604 31502
rect 37548 30482 37604 30492
rect 37884 30994 37940 32396
rect 37996 31892 38052 31902
rect 37996 31778 38052 31836
rect 38108 31890 38164 32620
rect 38220 32452 38276 32462
rect 38220 32358 38276 32396
rect 38108 31838 38110 31890
rect 38162 31838 38164 31890
rect 38108 31826 38164 31838
rect 37996 31726 37998 31778
rect 38050 31726 38052 31778
rect 37996 31714 38052 31726
rect 38220 31556 38276 31566
rect 38220 31462 38276 31500
rect 38332 31332 38388 32844
rect 38556 32004 38612 32014
rect 38556 31778 38612 31948
rect 38556 31726 38558 31778
rect 38610 31726 38612 31778
rect 38556 31714 38612 31726
rect 38668 31892 38724 33070
rect 38668 31444 38724 31836
rect 38780 31556 38836 33294
rect 38780 31490 38836 31500
rect 39004 31554 39060 34076
rect 39116 33908 39172 35646
rect 39116 33842 39172 33852
rect 39004 31502 39006 31554
rect 39058 31502 39060 31554
rect 38668 31378 38724 31388
rect 37884 30942 37886 30994
rect 37938 30942 37940 30994
rect 36316 29426 36372 29438
rect 36316 29374 36318 29426
rect 36370 29374 36372 29426
rect 36316 28868 36372 29374
rect 36316 28802 36372 28812
rect 36428 28980 36484 30156
rect 36428 28754 36484 28924
rect 36428 28702 36430 28754
rect 36482 28702 36484 28754
rect 36428 28690 36484 28702
rect 36540 29986 36596 29998
rect 36540 29934 36542 29986
rect 36594 29934 36596 29986
rect 36540 28756 36596 29934
rect 36540 28690 36596 28700
rect 36764 29538 36820 29550
rect 36764 29486 36766 29538
rect 36818 29486 36820 29538
rect 36764 28420 36820 29486
rect 36988 29092 37044 30156
rect 37100 30436 37156 30446
rect 37100 30210 37156 30380
rect 37884 30436 37940 30942
rect 38220 31276 38388 31332
rect 38220 30996 38276 31276
rect 38556 31106 38612 31118
rect 38556 31054 38558 31106
rect 38610 31054 38612 31106
rect 38332 30996 38388 31006
rect 38220 30994 38388 30996
rect 38220 30942 38334 30994
rect 38386 30942 38388 30994
rect 38220 30940 38388 30942
rect 37884 30370 37940 30380
rect 37100 30158 37102 30210
rect 37154 30158 37156 30210
rect 37100 29092 37156 30158
rect 37324 30324 37380 30334
rect 37212 29428 37268 29438
rect 37324 29428 37380 30268
rect 37772 30100 37828 30110
rect 37436 30098 37828 30100
rect 37436 30046 37774 30098
rect 37826 30046 37828 30098
rect 37436 30044 37828 30046
rect 37436 29650 37492 30044
rect 37772 30034 37828 30044
rect 38332 29876 38388 30940
rect 38332 29810 38388 29820
rect 38444 30882 38500 30894
rect 38444 30830 38446 30882
rect 38498 30830 38500 30882
rect 38444 29652 38500 30830
rect 38556 30324 38612 31054
rect 38556 30258 38612 30268
rect 38892 30996 38948 31006
rect 39004 30996 39060 31502
rect 38892 30994 39060 30996
rect 38892 30942 38894 30994
rect 38946 30942 39060 30994
rect 38892 30940 39060 30942
rect 37436 29598 37438 29650
rect 37490 29598 37492 29650
rect 37436 29586 37492 29598
rect 37772 29596 38500 29652
rect 37772 29538 37828 29596
rect 37772 29486 37774 29538
rect 37826 29486 37828 29538
rect 37772 29474 37828 29486
rect 37436 29428 37492 29438
rect 37324 29426 37492 29428
rect 37324 29374 37438 29426
rect 37490 29374 37492 29426
rect 37324 29372 37492 29374
rect 37212 29334 37268 29372
rect 37436 29362 37492 29372
rect 38780 29426 38836 29438
rect 38780 29374 38782 29426
rect 38834 29374 38836 29426
rect 38108 29316 38164 29326
rect 38108 29314 38276 29316
rect 38108 29262 38110 29314
rect 38162 29262 38276 29314
rect 38108 29260 38276 29262
rect 38108 29250 38164 29260
rect 38108 29092 38164 29102
rect 37100 29036 37380 29092
rect 36988 29026 37044 29036
rect 36764 28354 36820 28364
rect 36876 28980 36932 28990
rect 36428 28196 36484 28206
rect 36484 28140 36820 28196
rect 36428 28130 36484 28140
rect 36764 27970 36820 28140
rect 36764 27918 36766 27970
rect 36818 27918 36820 27970
rect 36764 27906 36820 27918
rect 36428 26290 36484 26302
rect 36428 26238 36430 26290
rect 36482 26238 36484 26290
rect 36428 26180 36484 26238
rect 36428 26114 36484 26124
rect 34860 25396 34916 25406
rect 34860 24946 34916 25340
rect 35420 25396 35476 25406
rect 35420 25302 35476 25340
rect 35532 25394 35588 25406
rect 35532 25342 35534 25394
rect 35586 25342 35588 25394
rect 35196 25284 35252 25294
rect 35196 25190 35252 25228
rect 34860 24894 34862 24946
rect 34914 24894 34916 24946
rect 34748 24836 34804 24846
rect 34860 24836 34916 24894
rect 34804 24780 34916 24836
rect 34972 25172 35028 25182
rect 34748 24770 34804 24780
rect 34748 24612 34804 24622
rect 34748 24518 34804 24556
rect 34972 22594 35028 25116
rect 35532 25060 35588 25342
rect 35084 25004 35588 25060
rect 35084 24724 35140 25004
rect 35084 24630 35140 24668
rect 35868 24612 35924 24622
rect 35868 24518 35924 24556
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35868 23938 35924 23950
rect 35868 23886 35870 23938
rect 35922 23886 35924 23938
rect 35196 23828 35252 23838
rect 34972 22542 34974 22594
rect 35026 22542 35028 22594
rect 34972 22530 35028 22542
rect 35084 23826 35252 23828
rect 35084 23774 35198 23826
rect 35250 23774 35252 23826
rect 35084 23772 35252 23774
rect 35084 22482 35140 23772
rect 35196 23762 35252 23772
rect 35756 23716 35812 23726
rect 35756 23378 35812 23660
rect 35868 23604 35924 23886
rect 35868 23538 35924 23548
rect 35756 23326 35758 23378
rect 35810 23326 35812 23378
rect 35756 23314 35812 23326
rect 35308 23044 35364 23054
rect 35980 23044 36036 23054
rect 35308 23042 36036 23044
rect 35308 22990 35310 23042
rect 35362 22990 35982 23042
rect 36034 22990 36036 23042
rect 35308 22988 36036 22990
rect 35308 22978 35364 22988
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35084 22430 35086 22482
rect 35138 22430 35140 22482
rect 35084 22418 35140 22430
rect 35308 22372 35364 22382
rect 35532 22372 35588 22988
rect 35980 22978 36036 22988
rect 36092 22820 36148 25452
rect 36540 25284 36596 25294
rect 36540 25190 36596 25228
rect 35980 22764 36148 22820
rect 36204 23042 36260 23054
rect 36204 22990 36206 23042
rect 36258 22990 36260 23042
rect 35308 22370 35588 22372
rect 35308 22318 35310 22370
rect 35362 22318 35588 22370
rect 35308 22316 35588 22318
rect 35308 22306 35364 22316
rect 34860 21476 34916 21486
rect 34860 21382 34916 21420
rect 34636 21196 35140 21252
rect 34524 21140 34580 21150
rect 34188 20860 34356 20916
rect 33964 20750 33966 20802
rect 34018 20750 34020 20802
rect 33964 20738 34020 20750
rect 34188 20692 34244 20702
rect 34188 20598 34244 20636
rect 33964 20580 34020 20590
rect 33964 20132 34020 20524
rect 34076 20132 34132 20142
rect 33964 20076 34076 20132
rect 34076 20038 34132 20076
rect 33740 19964 34020 20020
rect 33628 18498 33684 18508
rect 33852 19348 33908 19358
rect 33852 19234 33908 19292
rect 33852 19182 33854 19234
rect 33906 19182 33908 19234
rect 33852 18452 33908 19182
rect 33740 18396 33852 18452
rect 33404 17554 33572 17556
rect 33404 17502 33406 17554
rect 33458 17502 33572 17554
rect 33404 17500 33572 17502
rect 33628 17556 33684 17566
rect 33404 17490 33460 17500
rect 33628 17462 33684 17500
rect 33180 17388 33348 17444
rect 33068 16996 33124 17006
rect 33068 16882 33124 16940
rect 33068 16830 33070 16882
rect 33122 16830 33124 16882
rect 33068 16818 33124 16830
rect 33068 16548 33124 16558
rect 33068 16210 33124 16492
rect 33068 16158 33070 16210
rect 33122 16158 33124 16210
rect 33068 16100 33124 16158
rect 33068 16034 33124 16044
rect 33180 15540 33236 15550
rect 33180 15446 33236 15484
rect 33292 15538 33348 17388
rect 33628 16100 33684 16110
rect 33740 16100 33796 18396
rect 33852 18358 33908 18396
rect 33852 17780 33908 17790
rect 33852 17666 33908 17724
rect 33852 17614 33854 17666
rect 33906 17614 33908 17666
rect 33852 17602 33908 17614
rect 33964 17444 34020 19964
rect 34300 19348 34356 20860
rect 34412 20468 34468 20478
rect 34412 20130 34468 20412
rect 34412 20078 34414 20130
rect 34466 20078 34468 20130
rect 34412 20066 34468 20078
rect 34524 20130 34580 21084
rect 34636 20690 34692 20702
rect 34636 20638 34638 20690
rect 34690 20638 34692 20690
rect 34636 20356 34692 20638
rect 34636 20290 34692 20300
rect 34524 20078 34526 20130
rect 34578 20078 34580 20130
rect 34524 20066 34580 20078
rect 34636 20130 34692 20142
rect 34636 20078 34638 20130
rect 34690 20078 34692 20130
rect 34636 19460 34692 20078
rect 34636 19394 34692 19404
rect 34300 19282 34356 19292
rect 34188 19122 34244 19134
rect 34188 19070 34190 19122
rect 34242 19070 34244 19122
rect 34188 18900 34244 19070
rect 34524 19122 34580 19134
rect 34524 19070 34526 19122
rect 34578 19070 34580 19122
rect 34524 19012 34580 19070
rect 34972 19124 35028 19134
rect 34972 19030 35028 19068
rect 34524 18946 34580 18956
rect 34860 19010 34916 19022
rect 34860 18958 34862 19010
rect 34914 18958 34916 19010
rect 34188 18834 34244 18844
rect 34860 18564 34916 18958
rect 34076 18508 34916 18564
rect 34076 17554 34132 18508
rect 34524 18340 34580 18350
rect 34524 18338 34692 18340
rect 34524 18286 34526 18338
rect 34578 18286 34692 18338
rect 34524 18284 34692 18286
rect 34524 18274 34580 18284
rect 34636 17778 34692 18284
rect 35084 18228 35140 21196
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35420 20802 35476 20814
rect 35420 20750 35422 20802
rect 35474 20750 35476 20802
rect 35420 20580 35476 20750
rect 35420 20514 35476 20524
rect 35308 20132 35364 20142
rect 35308 20038 35364 20076
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35420 19460 35476 19470
rect 35420 19346 35476 19404
rect 35420 19294 35422 19346
rect 35474 19294 35476 19346
rect 35420 19282 35476 19294
rect 34636 17726 34638 17778
rect 34690 17726 34692 17778
rect 34636 17714 34692 17726
rect 34860 18172 35140 18228
rect 34524 17668 34580 17678
rect 34076 17502 34078 17554
rect 34130 17502 34132 17554
rect 34076 17490 34132 17502
rect 34188 17556 34244 17566
rect 34188 17462 34244 17500
rect 33628 16098 33796 16100
rect 33628 16046 33630 16098
rect 33682 16046 33796 16098
rect 33628 16044 33796 16046
rect 33852 17388 34020 17444
rect 33628 16034 33684 16044
rect 33292 15486 33294 15538
rect 33346 15486 33348 15538
rect 33292 15474 33348 15486
rect 33628 15876 33684 15886
rect 33404 15428 33460 15438
rect 33404 15334 33460 15372
rect 32844 15138 32900 15148
rect 33628 14644 33684 15820
rect 33628 14550 33684 14588
rect 33852 14530 33908 17388
rect 34300 15988 34356 15998
rect 34300 15894 34356 15932
rect 33852 14478 33854 14530
rect 33906 14478 33908 14530
rect 33628 13972 33684 13982
rect 33852 13972 33908 14478
rect 33628 13970 33908 13972
rect 33628 13918 33630 13970
rect 33682 13918 33908 13970
rect 33628 13916 33908 13918
rect 33964 15314 34020 15326
rect 33964 15262 33966 15314
rect 34018 15262 34020 15314
rect 33964 13972 34020 15262
rect 34076 15202 34132 15214
rect 34076 15150 34078 15202
rect 34130 15150 34132 15202
rect 34076 14642 34132 15150
rect 34524 15148 34580 17612
rect 34860 15652 34916 18172
rect 35196 18060 35460 18070
rect 34972 18004 35028 18014
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35028 17948 35140 18004
rect 35196 17994 35460 18004
rect 34972 17938 35028 17948
rect 35084 17778 35140 17948
rect 35084 17726 35086 17778
rect 35138 17726 35140 17778
rect 35084 17714 35140 17726
rect 35420 16884 35476 16894
rect 35420 16770 35476 16828
rect 35420 16718 35422 16770
rect 35474 16718 35476 16770
rect 35420 16706 35476 16718
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 34860 15586 34916 15596
rect 35308 15988 35364 15998
rect 35308 15538 35364 15932
rect 35308 15486 35310 15538
rect 35362 15486 35364 15538
rect 35308 15474 35364 15486
rect 35420 15652 35476 15662
rect 35420 15538 35476 15596
rect 35420 15486 35422 15538
rect 35474 15486 35476 15538
rect 35420 15474 35476 15486
rect 34860 15316 34916 15326
rect 35196 15316 35252 15326
rect 34860 15314 35252 15316
rect 34860 15262 34862 15314
rect 34914 15262 35198 15314
rect 35250 15262 35252 15314
rect 34860 15260 35252 15262
rect 34860 15250 34916 15260
rect 35196 15250 35252 15260
rect 34076 14590 34078 14642
rect 34130 14590 34132 14642
rect 34076 14578 34132 14590
rect 34412 15092 34580 15148
rect 35532 15148 35588 22316
rect 35756 22370 35812 22382
rect 35756 22318 35758 22370
rect 35810 22318 35812 22370
rect 35756 22148 35812 22318
rect 35756 22082 35812 22092
rect 35644 19906 35700 19918
rect 35644 19854 35646 19906
rect 35698 19854 35700 19906
rect 35644 18788 35700 19854
rect 35868 19012 35924 19022
rect 35868 18918 35924 18956
rect 35980 18788 36036 22764
rect 36204 22708 36260 22990
rect 36652 23042 36708 23054
rect 36652 22990 36654 23042
rect 36706 22990 36708 23042
rect 36652 22930 36708 22990
rect 36876 23044 36932 28924
rect 37100 28644 37156 28654
rect 37100 28550 37156 28588
rect 36988 28532 37044 28542
rect 36988 28438 37044 28476
rect 37212 28420 37268 28458
rect 37212 28354 37268 28364
rect 37212 28196 37268 28206
rect 37212 27074 37268 28140
rect 37324 27860 37380 29036
rect 37436 28980 37492 28990
rect 37492 28924 37604 28980
rect 37436 28914 37492 28924
rect 37548 28868 37604 28924
rect 37548 28812 37716 28868
rect 37436 28756 37492 28766
rect 37492 28700 37604 28756
rect 37436 28690 37492 28700
rect 37436 27860 37492 27870
rect 37324 27858 37492 27860
rect 37324 27806 37438 27858
rect 37490 27806 37492 27858
rect 37324 27804 37492 27806
rect 37212 27022 37214 27074
rect 37266 27022 37268 27074
rect 37212 27010 37268 27022
rect 37436 27076 37492 27804
rect 37436 27010 37492 27020
rect 37548 26908 37604 28700
rect 37660 28642 37716 28812
rect 38108 28754 38164 29036
rect 38108 28702 38110 28754
rect 38162 28702 38164 28754
rect 38108 28690 38164 28702
rect 37660 28590 37662 28642
rect 37714 28590 37716 28642
rect 37660 28578 37716 28590
rect 38220 28420 38276 29260
rect 38780 29204 38836 29374
rect 38780 29138 38836 29148
rect 38556 28868 38612 28878
rect 38220 28354 38276 28364
rect 38444 28642 38500 28654
rect 38444 28590 38446 28642
rect 38498 28590 38500 28642
rect 38444 28196 38500 28590
rect 38444 28130 38500 28140
rect 37996 28084 38052 28094
rect 37996 28082 38276 28084
rect 37996 28030 37998 28082
rect 38050 28030 38276 28082
rect 37996 28028 38276 28030
rect 37996 28018 38052 28028
rect 38220 27972 38276 28028
rect 38556 28082 38612 28812
rect 38556 28030 38558 28082
rect 38610 28030 38612 28082
rect 38556 27972 38612 28030
rect 38220 27916 38612 27972
rect 38108 27858 38164 27870
rect 38108 27806 38110 27858
rect 38162 27806 38164 27858
rect 37996 27634 38052 27646
rect 37996 27582 37998 27634
rect 38050 27582 38052 27634
rect 37884 26962 37940 26974
rect 37884 26910 37886 26962
rect 37938 26910 37940 26962
rect 37884 26908 37940 26910
rect 37436 26852 37604 26908
rect 37660 26852 37940 26908
rect 37212 26628 37268 26638
rect 36988 26516 37044 26526
rect 36988 25508 37044 26460
rect 37212 26290 37268 26572
rect 37212 26238 37214 26290
rect 37266 26238 37268 26290
rect 37212 26226 37268 26238
rect 37436 25508 37492 26852
rect 37660 26514 37716 26852
rect 37660 26462 37662 26514
rect 37714 26462 37716 26514
rect 37660 26450 37716 26462
rect 37548 26402 37604 26414
rect 37548 26350 37550 26402
rect 37602 26350 37604 26402
rect 37548 26180 37604 26350
rect 37772 26404 37828 26414
rect 37996 26404 38052 27582
rect 38108 26628 38164 27806
rect 38892 26908 38948 30940
rect 39228 28868 39284 35868
rect 39340 35830 39396 35868
rect 39900 35812 39956 35822
rect 40124 35812 40180 36206
rect 39900 35810 40124 35812
rect 39900 35758 39902 35810
rect 39954 35758 40124 35810
rect 39900 35756 40124 35758
rect 39900 35746 39956 35756
rect 40124 35746 40180 35756
rect 40348 36260 40404 36876
rect 40348 35586 40404 36204
rect 40348 35534 40350 35586
rect 40402 35534 40404 35586
rect 40348 35252 40404 35534
rect 40348 35186 40404 35196
rect 39676 34132 39732 34142
rect 39676 34038 39732 34076
rect 40012 34130 40068 34142
rect 40012 34078 40014 34130
rect 40066 34078 40068 34130
rect 39340 33348 39396 33358
rect 39340 32452 39396 33292
rect 39340 32386 39396 32396
rect 40012 32564 40068 34078
rect 40236 34130 40292 34142
rect 40236 34078 40238 34130
rect 40290 34078 40292 34130
rect 40124 34018 40180 34030
rect 40124 33966 40126 34018
rect 40178 33966 40180 34018
rect 40124 33908 40180 33966
rect 40236 34020 40292 34078
rect 40236 33964 40404 34020
rect 40124 33852 40292 33908
rect 40124 33684 40180 33694
rect 40124 33458 40180 33628
rect 40124 33406 40126 33458
rect 40178 33406 40180 33458
rect 40124 33394 40180 33406
rect 40236 32676 40292 33852
rect 40236 32610 40292 32620
rect 40348 32788 40404 33964
rect 40012 32004 40068 32508
rect 40236 32452 40292 32462
rect 40012 31938 40068 31948
rect 40124 32450 40292 32452
rect 40124 32398 40238 32450
rect 40290 32398 40292 32450
rect 40124 32396 40292 32398
rect 39340 31892 39396 31902
rect 39396 31836 39620 31892
rect 39340 31798 39396 31836
rect 39340 31556 39396 31566
rect 39340 30994 39396 31500
rect 39340 30942 39342 30994
rect 39394 30942 39396 30994
rect 39340 30930 39396 30942
rect 39564 30994 39620 31836
rect 39564 30942 39566 30994
rect 39618 30942 39620 30994
rect 39564 30930 39620 30942
rect 40124 30436 40180 32396
rect 40236 32386 40292 32396
rect 40348 32228 40404 32732
rect 40460 32452 40516 37772
rect 40572 36596 40628 42588
rect 40908 41860 40964 41870
rect 40684 41186 40740 41198
rect 40684 41134 40686 41186
rect 40738 41134 40740 41186
rect 40684 40628 40740 41134
rect 40684 40562 40740 40572
rect 40796 40962 40852 40974
rect 40796 40910 40798 40962
rect 40850 40910 40852 40962
rect 40796 38948 40852 40910
rect 40796 38882 40852 38892
rect 40908 38946 40964 41804
rect 41020 40404 41076 42812
rect 41356 42802 41412 42812
rect 41804 42644 41860 42654
rect 41580 42642 41860 42644
rect 41580 42590 41806 42642
rect 41858 42590 41860 42642
rect 41580 42588 41860 42590
rect 41468 42082 41524 42094
rect 41468 42030 41470 42082
rect 41522 42030 41524 42082
rect 41132 41972 41188 41982
rect 41132 41878 41188 41916
rect 41468 41972 41524 42030
rect 41468 41906 41524 41916
rect 41132 41074 41188 41086
rect 41132 41022 41134 41074
rect 41186 41022 41188 41074
rect 41132 40852 41188 41022
rect 41132 40786 41188 40796
rect 41468 40962 41524 40974
rect 41468 40910 41470 40962
rect 41522 40910 41524 40962
rect 41468 40404 41524 40910
rect 41020 40402 41300 40404
rect 41020 40350 41022 40402
rect 41074 40350 41300 40402
rect 41020 40348 41300 40350
rect 41020 40338 41076 40348
rect 41132 39620 41188 39630
rect 41244 39620 41300 40348
rect 41468 40338 41524 40348
rect 41580 40180 41636 42588
rect 41804 42578 41860 42588
rect 41804 41860 41860 41870
rect 41804 41766 41860 41804
rect 41692 41748 41748 41758
rect 41692 40514 41748 41692
rect 41692 40462 41694 40514
rect 41746 40462 41748 40514
rect 41692 40450 41748 40462
rect 41804 41188 41860 41198
rect 41132 39618 41300 39620
rect 41132 39566 41134 39618
rect 41186 39566 41300 39618
rect 41132 39564 41300 39566
rect 41468 40124 41636 40180
rect 41020 39060 41076 39070
rect 41020 38966 41076 39004
rect 40908 38894 40910 38946
rect 40962 38894 40964 38946
rect 40908 38882 40964 38894
rect 41132 38050 41188 39564
rect 41468 39060 41524 40124
rect 41580 39956 41636 39966
rect 41580 39618 41636 39900
rect 41580 39566 41582 39618
rect 41634 39566 41636 39618
rect 41580 39554 41636 39566
rect 41692 39620 41748 39630
rect 41804 39620 41860 41132
rect 41692 39618 41860 39620
rect 41692 39566 41694 39618
rect 41746 39566 41860 39618
rect 41692 39564 41860 39566
rect 41468 38994 41524 39004
rect 41580 38724 41636 38734
rect 41692 38724 41748 39564
rect 41916 39284 41972 44940
rect 42140 44210 42196 44222
rect 42140 44158 42142 44210
rect 42194 44158 42196 44210
rect 42140 42196 42196 44158
rect 42140 42130 42196 42140
rect 42140 41970 42196 41982
rect 42140 41918 42142 41970
rect 42194 41918 42196 41970
rect 42140 39732 42196 41918
rect 42364 40404 42420 45838
rect 42700 45778 42756 45790
rect 42700 45726 42702 45778
rect 42754 45726 42756 45778
rect 42700 43540 42756 45726
rect 42812 45668 42868 45678
rect 42812 45574 42868 45612
rect 42924 45666 42980 45678
rect 42924 45614 42926 45666
rect 42978 45614 42980 45666
rect 42924 43876 42980 45614
rect 43036 44548 43092 46732
rect 44380 46004 44436 49200
rect 44604 46116 44660 46126
rect 44604 46022 44660 46060
rect 44380 45948 44548 46004
rect 43932 45890 43988 45902
rect 43932 45838 43934 45890
rect 43986 45838 43988 45890
rect 43260 45556 43316 45566
rect 43148 44548 43204 44558
rect 43036 44492 43148 44548
rect 43148 44482 43204 44492
rect 43036 43876 43092 43886
rect 42924 43820 43036 43876
rect 43036 43810 43092 43820
rect 43260 43652 43316 45500
rect 43148 43596 43316 43652
rect 43820 44994 43876 45006
rect 43820 44942 43822 44994
rect 43874 44942 43876 44994
rect 42700 43474 42756 43484
rect 43036 43538 43092 43550
rect 43036 43486 43038 43538
rect 43090 43486 43092 43538
rect 42476 42868 42532 42878
rect 42476 42754 42532 42812
rect 42476 42702 42478 42754
rect 42530 42702 42532 42754
rect 42476 42690 42532 42702
rect 43036 42084 43092 43486
rect 43148 42642 43204 43596
rect 43260 43428 43316 43438
rect 43260 42866 43316 43372
rect 43260 42814 43262 42866
rect 43314 42814 43316 42866
rect 43260 42802 43316 42814
rect 43708 42868 43764 42906
rect 43708 42802 43764 42812
rect 43148 42590 43150 42642
rect 43202 42590 43204 42642
rect 43148 42532 43204 42590
rect 43372 42644 43428 42654
rect 43372 42642 43652 42644
rect 43372 42590 43374 42642
rect 43426 42590 43652 42642
rect 43372 42588 43652 42590
rect 43372 42578 43428 42588
rect 43148 42466 43204 42476
rect 43372 42084 43428 42094
rect 43036 42082 43428 42084
rect 43036 42030 43374 42082
rect 43426 42030 43428 42082
rect 43036 42028 43428 42030
rect 42588 41972 42644 41982
rect 42476 41188 42532 41198
rect 42476 41094 42532 41132
rect 42588 40852 42644 41916
rect 42364 40348 42532 40404
rect 42028 39676 42196 39732
rect 42364 40180 42420 40190
rect 42028 39618 42084 39676
rect 42028 39566 42030 39618
rect 42082 39566 42084 39618
rect 42028 39508 42084 39566
rect 42028 39442 42084 39452
rect 42252 39618 42308 39630
rect 42252 39566 42254 39618
rect 42306 39566 42308 39618
rect 42252 39284 42308 39566
rect 42364 39396 42420 40124
rect 42476 39956 42532 40348
rect 42476 39890 42532 39900
rect 42476 39732 42532 39742
rect 42588 39732 42644 40796
rect 42476 39730 42644 39732
rect 42476 39678 42478 39730
rect 42530 39678 42644 39730
rect 42476 39676 42644 39678
rect 42700 41970 42756 41982
rect 42700 41918 42702 41970
rect 42754 41918 42756 41970
rect 42700 40292 42756 41918
rect 42924 41970 42980 41982
rect 42924 41918 42926 41970
rect 42978 41918 42980 41970
rect 42700 39730 42756 40236
rect 42700 39678 42702 39730
rect 42754 39678 42756 39730
rect 42476 39666 42532 39676
rect 42700 39666 42756 39678
rect 42812 41748 42868 41758
rect 42812 41186 42868 41692
rect 42924 41300 42980 41918
rect 43372 41972 43428 42028
rect 43372 41906 43428 41916
rect 43484 42084 43540 42094
rect 42924 41234 42980 41244
rect 42812 41134 42814 41186
rect 42866 41134 42868 41186
rect 42812 39620 42868 41134
rect 43484 41186 43540 42028
rect 43484 41134 43486 41186
rect 43538 41134 43540 41186
rect 43372 40628 43428 40638
rect 43036 39620 43092 39630
rect 43372 39620 43428 40572
rect 43484 40516 43540 41134
rect 43484 40450 43540 40460
rect 42812 39618 43092 39620
rect 42812 39566 43038 39618
rect 43090 39566 43092 39618
rect 42812 39564 43092 39566
rect 43036 39554 43092 39564
rect 43148 39618 43428 39620
rect 43148 39566 43374 39618
rect 43426 39566 43428 39618
rect 43148 39564 43428 39566
rect 42588 39508 42644 39518
rect 42476 39396 42532 39406
rect 42364 39394 42532 39396
rect 42364 39342 42478 39394
rect 42530 39342 42532 39394
rect 42364 39340 42532 39342
rect 42476 39330 42532 39340
rect 41916 39228 42196 39284
rect 42028 39060 42084 39070
rect 42140 39060 42196 39228
rect 42252 39218 42308 39228
rect 42364 39060 42420 39070
rect 42140 39058 42420 39060
rect 42140 39006 42366 39058
rect 42418 39006 42420 39058
rect 42140 39004 42420 39006
rect 42028 38966 42084 39004
rect 42364 38994 42420 39004
rect 42476 38948 42532 38958
rect 42476 38854 42532 38892
rect 41580 38722 41748 38724
rect 41580 38670 41582 38722
rect 41634 38670 41748 38722
rect 41580 38668 41748 38670
rect 42588 38836 42644 39452
rect 43148 39396 43204 39564
rect 43372 39554 43428 39564
rect 42588 38668 42644 38780
rect 42924 39340 43204 39396
rect 43260 39394 43316 39406
rect 43260 39342 43262 39394
rect 43314 39342 43316 39394
rect 41580 38658 41636 38668
rect 42588 38612 42756 38668
rect 41132 37998 41134 38050
rect 41186 37998 41188 38050
rect 40684 37938 40740 37950
rect 40684 37886 40686 37938
rect 40738 37886 40740 37938
rect 40684 37604 40740 37886
rect 40796 37940 40852 37950
rect 40796 37846 40852 37884
rect 41132 37828 41188 37998
rect 41916 37940 41972 37950
rect 41916 37846 41972 37884
rect 41804 37828 41860 37838
rect 41132 37762 41188 37772
rect 41692 37772 41804 37828
rect 40684 37548 41076 37604
rect 41020 37490 41076 37548
rect 41020 37438 41022 37490
rect 41074 37438 41076 37490
rect 41020 37426 41076 37438
rect 41132 37380 41188 37390
rect 41132 37286 41188 37324
rect 41692 37266 41748 37772
rect 41804 37762 41860 37772
rect 41692 37214 41694 37266
rect 41746 37214 41748 37266
rect 40796 36596 40852 36606
rect 40572 36594 40852 36596
rect 40572 36542 40798 36594
rect 40850 36542 40852 36594
rect 40572 36540 40852 36542
rect 40796 36530 40852 36540
rect 41580 36482 41636 36494
rect 41580 36430 41582 36482
rect 41634 36430 41636 36482
rect 41132 36258 41188 36270
rect 41132 36206 41134 36258
rect 41186 36206 41188 36258
rect 41132 36148 41188 36206
rect 41132 36082 41188 36092
rect 41244 36258 41300 36270
rect 41244 36206 41246 36258
rect 41298 36206 41300 36258
rect 41244 35812 41300 36206
rect 41356 36258 41412 36270
rect 41356 36206 41358 36258
rect 41410 36206 41412 36258
rect 41356 36036 41412 36206
rect 41468 36260 41524 36270
rect 41468 36166 41524 36204
rect 41356 35970 41412 35980
rect 41244 35756 41412 35812
rect 41244 35588 41300 35598
rect 41244 35494 41300 35532
rect 41356 35364 41412 35756
rect 41468 35698 41524 35710
rect 41468 35646 41470 35698
rect 41522 35646 41524 35698
rect 41468 35364 41524 35646
rect 40908 35308 41524 35364
rect 40796 35028 40852 35038
rect 40908 35028 40964 35308
rect 41580 35252 41636 36430
rect 41692 35924 41748 37214
rect 41916 37266 41972 37278
rect 41916 37214 41918 37266
rect 41970 37214 41972 37266
rect 41916 37156 41972 37214
rect 42700 37266 42756 38612
rect 42700 37214 42702 37266
rect 42754 37214 42756 37266
rect 42700 37156 42756 37214
rect 41972 37100 42308 37156
rect 41916 37090 41972 37100
rect 42140 36484 42196 36494
rect 42140 36148 42196 36428
rect 42252 36482 42308 37100
rect 42700 37090 42756 37100
rect 42252 36430 42254 36482
rect 42306 36430 42308 36482
rect 42252 36418 42308 36430
rect 42364 36372 42420 36382
rect 42364 36278 42420 36316
rect 42700 36370 42756 36382
rect 42700 36318 42702 36370
rect 42754 36318 42756 36370
rect 42476 36260 42532 36270
rect 42476 36166 42532 36204
rect 42196 36092 42308 36148
rect 42140 36082 42196 36092
rect 41692 35868 42196 35924
rect 41692 35700 41748 35710
rect 41692 35606 41748 35644
rect 41804 35698 41860 35710
rect 41804 35646 41806 35698
rect 41858 35646 41860 35698
rect 41356 35196 41636 35252
rect 41244 35028 41300 35038
rect 40796 35026 40964 35028
rect 40796 34974 40798 35026
rect 40850 34974 40964 35026
rect 40796 34972 40964 34974
rect 41020 35026 41300 35028
rect 41020 34974 41246 35026
rect 41298 34974 41300 35026
rect 41020 34972 41300 34974
rect 40796 34962 40852 34972
rect 41020 34242 41076 34972
rect 41244 34962 41300 34972
rect 41020 34190 41022 34242
rect 41074 34190 41076 34242
rect 41020 34178 41076 34190
rect 41244 34690 41300 34702
rect 41244 34638 41246 34690
rect 41298 34638 41300 34690
rect 40908 33906 40964 33918
rect 40908 33854 40910 33906
rect 40962 33854 40964 33906
rect 40908 33684 40964 33854
rect 41244 33906 41300 34638
rect 41244 33854 41246 33906
rect 41298 33854 41300 33906
rect 41244 33842 41300 33854
rect 41356 34690 41412 35196
rect 41804 35140 41860 35646
rect 41692 35084 41860 35140
rect 41356 34638 41358 34690
rect 41410 34638 41412 34690
rect 40908 33618 40964 33628
rect 41356 33460 41412 34638
rect 41580 34690 41636 34702
rect 41580 34638 41582 34690
rect 41634 34638 41636 34690
rect 41468 34132 41524 34142
rect 41468 34038 41524 34076
rect 41356 33394 41412 33404
rect 41580 32900 41636 34638
rect 41692 33796 41748 35084
rect 41804 34916 41860 34926
rect 41916 34916 41972 35868
rect 42140 35810 42196 35868
rect 42140 35758 42142 35810
rect 42194 35758 42196 35810
rect 42140 35746 42196 35758
rect 41804 34914 41916 34916
rect 41804 34862 41806 34914
rect 41858 34862 41916 34914
rect 41804 34860 41916 34862
rect 41804 34850 41860 34860
rect 41916 34822 41972 34860
rect 42252 34468 42308 36092
rect 42476 36036 42532 36046
rect 42476 35698 42532 35980
rect 42476 35646 42478 35698
rect 42530 35646 42532 35698
rect 42476 35634 42532 35646
rect 42588 35586 42644 35598
rect 42588 35534 42590 35586
rect 42642 35534 42644 35586
rect 42476 35028 42532 35038
rect 42588 35028 42644 35534
rect 42476 35026 42644 35028
rect 42476 34974 42478 35026
rect 42530 34974 42644 35026
rect 42476 34972 42644 34974
rect 42700 35586 42756 36318
rect 42700 35534 42702 35586
rect 42754 35534 42756 35586
rect 42476 34962 42532 34972
rect 42588 34692 42644 34702
rect 42588 34598 42644 34636
rect 42028 34412 42308 34468
rect 42028 34354 42084 34412
rect 42028 34302 42030 34354
rect 42082 34302 42084 34354
rect 42028 33906 42084 34302
rect 42252 34020 42308 34030
rect 42700 34020 42756 35534
rect 42252 34018 42756 34020
rect 42252 33966 42254 34018
rect 42306 33966 42756 34018
rect 42252 33964 42756 33966
rect 42812 35924 42868 35934
rect 42252 33954 42308 33964
rect 42028 33854 42030 33906
rect 42082 33854 42084 33906
rect 42028 33842 42084 33854
rect 41692 33730 41748 33740
rect 42252 33460 42308 33470
rect 42252 33366 42308 33404
rect 41580 32834 41636 32844
rect 41916 33012 41972 33022
rect 41468 32788 41524 32798
rect 40908 32676 40964 32686
rect 40908 32582 40964 32620
rect 41468 32674 41524 32732
rect 41468 32622 41470 32674
rect 41522 32622 41524 32674
rect 41468 32610 41524 32622
rect 41132 32564 41188 32574
rect 40572 32452 40628 32462
rect 40460 32396 40572 32452
rect 40236 32172 40404 32228
rect 40236 31106 40292 32172
rect 40348 31220 40404 31230
rect 40404 31164 40516 31220
rect 40348 31154 40404 31164
rect 40236 31054 40238 31106
rect 40290 31054 40292 31106
rect 40236 31042 40292 31054
rect 39788 30324 39844 30334
rect 39900 30324 39956 30334
rect 39844 30322 39956 30324
rect 39844 30270 39902 30322
rect 39954 30270 39956 30322
rect 39844 30268 39956 30270
rect 39228 28802 39284 28812
rect 39564 29428 39620 29438
rect 39228 28532 39284 28542
rect 39116 28530 39284 28532
rect 39116 28478 39230 28530
rect 39282 28478 39284 28530
rect 39116 28476 39284 28478
rect 39004 28420 39060 28430
rect 39004 27970 39060 28364
rect 39116 28082 39172 28476
rect 39228 28466 39284 28476
rect 39116 28030 39118 28082
rect 39170 28030 39172 28082
rect 39116 28018 39172 28030
rect 39340 28084 39396 28094
rect 39004 27918 39006 27970
rect 39058 27918 39060 27970
rect 39004 27906 39060 27918
rect 39340 27860 39396 28028
rect 39564 28082 39620 29372
rect 39564 28030 39566 28082
rect 39618 28030 39620 28082
rect 39564 28018 39620 28030
rect 39788 28082 39844 30268
rect 39900 30258 39956 30268
rect 39788 28030 39790 28082
rect 39842 28030 39844 28082
rect 39788 28018 39844 28030
rect 39900 29876 39956 29886
rect 39900 27970 39956 29820
rect 40012 29540 40068 29550
rect 40012 29446 40068 29484
rect 40124 28084 40180 30380
rect 40236 29428 40292 29438
rect 40236 29314 40292 29372
rect 40236 29262 40238 29314
rect 40290 29262 40292 29314
rect 40236 29250 40292 29262
rect 40460 28868 40516 31164
rect 40348 28084 40404 28094
rect 40180 28082 40404 28084
rect 40180 28030 40350 28082
rect 40402 28030 40404 28082
rect 40180 28028 40404 28030
rect 40124 27990 40180 28028
rect 40348 28018 40404 28028
rect 39900 27918 39902 27970
rect 39954 27918 39956 27970
rect 39900 27906 39956 27918
rect 38108 26562 38164 26572
rect 38780 26852 38948 26908
rect 39116 27858 39396 27860
rect 39116 27806 39342 27858
rect 39394 27806 39396 27858
rect 39116 27804 39396 27806
rect 38668 26516 38724 26526
rect 38668 26422 38724 26460
rect 37772 26402 38052 26404
rect 37772 26350 37774 26402
rect 37826 26350 38052 26402
rect 37772 26348 38052 26350
rect 38220 26404 38276 26414
rect 37772 26338 37828 26348
rect 38108 26180 38164 26190
rect 37548 26178 38164 26180
rect 37548 26126 38110 26178
rect 38162 26126 38164 26178
rect 37548 26124 38164 26126
rect 38108 26114 38164 26124
rect 37548 25508 37604 25518
rect 36988 25506 37380 25508
rect 36988 25454 36990 25506
rect 37042 25454 37380 25506
rect 36988 25452 37380 25454
rect 37436 25452 37548 25508
rect 36988 25442 37044 25452
rect 37100 25282 37156 25294
rect 37100 25230 37102 25282
rect 37154 25230 37156 25282
rect 37100 25172 37156 25230
rect 37100 25106 37156 25116
rect 37212 25282 37268 25294
rect 37212 25230 37214 25282
rect 37266 25230 37268 25282
rect 37212 24724 37268 25230
rect 36988 24668 37268 24724
rect 36988 24612 37044 24668
rect 36988 24050 37044 24556
rect 37212 24164 37268 24174
rect 37324 24164 37380 25452
rect 37548 25442 37604 25452
rect 37212 24162 37380 24164
rect 37212 24110 37214 24162
rect 37266 24110 37380 24162
rect 37212 24108 37380 24110
rect 37436 25284 37492 25294
rect 37212 24098 37268 24108
rect 36988 23998 36990 24050
rect 37042 23998 37044 24050
rect 36988 23986 37044 23998
rect 37100 23044 37156 23054
rect 36876 23042 37156 23044
rect 36876 22990 37102 23042
rect 37154 22990 37156 23042
rect 36876 22988 37156 22990
rect 36652 22878 36654 22930
rect 36706 22878 36708 22930
rect 36652 22866 36708 22878
rect 36092 22652 36260 22708
rect 36092 22036 36148 22652
rect 36092 21970 36148 21980
rect 36204 22146 36260 22158
rect 36204 22094 36206 22146
rect 36258 22094 36260 22146
rect 36204 21588 36260 22094
rect 36316 22146 36372 22158
rect 36316 22094 36318 22146
rect 36370 22094 36372 22146
rect 36316 21700 36372 22094
rect 36428 22146 36484 22158
rect 36428 22094 36430 22146
rect 36482 22094 36484 22146
rect 36428 21812 36484 22094
rect 36988 22148 37044 22988
rect 37100 22978 37156 22988
rect 37212 22484 37268 22494
rect 36988 22082 37044 22092
rect 37100 22482 37268 22484
rect 37100 22430 37214 22482
rect 37266 22430 37268 22482
rect 37100 22428 37268 22430
rect 36428 21746 36484 21756
rect 36316 21634 36372 21644
rect 36204 21522 36260 21532
rect 36988 21474 37044 21486
rect 36988 21422 36990 21474
rect 37042 21422 37044 21474
rect 36316 20804 36372 20814
rect 36316 20710 36372 20748
rect 36988 20804 37044 21422
rect 36988 20710 37044 20748
rect 37100 20580 37156 22428
rect 37212 22418 37268 22428
rect 37436 22260 37492 25228
rect 37772 25172 37828 25182
rect 37828 25116 37940 25172
rect 37772 25106 37828 25116
rect 37884 24162 37940 25116
rect 37884 24110 37886 24162
rect 37938 24110 37940 24162
rect 37884 24098 37940 24110
rect 37996 24610 38052 24622
rect 37996 24558 37998 24610
rect 38050 24558 38052 24610
rect 37996 24050 38052 24558
rect 37996 23998 37998 24050
rect 38050 23998 38052 24050
rect 37996 23986 38052 23998
rect 38220 23940 38276 26348
rect 38444 26292 38500 26302
rect 38444 26198 38500 26236
rect 38780 24948 38836 26852
rect 38892 26404 38948 26414
rect 38892 26310 38948 26348
rect 39004 26292 39060 26302
rect 39004 26198 39060 26236
rect 38108 23938 38276 23940
rect 38108 23886 38222 23938
rect 38274 23886 38276 23938
rect 38108 23884 38276 23886
rect 37548 23828 37604 23838
rect 38108 23828 38164 23884
rect 38220 23874 38276 23884
rect 38668 24892 38836 24948
rect 39116 24948 39172 27804
rect 39340 27794 39396 27804
rect 40012 27186 40068 27198
rect 40012 27134 40014 27186
rect 40066 27134 40068 27186
rect 40012 26908 40068 27134
rect 40460 27186 40516 28812
rect 40460 27134 40462 27186
rect 40514 27134 40516 27186
rect 40460 27122 40516 27134
rect 39564 26852 40068 26908
rect 39564 26402 39620 26852
rect 39564 26350 39566 26402
rect 39618 26350 39620 26402
rect 39564 26338 39620 26350
rect 39452 26180 39508 26190
rect 39452 26086 39508 26124
rect 40012 26180 40068 26190
rect 40012 25732 40068 26124
rect 39228 25620 39284 25630
rect 39228 25526 39284 25564
rect 39788 25284 39844 25294
rect 39788 25190 39844 25228
rect 37548 23826 38164 23828
rect 37548 23774 37550 23826
rect 37602 23774 38164 23826
rect 37548 23772 38164 23774
rect 37548 23762 37604 23772
rect 38668 23716 38724 24892
rect 38780 24724 38836 24734
rect 38780 24630 38836 24668
rect 39116 24722 39172 24892
rect 39116 24670 39118 24722
rect 39170 24670 39172 24722
rect 39116 24658 39172 24670
rect 39676 24722 39732 24734
rect 39676 24670 39678 24722
rect 39730 24670 39732 24722
rect 38556 23660 38724 23716
rect 39676 23716 39732 24670
rect 38556 23492 38612 23660
rect 39676 23650 39732 23660
rect 40012 24724 40068 25676
rect 40236 25506 40292 25518
rect 40236 25454 40238 25506
rect 40290 25454 40292 25506
rect 40236 25284 40292 25454
rect 40236 25218 40292 25228
rect 40460 25282 40516 25294
rect 40460 25230 40462 25282
rect 40514 25230 40516 25282
rect 40460 25060 40516 25230
rect 40236 25004 40516 25060
rect 40236 24724 40292 25004
rect 40348 24836 40404 24846
rect 40348 24742 40404 24780
rect 40012 24722 40292 24724
rect 40012 24670 40014 24722
rect 40066 24670 40292 24722
rect 40012 24668 40292 24670
rect 40572 24724 40628 32396
rect 41020 30772 41076 30782
rect 40796 30212 40852 30222
rect 40796 30118 40852 30156
rect 41020 29316 41076 30716
rect 41132 29538 41188 32508
rect 41356 32450 41412 32462
rect 41356 32398 41358 32450
rect 41410 32398 41412 32450
rect 41356 31892 41412 32398
rect 41916 32450 41972 32956
rect 41916 32398 41918 32450
rect 41970 32398 41972 32450
rect 41916 32386 41972 32398
rect 41468 31892 41524 31902
rect 41356 31890 41524 31892
rect 41356 31838 41470 31890
rect 41522 31838 41524 31890
rect 41356 31836 41524 31838
rect 41468 31826 41524 31836
rect 42252 31892 42308 31902
rect 42252 31778 42308 31836
rect 42252 31726 42254 31778
rect 42306 31726 42308 31778
rect 41580 31556 41636 31566
rect 41468 30996 41524 31006
rect 41580 30996 41636 31500
rect 41468 30994 41636 30996
rect 41468 30942 41470 30994
rect 41522 30942 41636 30994
rect 41468 30940 41636 30942
rect 41468 30212 41524 30940
rect 41468 30146 41524 30156
rect 42252 30322 42308 31726
rect 42252 30270 42254 30322
rect 42306 30270 42308 30322
rect 41132 29486 41134 29538
rect 41186 29486 41188 29538
rect 41132 29474 41188 29486
rect 41356 29540 41412 29550
rect 42252 29540 42308 30270
rect 41244 29428 41300 29438
rect 41244 29334 41300 29372
rect 41020 29260 41188 29316
rect 41020 28084 41076 28094
rect 41020 27990 41076 28028
rect 40796 27074 40852 27086
rect 40796 27022 40798 27074
rect 40850 27022 40852 27074
rect 40796 26180 40852 27022
rect 40796 26114 40852 26124
rect 41020 26180 41076 26190
rect 40908 25506 40964 25518
rect 40908 25454 40910 25506
rect 40962 25454 40964 25506
rect 40908 25284 40964 25454
rect 40908 25218 40964 25228
rect 40908 24724 40964 24734
rect 40572 24722 40964 24724
rect 40572 24670 40910 24722
rect 40962 24670 40964 24722
rect 40572 24668 40964 24670
rect 40012 23604 40068 24668
rect 40908 24658 40964 24668
rect 40572 24052 40628 24062
rect 41020 24052 41076 26124
rect 40348 24050 41076 24052
rect 40348 23998 40574 24050
rect 40626 23998 41076 24050
rect 40348 23996 41076 23998
rect 41132 25282 41188 29260
rect 41132 25230 41134 25282
rect 41186 25230 41188 25282
rect 40124 23716 40180 23726
rect 40124 23622 40180 23660
rect 40012 23538 40068 23548
rect 38556 23426 38612 23436
rect 38108 23268 38164 23278
rect 37436 22194 37492 22204
rect 37996 23266 38164 23268
rect 37996 23214 38110 23266
rect 38162 23214 38164 23266
rect 37996 23212 38164 23214
rect 37100 20514 37156 20524
rect 37212 21812 37268 21822
rect 36092 20132 36148 20142
rect 36092 20038 36148 20076
rect 37212 20018 37268 21756
rect 37884 21812 37940 21822
rect 37324 21700 37380 21710
rect 37324 21606 37380 21644
rect 37660 21700 37716 21710
rect 37660 21586 37716 21644
rect 37884 21698 37940 21756
rect 37884 21646 37886 21698
rect 37938 21646 37940 21698
rect 37884 21634 37940 21646
rect 37660 21534 37662 21586
rect 37714 21534 37716 21586
rect 37660 21364 37716 21534
rect 37772 21476 37828 21486
rect 37772 21382 37828 21420
rect 37324 21308 37716 21364
rect 37324 20690 37380 21308
rect 37324 20638 37326 20690
rect 37378 20638 37380 20690
rect 37324 20626 37380 20638
rect 37884 20692 37940 20702
rect 37996 20692 38052 23212
rect 38108 23202 38164 23212
rect 38220 23156 38276 23166
rect 38108 21700 38164 21710
rect 38108 20802 38164 21644
rect 38220 20916 38276 23100
rect 38332 23154 38388 23166
rect 38332 23102 38334 23154
rect 38386 23102 38388 23154
rect 38332 21700 38388 23102
rect 38556 23154 38612 23166
rect 38556 23102 38558 23154
rect 38610 23102 38612 23154
rect 38444 23044 38500 23054
rect 38444 22950 38500 22988
rect 38332 21634 38388 21644
rect 38444 21812 38500 21822
rect 38332 20916 38388 20926
rect 38220 20914 38388 20916
rect 38220 20862 38334 20914
rect 38386 20862 38388 20914
rect 38220 20860 38388 20862
rect 38332 20850 38388 20860
rect 38108 20750 38110 20802
rect 38162 20750 38164 20802
rect 38108 20738 38164 20750
rect 38444 20802 38500 21756
rect 38444 20750 38446 20802
rect 38498 20750 38500 20802
rect 37884 20690 38052 20692
rect 37884 20638 37886 20690
rect 37938 20638 38052 20690
rect 37884 20636 38052 20638
rect 37884 20580 37940 20636
rect 37884 20514 37940 20524
rect 38444 20356 38500 20750
rect 38444 20290 38500 20300
rect 38444 20132 38500 20142
rect 38556 20132 38612 23102
rect 38892 23156 38948 23194
rect 38892 23090 38948 23100
rect 39004 23044 39060 23054
rect 39004 22260 39060 22988
rect 39116 23042 39172 23054
rect 39116 22990 39118 23042
rect 39170 22990 39172 23042
rect 39116 22484 39172 22990
rect 39228 22932 39284 22942
rect 39228 22838 39284 22876
rect 39340 22484 39396 22494
rect 39116 22482 39396 22484
rect 39116 22430 39342 22482
rect 39394 22430 39396 22482
rect 39116 22428 39396 22430
rect 39340 22418 39396 22428
rect 39004 21474 39060 22204
rect 40124 22370 40180 22382
rect 40124 22318 40126 22370
rect 40178 22318 40180 22370
rect 40124 21924 40180 22318
rect 40348 22036 40404 23996
rect 40572 23986 40628 23996
rect 41132 23940 41188 25230
rect 41244 28756 41300 28766
rect 41244 25172 41300 28700
rect 41356 28754 41412 29484
rect 42028 29484 42252 29540
rect 41916 29426 41972 29438
rect 41916 29374 41918 29426
rect 41970 29374 41972 29426
rect 41692 29316 41748 29326
rect 41692 29222 41748 29260
rect 41916 28980 41972 29374
rect 41692 28924 41972 28980
rect 41356 28702 41358 28754
rect 41410 28702 41412 28754
rect 41356 28644 41412 28702
rect 41356 28578 41412 28588
rect 41468 28868 41524 28878
rect 41468 28082 41524 28812
rect 41692 28642 41748 28924
rect 42028 28756 42084 29484
rect 42252 29474 42308 29484
rect 42364 31780 42420 31790
rect 42364 30882 42420 31724
rect 42700 31556 42756 31566
rect 42700 31462 42756 31500
rect 42364 30830 42366 30882
rect 42418 30830 42420 30882
rect 41692 28590 41694 28642
rect 41746 28590 41748 28642
rect 41692 28578 41748 28590
rect 41804 28700 42084 28756
rect 42140 29204 42196 29214
rect 41468 28030 41470 28082
rect 41522 28030 41524 28082
rect 41468 28018 41524 28030
rect 41804 28196 41860 28700
rect 41916 28532 41972 28542
rect 41916 28438 41972 28476
rect 42028 28532 42084 28542
rect 42140 28532 42196 29148
rect 42028 28530 42196 28532
rect 42028 28478 42030 28530
rect 42082 28478 42196 28530
rect 42028 28476 42196 28478
rect 42252 28980 42308 28990
rect 42028 28466 42084 28476
rect 41804 27860 41860 28140
rect 42252 27972 42308 28924
rect 42364 28084 42420 30830
rect 42812 30548 42868 35868
rect 42924 35700 42980 39340
rect 43260 39060 43316 39342
rect 43316 39004 43428 39060
rect 43260 38994 43316 39004
rect 43036 38834 43092 38846
rect 43036 38782 43038 38834
rect 43090 38782 43092 38834
rect 43036 38724 43092 38782
rect 43036 38658 43092 38668
rect 43148 38834 43204 38846
rect 43148 38782 43150 38834
rect 43202 38782 43204 38834
rect 43148 37828 43204 38782
rect 43260 38836 43316 38846
rect 43260 38742 43316 38780
rect 43148 37762 43204 37772
rect 43036 37378 43092 37390
rect 43036 37326 43038 37378
rect 43090 37326 43092 37378
rect 43036 36036 43092 37326
rect 43260 37268 43316 37278
rect 43036 35970 43092 35980
rect 43148 36932 43204 36942
rect 43148 36594 43204 36876
rect 43148 36542 43150 36594
rect 43202 36542 43204 36594
rect 43148 36484 43204 36542
rect 43148 35922 43204 36428
rect 43148 35870 43150 35922
rect 43202 35870 43204 35922
rect 43148 35858 43204 35870
rect 43260 35700 43316 37212
rect 43372 36372 43428 39004
rect 43484 38164 43540 38174
rect 43484 37490 43540 38108
rect 43596 37828 43652 42588
rect 43820 42196 43876 44942
rect 43932 43764 43988 45838
rect 44268 45780 44324 45790
rect 44156 45106 44212 45118
rect 44156 45054 44158 45106
rect 44210 45054 44212 45106
rect 44156 44884 44212 45054
rect 44156 44818 44212 44828
rect 44268 44660 44324 45724
rect 44380 45668 44436 45678
rect 44380 44882 44436 45612
rect 44380 44830 44382 44882
rect 44434 44830 44436 44882
rect 44380 44818 44436 44830
rect 44268 44604 44436 44660
rect 44268 44436 44324 44446
rect 43932 43698 43988 43708
rect 44044 44434 44324 44436
rect 44044 44382 44270 44434
rect 44322 44382 44324 44434
rect 44044 44380 44324 44382
rect 43932 43538 43988 43550
rect 43932 43486 43934 43538
rect 43986 43486 43988 43538
rect 43932 42754 43988 43486
rect 43932 42702 43934 42754
rect 43986 42702 43988 42754
rect 43932 42420 43988 42702
rect 43932 42354 43988 42364
rect 43708 42140 43876 42196
rect 43708 40404 43764 42140
rect 43820 41970 43876 41982
rect 44044 41972 44100 44380
rect 44268 44370 44324 44380
rect 44380 43652 44436 44604
rect 43820 41918 43822 41970
rect 43874 41918 43876 41970
rect 43820 41860 43876 41918
rect 43820 41188 43876 41804
rect 43820 41122 43876 41132
rect 43932 41916 44100 41972
rect 44156 43596 44436 43652
rect 43708 40338 43764 40348
rect 43932 40628 43988 41916
rect 44044 41748 44100 41758
rect 44044 41654 44100 41692
rect 44156 41410 44212 43596
rect 44380 43426 44436 43438
rect 44380 43374 44382 43426
rect 44434 43374 44436 43426
rect 44268 42532 44324 42542
rect 44268 42438 44324 42476
rect 44380 41972 44436 43374
rect 44492 42980 44548 45948
rect 45388 45668 45444 45678
rect 45276 45332 45332 45342
rect 44828 45220 44884 45230
rect 44828 45126 44884 45164
rect 44604 45106 44660 45118
rect 44604 45054 44606 45106
rect 44658 45054 44660 45106
rect 44604 43762 44660 45054
rect 44940 45108 44996 45118
rect 44940 45014 44996 45052
rect 45276 44994 45332 45276
rect 45276 44942 45278 44994
rect 45330 44942 45332 44994
rect 45276 44930 45332 44942
rect 45052 44322 45108 44334
rect 45052 44270 45054 44322
rect 45106 44270 45108 44322
rect 44604 43710 44606 43762
rect 44658 43710 44660 43762
rect 44604 43698 44660 43710
rect 44828 43876 44884 43886
rect 44492 42914 44548 42924
rect 44828 43650 44884 43820
rect 44828 43598 44830 43650
rect 44882 43598 44884 43650
rect 44828 42868 44884 43598
rect 44940 43540 44996 43550
rect 44940 43446 44996 43484
rect 45052 42980 45108 44270
rect 44828 42802 44884 42812
rect 44940 42924 45108 42980
rect 45276 43426 45332 43438
rect 45276 43374 45278 43426
rect 45330 43374 45332 43426
rect 44940 42644 44996 42924
rect 45164 42868 45220 42878
rect 45276 42868 45332 43374
rect 45220 42812 45332 42868
rect 45164 42802 45220 42812
rect 44268 41916 44436 41972
rect 44716 42588 44996 42644
rect 45052 42754 45108 42766
rect 45052 42702 45054 42754
rect 45106 42702 45108 42754
rect 44268 41748 44324 41916
rect 44268 41682 44324 41692
rect 44380 41746 44436 41758
rect 44380 41694 44382 41746
rect 44434 41694 44436 41746
rect 44156 41358 44158 41410
rect 44210 41358 44212 41410
rect 44156 41346 44212 41358
rect 43820 40292 43876 40302
rect 43820 40198 43876 40236
rect 43820 39620 43876 39630
rect 43932 39620 43988 40572
rect 44156 40964 44212 40974
rect 44156 40514 44212 40908
rect 44380 40740 44436 41694
rect 44380 40674 44436 40684
rect 44492 41300 44548 41310
rect 44156 40462 44158 40514
rect 44210 40462 44212 40514
rect 44156 40450 44212 40462
rect 44492 40402 44548 41244
rect 44604 40964 44660 40974
rect 44716 40964 44772 42588
rect 44828 41972 44884 41982
rect 44828 41878 44884 41916
rect 44940 41970 44996 41982
rect 44940 41918 44942 41970
rect 44994 41918 44996 41970
rect 44940 41636 44996 41918
rect 45052 41748 45108 42702
rect 45276 41860 45332 41870
rect 45276 41766 45332 41804
rect 45052 41682 45108 41692
rect 44940 41570 44996 41580
rect 44940 41076 44996 41086
rect 44940 40982 44996 41020
rect 45276 40964 45332 40974
rect 44660 40908 44772 40964
rect 45164 40962 45332 40964
rect 45164 40910 45278 40962
rect 45330 40910 45332 40962
rect 45164 40908 45332 40910
rect 44604 40898 44660 40908
rect 44492 40350 44494 40402
rect 44546 40350 44548 40402
rect 44492 40338 44548 40350
rect 44940 40404 44996 40414
rect 44940 40310 44996 40348
rect 44380 39732 44436 39742
rect 44380 39730 44548 39732
rect 44380 39678 44382 39730
rect 44434 39678 44548 39730
rect 44380 39676 44548 39678
rect 44380 39666 44436 39676
rect 43820 39618 43988 39620
rect 43820 39566 43822 39618
rect 43874 39566 43988 39618
rect 43820 39564 43988 39566
rect 44044 39618 44100 39630
rect 44044 39566 44046 39618
rect 44098 39566 44100 39618
rect 43820 39554 43876 39564
rect 43820 39396 43876 39406
rect 43820 39394 43988 39396
rect 43820 39342 43822 39394
rect 43874 39342 43988 39394
rect 43820 39340 43988 39342
rect 43820 39330 43876 39340
rect 43708 38834 43764 38846
rect 43708 38782 43710 38834
rect 43762 38782 43764 38834
rect 43708 38164 43764 38782
rect 43708 38098 43764 38108
rect 43820 38722 43876 38734
rect 43820 38670 43822 38722
rect 43874 38670 43876 38722
rect 43596 37762 43652 37772
rect 43820 37604 43876 38670
rect 43484 37438 43486 37490
rect 43538 37438 43540 37490
rect 43484 37426 43540 37438
rect 43708 37548 43876 37604
rect 43484 36372 43540 36382
rect 43372 36370 43540 36372
rect 43372 36318 43486 36370
rect 43538 36318 43540 36370
rect 43372 36316 43540 36318
rect 42924 35634 42980 35644
rect 43148 35644 43316 35700
rect 42924 34916 42980 34926
rect 42924 34802 42980 34860
rect 42924 34750 42926 34802
rect 42978 34750 42980 34802
rect 42924 34738 42980 34750
rect 43036 33122 43092 33134
rect 43036 33070 43038 33122
rect 43090 33070 43092 33122
rect 43036 33012 43092 33070
rect 43036 32946 43092 32956
rect 42812 30482 42868 30492
rect 43148 30212 43204 35644
rect 43260 34692 43316 34702
rect 43484 34692 43540 36316
rect 43596 36258 43652 36270
rect 43596 36206 43598 36258
rect 43650 36206 43652 36258
rect 43596 35924 43652 36206
rect 43708 36036 43764 37548
rect 43932 37380 43988 39340
rect 44044 39060 44100 39566
rect 44492 39620 44548 39676
rect 44492 39564 44772 39620
rect 44380 39508 44436 39518
rect 44380 39396 44436 39452
rect 44268 39340 44436 39396
rect 44044 38668 44100 39004
rect 44156 39284 44212 39294
rect 44156 38834 44212 39228
rect 44268 39058 44324 39340
rect 44268 39006 44270 39058
rect 44322 39006 44324 39058
rect 44268 38994 44324 39006
rect 44156 38782 44158 38834
rect 44210 38782 44212 38834
rect 44156 38770 44212 38782
rect 44492 38946 44548 38958
rect 44492 38894 44494 38946
rect 44546 38894 44548 38946
rect 44044 38612 44212 38668
rect 44044 38164 44100 38174
rect 44044 38070 44100 38108
rect 44156 37940 44212 38612
rect 43820 37324 43988 37380
rect 44044 37884 44212 37940
rect 43820 36372 43876 37324
rect 43932 37156 43988 37166
rect 43932 37062 43988 37100
rect 43820 36306 43876 36316
rect 43932 36260 43988 36270
rect 44044 36260 44100 37884
rect 44492 37492 44548 38894
rect 44716 38276 44772 39564
rect 44828 39508 44884 39518
rect 44828 39414 44884 39452
rect 44940 39396 44996 39406
rect 44940 39394 45108 39396
rect 44940 39342 44942 39394
rect 44994 39342 45108 39394
rect 44940 39340 45108 39342
rect 44940 39330 44996 39340
rect 45052 39172 45108 39340
rect 45052 39106 45108 39116
rect 44828 39060 44884 39070
rect 44828 38966 44884 39004
rect 45164 38948 45220 40908
rect 45276 40898 45332 40908
rect 45276 39730 45332 39742
rect 45276 39678 45278 39730
rect 45330 39678 45332 39730
rect 45276 39284 45332 39678
rect 45276 39218 45332 39228
rect 45388 39060 45444 45612
rect 45836 44548 45892 44558
rect 45836 44454 45892 44492
rect 45948 43652 46004 49200
rect 48412 47124 48468 47134
rect 46844 46004 46900 46014
rect 46844 46002 47348 46004
rect 46844 45950 46846 46002
rect 46898 45950 47348 46002
rect 46844 45948 47348 45950
rect 46844 45938 46900 45948
rect 46508 45780 46564 45790
rect 46508 45686 46564 45724
rect 46732 45666 46788 45678
rect 46732 45614 46734 45666
rect 46786 45614 46788 45666
rect 46732 45556 46788 45614
rect 46732 45490 46788 45500
rect 45948 43586 46004 43596
rect 46844 44884 46900 44894
rect 45612 43540 45668 43550
rect 45500 43204 45556 43214
rect 45500 41972 45556 43148
rect 45500 41906 45556 41916
rect 45612 41186 45668 43484
rect 45836 42980 45892 42990
rect 45836 42886 45892 42924
rect 46620 42532 46676 42542
rect 45612 41134 45614 41186
rect 45666 41134 45668 41186
rect 45500 40516 45556 40526
rect 45500 40402 45556 40460
rect 45500 40350 45502 40402
rect 45554 40350 45556 40402
rect 45500 40338 45556 40350
rect 45388 38994 45444 39004
rect 45164 38892 45332 38948
rect 44828 38836 44884 38846
rect 45276 38836 45332 38892
rect 45500 38836 45556 38846
rect 45612 38836 45668 41134
rect 46284 41860 46340 41870
rect 46284 40852 46340 41804
rect 45948 40516 46004 40526
rect 45836 40404 45892 40414
rect 45836 40310 45892 40348
rect 45276 38780 45444 38836
rect 44828 38668 44884 38780
rect 44828 38612 44996 38668
rect 45276 38666 45332 38678
rect 45276 38614 45278 38666
rect 45330 38614 45332 38666
rect 45276 38612 45332 38614
rect 44828 38276 44884 38286
rect 44716 38220 44828 38276
rect 44828 38210 44884 38220
rect 44940 38162 44996 38612
rect 45164 38556 45332 38612
rect 45164 38276 45220 38556
rect 45388 38500 45444 38780
rect 45556 38780 45668 38836
rect 45500 38770 45556 38780
rect 45164 38210 45220 38220
rect 45276 38444 45444 38500
rect 44940 38110 44942 38162
rect 44994 38110 44996 38162
rect 44940 38098 44996 38110
rect 45052 38164 45108 38174
rect 44492 37426 44548 37436
rect 44492 37266 44548 37278
rect 44492 37214 44494 37266
rect 44546 37214 44548 37266
rect 44492 36596 44548 37214
rect 44940 37156 44996 37166
rect 44940 37062 44996 37100
rect 43932 36258 44100 36260
rect 43932 36206 43934 36258
rect 43986 36206 44100 36258
rect 43932 36204 44100 36206
rect 44156 36540 44884 36596
rect 43820 36036 43876 36046
rect 43708 35980 43820 36036
rect 43820 35970 43876 35980
rect 43596 35858 43652 35868
rect 43596 35700 43652 35710
rect 43596 35606 43652 35644
rect 43260 34690 43540 34692
rect 43260 34638 43262 34690
rect 43314 34638 43540 34690
rect 43260 34636 43540 34638
rect 43260 30434 43316 34636
rect 43932 34580 43988 36204
rect 44156 35922 44212 36540
rect 44828 36482 44884 36540
rect 44828 36430 44830 36482
rect 44882 36430 44884 36482
rect 44828 36418 44884 36430
rect 44604 36372 44660 36382
rect 44660 36316 44772 36372
rect 44604 36306 44660 36316
rect 44268 36258 44324 36270
rect 44268 36206 44270 36258
rect 44322 36206 44324 36258
rect 44268 36036 44324 36206
rect 44268 35970 44324 35980
rect 44156 35870 44158 35922
rect 44210 35870 44212 35922
rect 44044 35588 44100 35598
rect 44044 34802 44100 35532
rect 44156 35026 44212 35870
rect 44716 35810 44772 36316
rect 45052 36260 45108 38108
rect 45164 37940 45220 37950
rect 45164 37846 45220 37884
rect 44828 36204 45108 36260
rect 45164 36260 45220 36270
rect 44828 35922 44884 36204
rect 45164 36166 45220 36204
rect 44828 35870 44830 35922
rect 44882 35870 44884 35922
rect 44828 35858 44884 35870
rect 44716 35758 44718 35810
rect 44770 35758 44772 35810
rect 44716 35746 44772 35758
rect 44156 34974 44158 35026
rect 44210 34974 44212 35026
rect 44156 34962 44212 34974
rect 44492 35588 44548 35598
rect 44044 34750 44046 34802
rect 44098 34750 44100 34802
rect 44044 34738 44100 34750
rect 44268 34804 44324 34814
rect 44268 34710 44324 34748
rect 44380 34692 44436 34702
rect 43932 34524 44212 34580
rect 43708 33346 43764 33358
rect 43708 33294 43710 33346
rect 43762 33294 43764 33346
rect 43372 33234 43428 33246
rect 43708 33236 43764 33294
rect 43372 33182 43374 33234
rect 43426 33182 43428 33234
rect 43372 33012 43428 33182
rect 43372 32946 43428 32956
rect 43596 33180 43708 33236
rect 43596 31778 43652 33180
rect 43708 33170 43764 33180
rect 43932 33234 43988 33246
rect 43932 33182 43934 33234
rect 43986 33182 43988 33234
rect 43820 33124 43876 33162
rect 43820 33058 43876 33068
rect 43932 32788 43988 33182
rect 43596 31726 43598 31778
rect 43650 31726 43652 31778
rect 43596 31714 43652 31726
rect 43820 32732 43988 32788
rect 43260 30382 43262 30434
rect 43314 30382 43316 30434
rect 43260 30370 43316 30382
rect 43372 30660 43428 30670
rect 43260 30212 43316 30222
rect 43148 30156 43260 30212
rect 43260 30146 43316 30156
rect 43372 29764 43428 30604
rect 43596 30548 43652 30558
rect 43820 30548 43876 32732
rect 44156 32676 44212 34524
rect 44380 34242 44436 34636
rect 44380 34190 44382 34242
rect 44434 34190 44436 34242
rect 44380 34178 44436 34190
rect 44492 34244 44548 35532
rect 45276 35140 45332 38444
rect 45724 37156 45780 37166
rect 45052 35084 45332 35140
rect 45388 37044 45444 37054
rect 45388 35698 45444 36988
rect 45500 36482 45556 36494
rect 45500 36430 45502 36482
rect 45554 36430 45556 36482
rect 45500 36036 45556 36430
rect 45500 35970 45556 35980
rect 45724 36258 45780 37100
rect 45836 36596 45892 36606
rect 45948 36596 46004 40460
rect 46284 40514 46340 40796
rect 46508 40628 46564 40638
rect 46508 40534 46564 40572
rect 46284 40462 46286 40514
rect 46338 40462 46340 40514
rect 46284 40450 46340 40462
rect 46396 38388 46452 38398
rect 45836 36594 46004 36596
rect 45836 36542 45838 36594
rect 45890 36542 46004 36594
rect 45836 36540 46004 36542
rect 46060 38276 46116 38286
rect 45836 36530 45892 36540
rect 46060 36482 46116 38220
rect 46060 36430 46062 36482
rect 46114 36430 46116 36482
rect 46060 36418 46116 36430
rect 45724 36206 45726 36258
rect 45778 36206 45780 36258
rect 45388 35646 45390 35698
rect 45442 35646 45444 35698
rect 45388 35252 45444 35646
rect 44940 34692 44996 34702
rect 44940 34598 44996 34636
rect 44492 34188 44884 34244
rect 44828 33460 44884 34188
rect 44940 33460 44996 33470
rect 44828 33458 44996 33460
rect 44828 33406 44942 33458
rect 44994 33406 44996 33458
rect 44828 33404 44996 33406
rect 44828 33236 44884 33246
rect 44828 33142 44884 33180
rect 43932 32620 44212 32676
rect 44380 33124 44436 33134
rect 43932 32002 43988 32620
rect 44044 32452 44100 32462
rect 44044 32450 44324 32452
rect 44044 32398 44046 32450
rect 44098 32398 44324 32450
rect 44044 32396 44324 32398
rect 44044 32386 44100 32396
rect 43932 31950 43934 32002
rect 43986 31950 43988 32002
rect 43932 31938 43988 31950
rect 44156 31890 44212 31902
rect 44156 31838 44158 31890
rect 44210 31838 44212 31890
rect 43932 31778 43988 31790
rect 43932 31726 43934 31778
rect 43986 31726 43988 31778
rect 43932 31556 43988 31726
rect 43932 31490 43988 31500
rect 44156 30994 44212 31838
rect 44268 31218 44324 32396
rect 44380 31890 44436 33068
rect 44380 31838 44382 31890
rect 44434 31838 44436 31890
rect 44380 31826 44436 31838
rect 44716 32562 44772 32574
rect 44716 32510 44718 32562
rect 44770 32510 44772 32562
rect 44716 31892 44772 32510
rect 44716 31826 44772 31836
rect 44268 31166 44270 31218
rect 44322 31166 44324 31218
rect 44268 31154 44324 31166
rect 44380 31668 44436 31678
rect 44156 30942 44158 30994
rect 44210 30942 44212 30994
rect 44156 30930 44212 30942
rect 44380 30994 44436 31612
rect 44828 31556 44884 31566
rect 44828 31462 44884 31500
rect 44940 31444 44996 33404
rect 44940 31378 44996 31388
rect 44380 30942 44382 30994
rect 44434 30942 44436 30994
rect 44380 30930 44436 30942
rect 44492 31276 44884 31332
rect 43932 30772 43988 30782
rect 43932 30678 43988 30716
rect 43652 30492 43764 30548
rect 43820 30492 43988 30548
rect 43596 30482 43652 30492
rect 43260 29708 43428 29764
rect 43484 30210 43540 30222
rect 43484 30158 43486 30210
rect 43538 30158 43540 30210
rect 42812 29538 42868 29550
rect 42812 29486 42814 29538
rect 42866 29486 42868 29538
rect 42700 29316 42756 29326
rect 42700 29222 42756 29260
rect 42588 29204 42644 29214
rect 42588 29110 42644 29148
rect 42700 28868 42756 28878
rect 42700 28530 42756 28812
rect 42812 28644 42868 29486
rect 43260 29204 43316 29708
rect 43372 29540 43428 29550
rect 43372 29426 43428 29484
rect 43372 29374 43374 29426
rect 43426 29374 43428 29426
rect 43372 29362 43428 29374
rect 43260 29148 43428 29204
rect 42812 28578 42868 28588
rect 43260 28644 43316 28654
rect 42700 28478 42702 28530
rect 42754 28478 42756 28530
rect 42700 28466 42756 28478
rect 42924 28532 42980 28542
rect 42924 28530 43204 28532
rect 42924 28478 42926 28530
rect 42978 28478 43204 28530
rect 42924 28476 43204 28478
rect 42924 28466 42980 28476
rect 42364 28018 42420 28028
rect 42812 28418 42868 28430
rect 42812 28366 42814 28418
rect 42866 28366 42868 28418
rect 41580 27858 41860 27860
rect 41580 27806 41806 27858
rect 41858 27806 41860 27858
rect 41580 27804 41860 27806
rect 41468 27076 41524 27086
rect 41580 27076 41636 27804
rect 41804 27794 41860 27804
rect 42028 27916 42308 27972
rect 41468 27074 41636 27076
rect 41468 27022 41470 27074
rect 41522 27022 41636 27074
rect 41468 27020 41636 27022
rect 41468 26908 41524 27020
rect 41244 25106 41300 25116
rect 41356 26852 41524 26908
rect 42028 26908 42084 27916
rect 42588 27746 42644 27758
rect 42588 27694 42590 27746
rect 42642 27694 42644 27746
rect 42140 27188 42196 27198
rect 42140 27094 42196 27132
rect 42028 26852 42308 26908
rect 40908 23884 41188 23940
rect 41244 24836 41300 24846
rect 40572 22932 40628 22942
rect 40572 22594 40628 22876
rect 40572 22542 40574 22594
rect 40626 22542 40628 22594
rect 40572 22530 40628 22542
rect 40796 22484 40852 22494
rect 40684 22428 40796 22484
rect 40460 22260 40516 22270
rect 40460 22166 40516 22204
rect 40572 22260 40628 22270
rect 40684 22260 40740 22428
rect 40796 22418 40852 22428
rect 40572 22258 40740 22260
rect 40572 22206 40574 22258
rect 40626 22206 40740 22258
rect 40572 22204 40740 22206
rect 40572 22194 40628 22204
rect 40348 21980 40516 22036
rect 40124 21858 40180 21868
rect 39004 21422 39006 21474
rect 39058 21422 39060 21474
rect 39004 21410 39060 21422
rect 39228 21586 39284 21598
rect 39228 21534 39230 21586
rect 39282 21534 39284 21586
rect 39228 20916 39284 21534
rect 39788 21476 39844 21486
rect 39788 21382 39844 21420
rect 39228 20822 39284 20860
rect 38444 20130 38612 20132
rect 38444 20078 38446 20130
rect 38498 20078 38612 20130
rect 38444 20076 38612 20078
rect 38444 20066 38500 20076
rect 37212 19966 37214 20018
rect 37266 19966 37268 20018
rect 37212 19954 37268 19966
rect 38556 20020 38612 20076
rect 38780 20132 38836 20142
rect 38780 20038 38836 20076
rect 38556 19954 38612 19964
rect 39004 20020 39060 20030
rect 39004 19926 39060 19964
rect 36540 19906 36596 19918
rect 36540 19854 36542 19906
rect 36594 19854 36596 19906
rect 36540 19460 36596 19854
rect 37436 19906 37492 19918
rect 37436 19854 37438 19906
rect 37490 19854 37492 19906
rect 37436 19460 37492 19854
rect 37884 19908 37940 19918
rect 37884 19906 38052 19908
rect 37884 19854 37886 19906
rect 37938 19854 38052 19906
rect 37884 19852 38052 19854
rect 37884 19842 37940 19852
rect 37548 19796 37604 19806
rect 37548 19794 37828 19796
rect 37548 19742 37550 19794
rect 37602 19742 37828 19794
rect 37548 19740 37828 19742
rect 37548 19730 37604 19740
rect 37772 19572 37828 19740
rect 37772 19516 37940 19572
rect 37436 19404 37828 19460
rect 36540 19394 36596 19404
rect 37772 19346 37828 19404
rect 37772 19294 37774 19346
rect 37826 19294 37828 19346
rect 37772 19282 37828 19294
rect 36988 19234 37044 19246
rect 36988 19182 36990 19234
rect 37042 19182 37044 19234
rect 36652 19124 36708 19134
rect 35644 18722 35700 18732
rect 35868 18732 36036 18788
rect 36316 19010 36372 19022
rect 36316 18958 36318 19010
rect 36370 18958 36372 19010
rect 35644 17666 35700 17678
rect 35644 17614 35646 17666
rect 35698 17614 35700 17666
rect 35644 15428 35700 17614
rect 35756 17666 35812 17678
rect 35756 17614 35758 17666
rect 35810 17614 35812 17666
rect 35756 15540 35812 17614
rect 35868 15652 35924 18732
rect 35868 15586 35924 15596
rect 35980 17666 36036 17678
rect 35980 17614 35982 17666
rect 36034 17614 36036 17666
rect 35756 15474 35812 15484
rect 35980 15540 36036 17614
rect 36316 17668 36372 18958
rect 36652 18676 36708 19068
rect 36652 18338 36708 18620
rect 36652 18286 36654 18338
rect 36706 18286 36708 18338
rect 36652 18274 36708 18286
rect 36988 18452 37044 19182
rect 36316 17602 36372 17612
rect 36092 17556 36148 17566
rect 36092 17554 36260 17556
rect 36092 17502 36094 17554
rect 36146 17502 36260 17554
rect 36092 17500 36260 17502
rect 36092 17490 36148 17500
rect 35980 15474 36036 15484
rect 36092 16884 36148 16894
rect 35644 15362 35700 15372
rect 35980 15204 36036 15242
rect 35532 15092 35812 15148
rect 35980 15138 36036 15148
rect 36092 15148 36148 16828
rect 36204 16212 36260 17500
rect 36540 16884 36596 16894
rect 36540 16790 36596 16828
rect 36988 16884 37044 18396
rect 37100 19012 37156 19022
rect 37100 18340 37156 18956
rect 37660 18564 37716 18574
rect 37884 18564 37940 19516
rect 37996 19348 38052 19852
rect 39564 19906 39620 19918
rect 39564 19854 39566 19906
rect 39618 19854 39620 19906
rect 38108 19794 38164 19806
rect 38108 19742 38110 19794
rect 38162 19742 38164 19794
rect 38108 19684 38164 19742
rect 38108 19628 38388 19684
rect 37996 18676 38052 19292
rect 38108 18676 38164 18686
rect 37996 18674 38164 18676
rect 37996 18622 38110 18674
rect 38162 18622 38164 18674
rect 37996 18620 38164 18622
rect 38108 18610 38164 18620
rect 37884 18508 38052 18564
rect 37660 18452 37716 18508
rect 37548 18450 37716 18452
rect 37548 18398 37662 18450
rect 37714 18398 37716 18450
rect 37548 18396 37716 18398
rect 37996 18452 38052 18508
rect 38332 18562 38388 19628
rect 38892 18676 38948 18686
rect 38892 18582 38948 18620
rect 38332 18510 38334 18562
rect 38386 18510 38388 18562
rect 38220 18452 38276 18462
rect 37996 18450 38276 18452
rect 37996 18398 38222 18450
rect 38274 18398 38276 18450
rect 37996 18396 38276 18398
rect 37100 18338 37380 18340
rect 37100 18286 37102 18338
rect 37154 18286 37380 18338
rect 37100 18284 37380 18286
rect 37100 18274 37156 18284
rect 36988 16818 37044 16828
rect 37100 16996 37156 17006
rect 36316 16212 36372 16222
rect 36204 16156 36316 16212
rect 36316 16146 36372 16156
rect 36428 16212 36484 16222
rect 36428 16210 36596 16212
rect 36428 16158 36430 16210
rect 36482 16158 36596 16210
rect 36428 16156 36596 16158
rect 36428 16146 36484 16156
rect 36428 15316 36484 15326
rect 36428 15222 36484 15260
rect 36092 15092 36372 15148
rect 34188 14532 34244 14542
rect 34188 14438 34244 14476
rect 33964 13916 34356 13972
rect 33628 13906 33684 13916
rect 33292 13748 33348 13758
rect 33068 13636 33124 13646
rect 32620 13074 32788 13076
rect 32620 13022 32622 13074
rect 32674 13022 32788 13074
rect 32620 13020 32788 13022
rect 32956 13634 33124 13636
rect 32956 13582 33070 13634
rect 33122 13582 33124 13634
rect 32956 13580 33124 13582
rect 32620 13010 32676 13020
rect 32508 12796 32676 12852
rect 32396 10782 32398 10834
rect 32450 10782 32452 10834
rect 32396 10770 32452 10782
rect 32508 10500 32564 10510
rect 32508 9826 32564 10444
rect 32508 9774 32510 9826
rect 32562 9774 32564 9826
rect 32508 9762 32564 9774
rect 32620 9380 32676 12796
rect 32956 10500 33012 13580
rect 33068 13570 33124 13580
rect 33180 13524 33236 13534
rect 33180 12850 33236 13468
rect 33180 12798 33182 12850
rect 33234 12798 33236 12850
rect 33180 12628 33236 12798
rect 33068 12516 33124 12526
rect 33068 12178 33124 12460
rect 33068 12126 33070 12178
rect 33122 12126 33124 12178
rect 33068 12114 33124 12126
rect 33180 11844 33236 12572
rect 33180 11778 33236 11788
rect 33292 13522 33348 13692
rect 33964 13748 34020 13758
rect 33964 13654 34020 13692
rect 34188 13746 34244 13758
rect 34188 13694 34190 13746
rect 34242 13694 34244 13746
rect 33292 13470 33294 13522
rect 33346 13470 33348 13522
rect 33292 11954 33348 13470
rect 34076 13634 34132 13646
rect 34076 13582 34078 13634
rect 34130 13582 34132 13634
rect 34076 13188 34132 13582
rect 33740 13186 34132 13188
rect 33740 13134 34078 13186
rect 34130 13134 34132 13186
rect 33740 13132 34132 13134
rect 33516 13076 33572 13086
rect 33516 12982 33572 13020
rect 33404 12964 33460 12974
rect 33404 12870 33460 12908
rect 33740 12962 33796 13132
rect 34076 13122 34132 13132
rect 34188 13188 34244 13694
rect 34300 13188 34356 13916
rect 34412 13412 34468 15092
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 34524 14532 34580 14542
rect 34524 14438 34580 14476
rect 35196 14530 35252 14542
rect 35196 14478 35198 14530
rect 35250 14478 35252 14530
rect 34860 14420 34916 14430
rect 34636 14418 34916 14420
rect 34636 14366 34862 14418
rect 34914 14366 34916 14418
rect 34636 14364 34916 14366
rect 34524 13746 34580 13758
rect 34524 13694 34526 13746
rect 34578 13694 34580 13746
rect 34524 13524 34580 13694
rect 34524 13458 34580 13468
rect 34412 13346 34468 13356
rect 34412 13188 34468 13198
rect 34300 13132 34412 13188
rect 34188 13122 34244 13132
rect 34412 13122 34468 13132
rect 34524 13188 34580 13198
rect 34636 13188 34692 14364
rect 34860 14354 34916 14364
rect 34972 14420 35028 14430
rect 34524 13186 34692 13188
rect 34524 13134 34526 13186
rect 34578 13134 34692 13186
rect 34524 13132 34692 13134
rect 34748 13748 34804 13758
rect 34524 13122 34580 13132
rect 33740 12910 33742 12962
rect 33794 12910 33796 12962
rect 33740 12898 33796 12910
rect 34188 12964 34244 12974
rect 34412 12964 34468 12974
rect 34244 12908 34356 12964
rect 34188 12870 34244 12908
rect 34076 12740 34132 12750
rect 34076 12404 34132 12684
rect 33964 12402 34132 12404
rect 33964 12350 34078 12402
rect 34130 12350 34132 12402
rect 33964 12348 34132 12350
rect 33292 11902 33294 11954
rect 33346 11902 33348 11954
rect 33292 10724 33348 11902
rect 33628 11954 33684 11966
rect 33628 11902 33630 11954
rect 33682 11902 33684 11954
rect 33628 11508 33684 11902
rect 33740 11844 33796 11854
rect 33796 11788 33908 11844
rect 33740 11778 33796 11788
rect 33628 11442 33684 11452
rect 33740 11506 33796 11518
rect 33740 11454 33742 11506
rect 33794 11454 33796 11506
rect 33740 11284 33796 11454
rect 33740 11218 33796 11228
rect 33852 10948 33908 11788
rect 33292 10658 33348 10668
rect 33740 10892 33908 10948
rect 33180 10500 33236 10510
rect 32956 10498 33236 10500
rect 32956 10446 33182 10498
rect 33234 10446 33236 10498
rect 32956 10444 33236 10446
rect 33180 10276 33236 10444
rect 33628 10500 33684 10510
rect 33628 10406 33684 10444
rect 33180 10210 33236 10220
rect 33292 10164 33348 10174
rect 33180 9716 33236 9726
rect 33180 9622 33236 9660
rect 32620 9324 32900 9380
rect 32508 8932 32564 8942
rect 32284 8930 32676 8932
rect 32284 8878 32510 8930
rect 32562 8878 32676 8930
rect 32284 8876 32676 8878
rect 32508 8866 32564 8876
rect 32060 8370 32228 8372
rect 32060 8318 32062 8370
rect 32114 8318 32228 8370
rect 32060 8316 32228 8318
rect 32508 8370 32564 8382
rect 32508 8318 32510 8370
rect 32562 8318 32564 8370
rect 32060 8306 32116 8316
rect 32284 8260 32340 8270
rect 32172 8204 32284 8260
rect 32172 7474 32228 8204
rect 32284 8194 32340 8204
rect 32284 7812 32340 7822
rect 32284 7698 32340 7756
rect 32284 7646 32286 7698
rect 32338 7646 32340 7698
rect 32284 7634 32340 7646
rect 32172 7422 32174 7474
rect 32226 7422 32228 7474
rect 32172 7364 32228 7422
rect 32172 7298 32228 7308
rect 31164 7196 31556 7252
rect 30828 7084 30996 7140
rect 30828 6578 30884 6590
rect 30828 6526 30830 6578
rect 30882 6526 30884 6578
rect 30828 6020 30884 6526
rect 30940 6356 30996 7084
rect 30940 6290 30996 6300
rect 30828 5954 30884 5964
rect 31052 5906 31108 5918
rect 31052 5854 31054 5906
rect 31106 5854 31108 5906
rect 30828 5796 30884 5806
rect 30828 5702 30884 5740
rect 31052 5684 31108 5854
rect 31052 5618 31108 5628
rect 30716 5516 30884 5572
rect 30156 5234 30548 5236
rect 30156 5182 30158 5234
rect 30210 5182 30548 5234
rect 30156 5180 30548 5182
rect 30156 5170 30212 5180
rect 29708 5124 29764 5134
rect 29596 5122 29764 5124
rect 29596 5070 29710 5122
rect 29762 5070 29764 5122
rect 29596 5068 29764 5070
rect 29708 5058 29764 5068
rect 30492 5124 30548 5180
rect 30492 5122 30772 5124
rect 30492 5070 30494 5122
rect 30546 5070 30772 5122
rect 30492 5068 30772 5070
rect 30492 5058 30548 5068
rect 29372 5012 29428 5022
rect 29372 4918 29428 4956
rect 30268 5012 30324 5022
rect 30268 4226 30324 4956
rect 30716 4562 30772 5068
rect 30716 4510 30718 4562
rect 30770 4510 30772 4562
rect 30716 4498 30772 4510
rect 30268 4174 30270 4226
rect 30322 4174 30324 4226
rect 30268 4162 30324 4174
rect 30828 3388 30884 5516
rect 31164 4116 31220 7196
rect 32284 6916 32340 6926
rect 31724 6804 31780 6814
rect 31276 6690 31332 6702
rect 31276 6638 31278 6690
rect 31330 6638 31332 6690
rect 31276 6580 31332 6638
rect 31500 6692 31556 6702
rect 31500 6598 31556 6636
rect 31276 6514 31332 6524
rect 31724 6130 31780 6748
rect 32172 6690 32228 6702
rect 32172 6638 32174 6690
rect 32226 6638 32228 6690
rect 31836 6468 31892 6478
rect 32172 6468 32228 6638
rect 31836 6466 32228 6468
rect 31836 6414 31838 6466
rect 31890 6414 32228 6466
rect 31836 6412 32228 6414
rect 31836 6402 31892 6412
rect 31724 6078 31726 6130
rect 31778 6078 31780 6130
rect 31500 5906 31556 5918
rect 31500 5854 31502 5906
rect 31554 5854 31556 5906
rect 31500 5796 31556 5854
rect 31500 5348 31556 5740
rect 31500 5282 31556 5292
rect 31612 5906 31668 5918
rect 31612 5854 31614 5906
rect 31666 5854 31668 5906
rect 31388 5236 31444 5246
rect 31276 5010 31332 5022
rect 31276 4958 31278 5010
rect 31330 4958 31332 5010
rect 31276 4562 31332 4958
rect 31276 4510 31278 4562
rect 31330 4510 31332 4562
rect 31276 4498 31332 4510
rect 31388 4450 31444 5180
rect 31612 5012 31668 5854
rect 31612 4946 31668 4956
rect 31724 4562 31780 6078
rect 31948 6244 32004 6254
rect 31948 6018 32004 6188
rect 31948 5966 31950 6018
rect 32002 5966 32004 6018
rect 31948 5954 32004 5966
rect 32172 5684 32228 6412
rect 32060 5124 32116 5134
rect 31724 4510 31726 4562
rect 31778 4510 31780 4562
rect 31724 4498 31780 4510
rect 31836 4564 31892 4574
rect 32060 4564 32116 5068
rect 31836 4562 32116 4564
rect 31836 4510 31838 4562
rect 31890 4510 32116 4562
rect 31836 4508 32116 4510
rect 31836 4498 31892 4508
rect 31388 4398 31390 4450
rect 31442 4398 31444 4450
rect 31388 4386 31444 4398
rect 31948 4340 32004 4350
rect 32172 4340 32228 5628
rect 31948 4338 32228 4340
rect 31948 4286 31950 4338
rect 32002 4286 32228 4338
rect 31948 4284 32228 4286
rect 32284 4338 32340 6860
rect 32396 6804 32452 6814
rect 32396 6710 32452 6748
rect 32508 6804 32564 8318
rect 32620 8372 32676 8876
rect 32620 7364 32676 8316
rect 32620 7298 32676 7308
rect 32732 7028 32788 7038
rect 32620 6804 32676 6814
rect 32508 6748 32620 6804
rect 32508 6468 32564 6748
rect 32620 6738 32676 6748
rect 32284 4286 32286 4338
rect 32338 4286 32340 4338
rect 31948 4274 32004 4284
rect 32284 4274 32340 4286
rect 32396 6412 32564 6468
rect 32732 6690 32788 6972
rect 32732 6638 32734 6690
rect 32786 6638 32788 6690
rect 31164 4050 31220 4060
rect 32396 3388 32452 6412
rect 32508 5908 32564 5918
rect 32508 5794 32564 5852
rect 32508 5742 32510 5794
rect 32562 5742 32564 5794
rect 32508 5572 32564 5742
rect 32732 5796 32788 6638
rect 32844 5908 32900 9324
rect 33292 8930 33348 10108
rect 33292 8878 33294 8930
rect 33346 8878 33348 8930
rect 33292 8260 33348 8878
rect 33292 8194 33348 8204
rect 32956 8036 33012 8046
rect 33292 8036 33348 8046
rect 32956 8034 33348 8036
rect 32956 7982 32958 8034
rect 33010 7982 33294 8034
rect 33346 7982 33348 8034
rect 32956 7980 33348 7982
rect 32956 7588 33012 7980
rect 33292 7970 33348 7980
rect 33292 7812 33348 7822
rect 33068 7588 33124 7598
rect 32956 7532 33068 7588
rect 33068 7494 33124 7532
rect 33068 6692 33124 6702
rect 33068 6598 33124 6636
rect 33292 6690 33348 7756
rect 33740 7700 33796 10892
rect 33964 10724 34020 12348
rect 34076 12338 34132 12348
rect 34076 11620 34132 11630
rect 34076 11526 34132 11564
rect 34076 11396 34132 11406
rect 34300 11396 34356 12908
rect 34412 12962 34692 12964
rect 34412 12910 34414 12962
rect 34466 12910 34692 12962
rect 34412 12908 34692 12910
rect 34412 12898 34468 12908
rect 34412 12404 34468 12414
rect 34412 12310 34468 12348
rect 34636 11732 34692 12908
rect 34748 12740 34804 13692
rect 34972 13746 35028 14364
rect 34972 13694 34974 13746
rect 35026 13694 35028 13746
rect 34972 13682 35028 13694
rect 35196 13524 35252 14478
rect 35420 14418 35476 14430
rect 35420 14366 35422 14418
rect 35474 14366 35476 14418
rect 35308 14306 35364 14318
rect 35308 14254 35310 14306
rect 35362 14254 35364 14306
rect 35308 13524 35364 14254
rect 35420 14308 35476 14366
rect 35420 13748 35476 14252
rect 35420 13682 35476 13692
rect 35644 13634 35700 13646
rect 35644 13582 35646 13634
rect 35698 13582 35700 13634
rect 35308 13468 35588 13524
rect 35196 13458 35252 13468
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35084 12964 35140 12974
rect 35084 12870 35140 12908
rect 35532 12962 35588 13468
rect 35532 12910 35534 12962
rect 35586 12910 35588 12962
rect 35532 12898 35588 12910
rect 34748 12674 34804 12684
rect 34860 12850 34916 12862
rect 34860 12798 34862 12850
rect 34914 12798 34916 12850
rect 34860 12516 34916 12798
rect 35308 12740 35364 12750
rect 35644 12740 35700 13582
rect 35756 13188 35812 15092
rect 35980 14644 36036 14654
rect 35868 14306 35924 14318
rect 35868 14254 35870 14306
rect 35922 14254 35924 14306
rect 35868 14196 35924 14254
rect 35868 14130 35924 14140
rect 35756 13122 35812 13132
rect 35308 12738 35700 12740
rect 35308 12686 35310 12738
rect 35362 12686 35700 12738
rect 35308 12684 35700 12686
rect 35868 13074 35924 13086
rect 35868 13022 35870 13074
rect 35922 13022 35924 13074
rect 35308 12674 35364 12684
rect 34860 12450 34916 12460
rect 35868 12404 35924 13022
rect 35980 13076 36036 14588
rect 36316 14420 36372 15092
rect 36540 14532 36596 16156
rect 37100 16210 37156 16940
rect 37212 16770 37268 16782
rect 37212 16718 37214 16770
rect 37266 16718 37268 16770
rect 37212 16436 37268 16718
rect 37324 16548 37380 18284
rect 37324 16482 37380 16492
rect 37212 16370 37268 16380
rect 37100 16158 37102 16210
rect 37154 16158 37156 16210
rect 37100 16146 37156 16158
rect 37324 15540 37380 15550
rect 36372 14364 36484 14420
rect 36316 14326 36372 14364
rect 35980 13010 36036 13020
rect 36092 13748 36148 13758
rect 35868 12348 36036 12404
rect 34524 11396 34580 11406
rect 34300 11340 34524 11396
rect 34076 10948 34132 11340
rect 34524 11302 34580 11340
rect 34188 11284 34244 11294
rect 34188 11190 34244 11228
rect 34076 10882 34132 10892
rect 34524 11060 34580 11070
rect 34524 10836 34580 11004
rect 34636 10948 34692 11676
rect 34748 12178 34804 12190
rect 34748 12126 34750 12178
rect 34802 12126 34804 12178
rect 34748 11508 34804 12126
rect 34860 12180 34916 12190
rect 34860 12086 34916 12124
rect 34972 12178 35028 12190
rect 34972 12126 34974 12178
rect 35026 12126 35028 12178
rect 34972 12068 35028 12126
rect 34972 12002 35028 12012
rect 35420 12178 35476 12190
rect 35420 12126 35422 12178
rect 35474 12126 35476 12178
rect 34860 11956 34916 11966
rect 35420 11956 35476 12126
rect 35532 12180 35588 12190
rect 35532 12086 35588 12124
rect 35868 12178 35924 12190
rect 35868 12126 35870 12178
rect 35922 12126 35924 12178
rect 35644 12068 35700 12078
rect 35700 12012 35812 12068
rect 35644 12002 35700 12012
rect 35420 11900 35588 11956
rect 34860 11618 34916 11900
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 34860 11566 34862 11618
rect 34914 11566 34916 11618
rect 34860 11554 34916 11566
rect 34748 11442 34804 11452
rect 35084 11396 35140 11406
rect 35084 11302 35140 11340
rect 35532 11396 35588 11900
rect 35532 11302 35588 11340
rect 35756 11394 35812 12012
rect 35868 11956 35924 12126
rect 35980 11956 36036 12348
rect 36092 12178 36148 13692
rect 36204 12962 36260 12974
rect 36204 12910 36206 12962
rect 36258 12910 36260 12962
rect 36204 12404 36260 12910
rect 36204 12338 36260 12348
rect 36316 12628 36372 12638
rect 36092 12126 36094 12178
rect 36146 12126 36148 12178
rect 36092 12114 36148 12126
rect 36316 12180 36372 12572
rect 36316 12086 36372 12124
rect 35980 11900 36148 11956
rect 35868 11890 35924 11900
rect 35868 11508 35924 11518
rect 35868 11414 35924 11452
rect 35756 11342 35758 11394
rect 35810 11342 35812 11394
rect 35756 11330 35812 11342
rect 34748 11172 34804 11182
rect 34748 11078 34804 11116
rect 36092 11060 36148 11900
rect 36092 10994 36148 11004
rect 34860 10948 34916 10958
rect 34636 10892 34860 10948
rect 34524 10780 34692 10836
rect 34188 10724 34244 10734
rect 33964 10722 34244 10724
rect 33964 10670 34190 10722
rect 34242 10670 34244 10722
rect 33964 10668 34244 10670
rect 34188 9716 34244 10668
rect 34300 10722 34356 10734
rect 34300 10670 34302 10722
rect 34354 10670 34356 10722
rect 34300 10164 34356 10670
rect 34300 10098 34356 10108
rect 34524 10610 34580 10622
rect 34524 10558 34526 10610
rect 34578 10558 34580 10610
rect 34188 9650 34244 9660
rect 34412 8932 34468 8942
rect 33740 7606 33796 7644
rect 33852 8258 33908 8270
rect 33852 8206 33854 8258
rect 33906 8206 33908 8258
rect 33852 7924 33908 8206
rect 34188 8148 34244 8158
rect 34188 8054 34244 8092
rect 34412 8034 34468 8876
rect 34524 8258 34580 10558
rect 34524 8206 34526 8258
rect 34578 8206 34580 8258
rect 34524 8194 34580 8206
rect 34412 7982 34414 8034
rect 34466 7982 34468 8034
rect 34412 7970 34468 7982
rect 33404 7586 33460 7598
rect 33404 7534 33406 7586
rect 33458 7534 33460 7586
rect 33404 6916 33460 7534
rect 33852 7476 33908 7868
rect 33852 7410 33908 7420
rect 34300 7924 34356 7934
rect 34636 7924 34692 10780
rect 34860 10834 34916 10892
rect 34860 10782 34862 10834
rect 34914 10782 34916 10834
rect 34860 10770 34916 10782
rect 35532 10834 35588 10846
rect 35532 10782 35534 10834
rect 35586 10782 35588 10834
rect 35308 10724 35364 10734
rect 35308 10630 35364 10668
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35308 9940 35364 9950
rect 35308 9044 35364 9884
rect 35308 8978 35364 8988
rect 35420 8932 35476 8942
rect 35420 8838 35476 8876
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 34748 8372 34804 8382
rect 34748 8258 34804 8316
rect 34748 8206 34750 8258
rect 34802 8206 34804 8258
rect 34748 8194 34804 8206
rect 34972 8260 35028 8270
rect 34300 7362 34356 7868
rect 34300 7310 34302 7362
rect 34354 7310 34356 7362
rect 33516 6916 33572 6926
rect 33404 6860 33516 6916
rect 34300 6916 34356 7310
rect 34524 7868 34692 7924
rect 34860 8036 34916 8046
rect 34524 7028 34580 7868
rect 34636 7700 34692 7710
rect 34636 7588 34692 7644
rect 34748 7588 34804 7598
rect 34636 7586 34804 7588
rect 34636 7534 34750 7586
rect 34802 7534 34804 7586
rect 34636 7532 34804 7534
rect 34748 7522 34804 7532
rect 34524 6972 34692 7028
rect 34300 6860 34580 6916
rect 33292 6638 33294 6690
rect 33346 6638 33348 6690
rect 33292 6580 33348 6638
rect 33516 6692 33572 6860
rect 33628 6692 33684 6702
rect 33516 6690 33684 6692
rect 33516 6638 33630 6690
rect 33682 6638 33684 6690
rect 33516 6636 33684 6638
rect 33628 6626 33684 6636
rect 34300 6690 34356 6702
rect 34300 6638 34302 6690
rect 34354 6638 34356 6690
rect 33292 6514 33348 6524
rect 33180 6466 33236 6478
rect 33180 6414 33182 6466
rect 33234 6414 33236 6466
rect 32844 5842 32900 5852
rect 32956 6020 33012 6030
rect 32732 5730 32788 5740
rect 32508 5506 32564 5516
rect 32956 4228 33012 5964
rect 33068 5908 33124 5918
rect 33180 5908 33236 6414
rect 33628 6468 33684 6478
rect 33068 5906 33236 5908
rect 33068 5854 33070 5906
rect 33122 5854 33236 5906
rect 33068 5852 33236 5854
rect 33516 6018 33572 6030
rect 33516 5966 33518 6018
rect 33570 5966 33572 6018
rect 33068 5842 33124 5852
rect 33180 5684 33236 5694
rect 33180 5590 33236 5628
rect 33516 5460 33572 5966
rect 33516 5394 33572 5404
rect 33404 5348 33460 5358
rect 33404 5234 33460 5292
rect 33404 5182 33406 5234
rect 33458 5182 33460 5234
rect 33404 5170 33460 5182
rect 33068 4228 33124 4238
rect 32956 4226 33124 4228
rect 32956 4174 33070 4226
rect 33122 4174 33124 4226
rect 32956 4172 33124 4174
rect 33068 4162 33124 4172
rect 28700 3332 28980 3388
rect 28924 2996 28980 3332
rect 28924 2930 28980 2940
rect 30380 3332 30884 3388
rect 32284 3332 32452 3388
rect 27580 2706 27636 2716
rect 30380 1540 30436 3332
rect 32284 2324 32340 3332
rect 33628 3220 33684 6412
rect 34076 6466 34132 6478
rect 34076 6414 34078 6466
rect 34130 6414 34132 6466
rect 34076 6244 34132 6414
rect 34300 6468 34356 6638
rect 34300 6402 34356 6412
rect 33740 6188 34132 6244
rect 33740 6018 33796 6188
rect 33740 5966 33742 6018
rect 33794 5966 33796 6018
rect 33740 5954 33796 5966
rect 33740 5796 33796 5806
rect 33740 5348 33796 5740
rect 33852 5572 33908 6188
rect 34076 6132 34132 6188
rect 34076 6066 34132 6076
rect 33964 6020 34020 6030
rect 33964 5926 34020 5964
rect 34412 5908 34468 5918
rect 34412 5814 34468 5852
rect 34076 5794 34132 5806
rect 34076 5742 34078 5794
rect 34130 5742 34132 5794
rect 34076 5684 34132 5742
rect 34076 5618 34132 5628
rect 33852 5506 33908 5516
rect 34188 5572 34244 5582
rect 34076 5460 34132 5470
rect 33852 5348 33908 5358
rect 33740 5346 33908 5348
rect 33740 5294 33854 5346
rect 33906 5294 33908 5346
rect 33740 5292 33908 5294
rect 33852 5282 33908 5292
rect 33740 5124 33796 5134
rect 33740 5030 33796 5068
rect 34076 5010 34132 5404
rect 34188 5124 34244 5516
rect 34412 5124 34468 5134
rect 34188 5122 34468 5124
rect 34188 5070 34414 5122
rect 34466 5070 34468 5122
rect 34188 5068 34468 5070
rect 34412 5058 34468 5068
rect 34076 4958 34078 5010
rect 34130 4958 34132 5010
rect 34076 4946 34132 4958
rect 33628 3154 33684 3164
rect 34412 2660 34468 2670
rect 34524 2660 34580 6860
rect 34636 5460 34692 6972
rect 34860 6804 34916 7980
rect 34972 7588 35028 8204
rect 35532 8260 35588 10782
rect 36204 10724 36260 10734
rect 36204 10630 36260 10668
rect 35644 10610 35700 10622
rect 35644 10558 35646 10610
rect 35698 10558 35700 10610
rect 35644 10388 35700 10558
rect 35868 10610 35924 10622
rect 35868 10558 35870 10610
rect 35922 10558 35924 10610
rect 35644 10322 35700 10332
rect 35756 10500 35812 10510
rect 35756 9604 35812 10444
rect 35532 8194 35588 8204
rect 35644 9602 35812 9604
rect 35644 9550 35758 9602
rect 35810 9550 35812 9602
rect 35644 9548 35812 9550
rect 35644 9268 35700 9548
rect 35756 9538 35812 9548
rect 35868 10388 35924 10558
rect 36428 10500 36484 14364
rect 36540 13636 36596 14476
rect 36876 15314 36932 15326
rect 36876 15262 36878 15314
rect 36930 15262 36932 15314
rect 36876 14420 36932 15262
rect 37324 15148 37380 15484
rect 36876 14354 36932 14364
rect 37100 15092 37380 15148
rect 36988 14306 37044 14318
rect 36988 14254 36990 14306
rect 37042 14254 37044 14306
rect 36988 14084 37044 14254
rect 36988 14018 37044 14028
rect 37100 13748 37156 15092
rect 37324 14532 37380 14542
rect 37324 14438 37380 14476
rect 37100 13682 37156 13692
rect 36540 13570 36596 13580
rect 37100 12740 37156 12750
rect 37100 12646 37156 12684
rect 36988 12516 37044 12526
rect 36652 12404 36708 12414
rect 36652 12310 36708 12348
rect 36540 12178 36596 12190
rect 36540 12126 36542 12178
rect 36594 12126 36596 12178
rect 36540 11620 36596 12126
rect 36540 11554 36596 11564
rect 36876 12068 36932 12078
rect 36876 11508 36932 12012
rect 36876 11442 36932 11452
rect 36988 11844 37044 12460
rect 36988 10834 37044 11788
rect 37100 12292 37156 12302
rect 37100 11506 37156 12236
rect 37548 11788 37604 18396
rect 37660 18386 37716 18396
rect 38220 18386 38276 18396
rect 38332 17108 38388 18510
rect 39004 18562 39060 18574
rect 39004 18510 39006 18562
rect 39058 18510 39060 18562
rect 39004 18452 39060 18510
rect 39564 18564 39620 19854
rect 40012 19906 40068 19918
rect 40012 19854 40014 19906
rect 40066 19854 40068 19906
rect 39564 18498 39620 18508
rect 39676 19796 39732 19806
rect 39004 18386 39060 18396
rect 39676 18450 39732 19740
rect 39900 19348 39956 19358
rect 39900 19254 39956 19292
rect 39676 18398 39678 18450
rect 39730 18398 39732 18450
rect 39676 18386 39732 18398
rect 39452 18340 39508 18350
rect 39116 18338 39508 18340
rect 39116 18286 39454 18338
rect 39506 18286 39508 18338
rect 39116 18284 39508 18286
rect 38892 18228 38948 18238
rect 39116 18228 39172 18284
rect 39452 18274 39508 18284
rect 38892 18226 39172 18228
rect 38892 18174 38894 18226
rect 38946 18174 39172 18226
rect 38892 18172 39172 18174
rect 38892 18162 38948 18172
rect 38332 17042 38388 17052
rect 38444 17778 38500 17790
rect 38444 17726 38446 17778
rect 38498 17726 38500 17778
rect 37772 16996 37828 17006
rect 37660 15988 37716 15998
rect 37660 15894 37716 15932
rect 37772 15538 37828 16940
rect 38444 16884 38500 17726
rect 39004 17668 39060 17678
rect 39004 16996 39060 17612
rect 40012 17668 40068 19854
rect 40236 19908 40292 19918
rect 40236 19346 40292 19852
rect 40236 19294 40238 19346
rect 40290 19294 40292 19346
rect 40236 19282 40292 19294
rect 40348 18340 40404 18350
rect 40348 18246 40404 18284
rect 40012 17602 40068 17612
rect 39004 16930 39060 16940
rect 40236 17108 40292 17118
rect 37884 16100 37940 16110
rect 37884 16006 37940 16044
rect 38444 16098 38500 16828
rect 40124 16884 40180 16894
rect 38444 16046 38446 16098
rect 38498 16046 38500 16098
rect 38444 16034 38500 16046
rect 39004 16772 39060 16782
rect 38108 15988 38164 15998
rect 38108 15894 38164 15932
rect 38780 15988 38836 15998
rect 37996 15876 38052 15886
rect 37996 15782 38052 15820
rect 38668 15764 38724 15774
rect 37772 15486 37774 15538
rect 37826 15486 37828 15538
rect 37772 15474 37828 15486
rect 38220 15652 38276 15662
rect 38220 15538 38276 15596
rect 38220 15486 38222 15538
rect 38274 15486 38276 15538
rect 38220 15474 38276 15486
rect 38668 15538 38724 15708
rect 38668 15486 38670 15538
rect 38722 15486 38724 15538
rect 38668 15474 38724 15486
rect 38780 15204 38836 15932
rect 39004 15148 39060 16716
rect 39340 16772 39396 16782
rect 39676 16772 39732 16782
rect 39340 16770 39732 16772
rect 39340 16718 39342 16770
rect 39394 16718 39678 16770
rect 39730 16718 39732 16770
rect 39340 16716 39732 16718
rect 39228 16212 39284 16222
rect 39228 16118 39284 16156
rect 39340 16100 39396 16716
rect 39676 16706 39732 16716
rect 39900 16660 39956 16670
rect 39900 16658 40068 16660
rect 39900 16606 39902 16658
rect 39954 16606 40068 16658
rect 39900 16604 40068 16606
rect 39900 16594 39956 16604
rect 39340 16034 39396 16044
rect 39788 16436 39844 16446
rect 39676 15876 39732 15886
rect 39676 15426 39732 15820
rect 39788 15538 39844 16380
rect 39788 15486 39790 15538
rect 39842 15486 39844 15538
rect 39788 15474 39844 15486
rect 39900 15540 39956 15550
rect 39900 15446 39956 15484
rect 39676 15374 39678 15426
rect 39730 15374 39732 15426
rect 39676 15362 39732 15374
rect 37772 14418 37828 14430
rect 37772 14366 37774 14418
rect 37826 14366 37828 14418
rect 37660 14308 37716 14318
rect 37772 14308 37828 14366
rect 38220 14420 38276 14430
rect 38220 14326 38276 14364
rect 37716 14252 37828 14308
rect 37884 14308 37940 14318
rect 37660 14242 37716 14252
rect 37772 13634 37828 13646
rect 37772 13582 37774 13634
rect 37826 13582 37828 13634
rect 37772 13524 37828 13582
rect 37772 13458 37828 13468
rect 37884 12962 37940 14252
rect 38444 14084 38500 14094
rect 38444 13748 38500 14028
rect 38332 13522 38388 13534
rect 38332 13470 38334 13522
rect 38386 13470 38388 13522
rect 38332 13076 38388 13470
rect 38444 13524 38500 13692
rect 38668 13746 38724 13758
rect 38668 13694 38670 13746
rect 38722 13694 38724 13746
rect 38668 13636 38724 13694
rect 38780 13748 38836 15148
rect 38892 15092 39060 15148
rect 39900 15204 39956 15214
rect 38892 14532 38948 15092
rect 39788 14756 39844 14766
rect 39900 14756 39956 15148
rect 40012 14756 40068 16604
rect 39788 14754 40068 14756
rect 39788 14702 39790 14754
rect 39842 14702 40068 14754
rect 39788 14700 40068 14702
rect 39788 14690 39844 14700
rect 38892 14438 38948 14476
rect 39452 14420 39508 14430
rect 39676 14420 39732 14430
rect 39452 14418 39732 14420
rect 39452 14366 39454 14418
rect 39506 14366 39678 14418
rect 39730 14366 39732 14418
rect 39452 14364 39732 14366
rect 39452 14354 39508 14364
rect 39676 14354 39732 14364
rect 39116 14306 39172 14318
rect 39116 14254 39118 14306
rect 39170 14254 39172 14306
rect 39116 14084 39172 14254
rect 39340 14306 39396 14318
rect 39340 14254 39342 14306
rect 39394 14254 39396 14306
rect 39340 14196 39396 14254
rect 39340 14140 39844 14196
rect 39116 14028 39620 14084
rect 38892 13748 38948 13758
rect 38780 13746 38948 13748
rect 38780 13694 38894 13746
rect 38946 13694 38948 13746
rect 38780 13692 38948 13694
rect 38892 13682 38948 13692
rect 39228 13748 39284 13758
rect 39228 13654 39284 13692
rect 39564 13746 39620 14028
rect 39564 13694 39566 13746
rect 39618 13694 39620 13746
rect 38668 13580 38836 13636
rect 38780 13524 38836 13580
rect 39340 13634 39396 13646
rect 39340 13582 39342 13634
rect 39394 13582 39396 13634
rect 39340 13524 39396 13582
rect 38444 13468 38724 13524
rect 38780 13468 39396 13524
rect 39452 13636 39508 13646
rect 38556 13076 38612 13086
rect 38332 13074 38612 13076
rect 38332 13022 38558 13074
rect 38610 13022 38612 13074
rect 38332 13020 38612 13022
rect 38556 13010 38612 13020
rect 37884 12910 37886 12962
rect 37938 12910 37940 12962
rect 37884 12898 37940 12910
rect 37100 11454 37102 11506
rect 37154 11454 37156 11506
rect 37100 11396 37156 11454
rect 37100 11330 37156 11340
rect 37324 11732 37604 11788
rect 38332 12852 38388 12862
rect 38332 11844 38388 12796
rect 36988 10782 36990 10834
rect 37042 10782 37044 10834
rect 36988 10770 37044 10782
rect 36428 10434 36484 10444
rect 36540 10610 36596 10622
rect 36540 10558 36542 10610
rect 36594 10558 36596 10610
rect 35084 8146 35140 8158
rect 35084 8094 35086 8146
rect 35138 8094 35140 8146
rect 35084 7812 35140 8094
rect 35420 8148 35476 8158
rect 35420 8054 35476 8092
rect 35196 8036 35252 8046
rect 35196 7942 35252 7980
rect 35532 8036 35588 8046
rect 35532 7942 35588 7980
rect 35644 7812 35700 9212
rect 35868 8708 35924 10332
rect 36540 10164 36596 10558
rect 36540 10098 36596 10108
rect 36988 10164 37044 10174
rect 36092 9828 36148 9838
rect 36092 9734 36148 9772
rect 36988 9826 37044 10108
rect 36988 9774 36990 9826
rect 37042 9774 37044 9826
rect 36988 9762 37044 9774
rect 37212 10052 37268 10062
rect 37212 9826 37268 9996
rect 37212 9774 37214 9826
rect 37266 9774 37268 9826
rect 37212 9762 37268 9774
rect 36652 9716 36708 9726
rect 36428 9604 36484 9614
rect 36428 9510 36484 9548
rect 36652 9266 36708 9660
rect 37100 9604 37156 9614
rect 36652 9214 36654 9266
rect 36706 9214 36708 9266
rect 36652 9202 36708 9214
rect 36876 9602 37156 9604
rect 36876 9550 37102 9602
rect 37154 9550 37156 9602
rect 36876 9548 37156 9550
rect 36092 9044 36148 9054
rect 36092 8950 36148 8988
rect 35868 8642 35924 8652
rect 35980 8484 36036 8494
rect 36316 8484 36372 8494
rect 35868 8428 35980 8484
rect 36036 8482 36372 8484
rect 36036 8430 36318 8482
rect 36370 8430 36372 8482
rect 36036 8428 36372 8430
rect 35868 8258 35924 8428
rect 35980 8418 36036 8428
rect 36316 8418 36372 8428
rect 35868 8206 35870 8258
rect 35922 8206 35924 8258
rect 35868 8194 35924 8206
rect 36204 8260 36260 8270
rect 36204 8166 36260 8204
rect 35756 8148 35812 8158
rect 35756 8054 35812 8092
rect 36316 8036 36372 8046
rect 35084 7746 35140 7756
rect 35420 7756 35700 7812
rect 35868 8034 36372 8036
rect 35868 7982 36318 8034
rect 36370 7982 36372 8034
rect 35868 7980 36372 7982
rect 35196 7588 35252 7598
rect 34972 7586 35252 7588
rect 34972 7534 35198 7586
rect 35250 7534 35252 7586
rect 34972 7532 35252 7534
rect 35196 7522 35252 7532
rect 35084 7308 35308 7364
rect 35084 6804 35140 7308
rect 35252 7252 35308 7308
rect 35420 7252 35476 7756
rect 35868 7700 35924 7980
rect 36316 7970 36372 7980
rect 35532 7644 35868 7700
rect 35532 7474 35588 7644
rect 35868 7606 35924 7644
rect 35532 7422 35534 7474
rect 35586 7422 35588 7474
rect 35532 7410 35588 7422
rect 36204 7588 36260 7598
rect 36204 7474 36260 7532
rect 36764 7588 36820 7598
rect 36876 7588 36932 9548
rect 37100 9538 37156 9548
rect 37212 9604 37268 9614
rect 37324 9604 37380 11732
rect 37436 11620 37492 11630
rect 37436 11526 37492 11564
rect 37548 11508 37604 11518
rect 37548 10722 37604 11452
rect 37996 11396 38052 11406
rect 37996 11302 38052 11340
rect 37548 10670 37550 10722
rect 37602 10670 37604 10722
rect 37548 10658 37604 10670
rect 37996 10612 38052 10622
rect 37660 10610 38052 10612
rect 37660 10558 37998 10610
rect 38050 10558 38052 10610
rect 37660 10556 38052 10558
rect 37660 10500 37716 10556
rect 37996 10546 38052 10556
rect 37268 9548 37380 9604
rect 37548 10444 37716 10500
rect 37548 9714 37604 10444
rect 37772 10388 37828 10398
rect 37772 10294 37828 10332
rect 38220 10386 38276 10398
rect 38220 10334 38222 10386
rect 38274 10334 38276 10386
rect 37548 9662 37550 9714
rect 37602 9662 37604 9714
rect 37100 9268 37156 9278
rect 37100 9174 37156 9212
rect 37100 8596 37156 8606
rect 37100 8372 37156 8540
rect 37212 8484 37268 9548
rect 37212 8418 37268 8428
rect 37100 8278 37156 8316
rect 36820 7532 36932 7588
rect 37100 8148 37156 8158
rect 36764 7494 36820 7532
rect 36204 7422 36206 7474
rect 36258 7422 36260 7474
rect 36204 7410 36260 7422
rect 36988 7474 37044 7486
rect 36988 7422 36990 7474
rect 37042 7422 37044 7474
rect 36428 7362 36484 7374
rect 36428 7310 36430 7362
rect 36482 7310 36484 7362
rect 35252 7196 35476 7252
rect 35532 7252 35588 7262
rect 36428 7252 36484 7310
rect 35532 7250 35812 7252
rect 35532 7198 35534 7250
rect 35586 7198 35812 7250
rect 35532 7196 35812 7198
rect 35532 7186 35588 7196
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35644 7028 35700 7038
rect 35196 7018 35460 7028
rect 35532 6972 35644 7028
rect 35308 6916 35364 6926
rect 35532 6916 35588 6972
rect 35644 6962 35700 6972
rect 35308 6914 35588 6916
rect 35308 6862 35310 6914
rect 35362 6862 35588 6914
rect 35308 6860 35588 6862
rect 35308 6850 35364 6860
rect 35756 6804 35812 7196
rect 36428 7186 36484 7196
rect 36876 7362 36932 7374
rect 36876 7310 36878 7362
rect 36930 7310 36932 7362
rect 35980 6804 36036 6814
rect 35084 6748 35252 6804
rect 34860 6356 34916 6748
rect 35196 6692 35252 6748
rect 35420 6748 35812 6804
rect 35868 6748 35980 6804
rect 35196 6636 35364 6692
rect 34860 6290 34916 6300
rect 35196 6468 35252 6478
rect 34748 6244 34804 6254
rect 34748 6130 34804 6188
rect 34748 6078 34750 6130
rect 34802 6078 34804 6130
rect 34748 6066 34804 6078
rect 35196 6130 35252 6412
rect 35196 6078 35198 6130
rect 35250 6078 35252 6130
rect 35196 6066 35252 6078
rect 35308 5796 35364 6636
rect 35420 6690 35476 6748
rect 35420 6638 35422 6690
rect 35474 6638 35476 6690
rect 35420 6626 35476 6638
rect 35756 6580 35812 6590
rect 35756 6244 35812 6524
rect 35756 6178 35812 6188
rect 35756 5908 35812 5918
rect 35868 5908 35924 6748
rect 35980 6738 36036 6748
rect 36876 6804 36932 7310
rect 36988 7252 37044 7422
rect 36988 7186 37044 7196
rect 37100 7476 37156 8092
rect 37436 8036 37492 8046
rect 37436 7942 37492 7980
rect 36876 6738 36932 6748
rect 36316 6692 36372 6702
rect 36316 6598 36372 6636
rect 37100 6690 37156 7420
rect 37212 7588 37268 7598
rect 37212 6916 37268 7532
rect 37548 7252 37604 9662
rect 37660 10164 37716 10174
rect 37660 9154 37716 10108
rect 37996 9828 38052 9838
rect 37996 9734 38052 9772
rect 37660 9102 37662 9154
rect 37714 9102 37716 9154
rect 37660 9090 37716 9102
rect 37772 9492 37828 9502
rect 37772 9044 37828 9436
rect 37884 9268 37940 9278
rect 37884 9266 38164 9268
rect 37884 9214 37886 9266
rect 37938 9214 38164 9266
rect 37884 9212 38164 9214
rect 37884 9202 37940 9212
rect 37884 9044 37940 9054
rect 37772 9042 37940 9044
rect 37772 8990 37886 9042
rect 37938 8990 37940 9042
rect 37772 8988 37940 8990
rect 37884 8978 37940 8988
rect 37772 8260 37828 8270
rect 37772 8166 37828 8204
rect 37996 8260 38052 8270
rect 37996 8166 38052 8204
rect 38108 7476 38164 9212
rect 38220 9042 38276 10334
rect 38220 8990 38222 9042
rect 38274 8990 38276 9042
rect 38220 7812 38276 8990
rect 38332 8596 38388 11788
rect 38556 12852 38612 12862
rect 38444 11170 38500 11182
rect 38444 11118 38446 11170
rect 38498 11118 38500 11170
rect 38444 11060 38500 11118
rect 38444 10994 38500 11004
rect 38556 10836 38612 12796
rect 38668 12068 38724 13468
rect 39004 13076 39060 13086
rect 39452 13076 39508 13580
rect 39564 13300 39620 13694
rect 39788 13746 39844 14140
rect 39788 13694 39790 13746
rect 39842 13694 39844 13746
rect 39564 13234 39620 13244
rect 39676 13524 39732 13534
rect 39060 13020 39172 13076
rect 39452 13020 39620 13076
rect 39004 13010 39060 13020
rect 39004 12404 39060 12414
rect 39004 12290 39060 12348
rect 39004 12238 39006 12290
rect 39058 12238 39060 12290
rect 39004 12226 39060 12238
rect 38668 12012 39060 12068
rect 39004 11506 39060 12012
rect 39004 11454 39006 11506
rect 39058 11454 39060 11506
rect 39004 11442 39060 11454
rect 38332 8530 38388 8540
rect 38444 10780 38612 10836
rect 38444 8372 38500 10780
rect 38892 10724 38948 10734
rect 38556 10722 38948 10724
rect 38556 10670 38894 10722
rect 38946 10670 38948 10722
rect 38556 10668 38948 10670
rect 38556 10164 38612 10668
rect 38892 10658 38948 10668
rect 38556 9154 38612 10108
rect 38668 10386 38724 10398
rect 38668 10334 38670 10386
rect 38722 10334 38724 10386
rect 38668 9716 38724 10334
rect 38668 9650 38724 9660
rect 39116 9380 39172 13020
rect 39228 10610 39284 10622
rect 39228 10558 39230 10610
rect 39282 10558 39284 10610
rect 39228 10500 39284 10558
rect 39228 10434 39284 10444
rect 39564 9714 39620 13020
rect 39676 11956 39732 13468
rect 39788 13076 39844 13694
rect 39788 13010 39844 13020
rect 39788 12180 39844 12190
rect 40124 12180 40180 16828
rect 40236 15540 40292 17052
rect 40236 15474 40292 15484
rect 40236 13748 40292 13758
rect 40236 13654 40292 13692
rect 40460 12964 40516 21980
rect 40908 21924 40964 23884
rect 41244 23828 41300 24780
rect 41356 24724 41412 26852
rect 41916 26180 41972 26190
rect 41916 26086 41972 26124
rect 42140 26180 42196 26190
rect 42140 26086 42196 26124
rect 42140 25844 42196 25854
rect 42140 25508 42196 25788
rect 41916 25394 41972 25406
rect 41916 25342 41918 25394
rect 41970 25342 41972 25394
rect 41580 25284 41636 25294
rect 41356 24658 41412 24668
rect 41468 24722 41524 24734
rect 41468 24670 41470 24722
rect 41522 24670 41524 24722
rect 41132 23714 41188 23726
rect 41132 23662 41134 23714
rect 41186 23662 41188 23714
rect 41132 23604 41188 23662
rect 41132 23538 41188 23548
rect 40572 21868 40964 21924
rect 41020 23154 41076 23166
rect 41020 23102 41022 23154
rect 41074 23102 41076 23154
rect 41020 21924 41076 23102
rect 41132 22484 41188 22494
rect 41132 22390 41188 22428
rect 40572 14084 40628 21868
rect 41020 21858 41076 21868
rect 41132 21700 41188 21710
rect 41244 21700 41300 23772
rect 41356 23716 41412 23726
rect 41468 23716 41524 24670
rect 41580 23938 41636 25228
rect 41580 23886 41582 23938
rect 41634 23886 41636 23938
rect 41580 23874 41636 23886
rect 41916 25172 41972 25342
rect 41412 23660 41524 23716
rect 41356 23650 41412 23660
rect 41132 21698 41300 21700
rect 41132 21646 41134 21698
rect 41186 21646 41300 21698
rect 41132 21644 41300 21646
rect 41580 23604 41636 23614
rect 40908 21476 40964 21486
rect 40908 21382 40964 21420
rect 41020 19908 41076 19918
rect 40908 19906 41076 19908
rect 40908 19854 41022 19906
rect 41074 19854 41076 19906
rect 40908 19852 41076 19854
rect 40908 18450 40964 19852
rect 41020 19842 41076 19852
rect 41132 19684 41188 21644
rect 41244 21364 41300 21374
rect 41244 21362 41412 21364
rect 41244 21310 41246 21362
rect 41298 21310 41412 21362
rect 41244 21308 41412 21310
rect 41244 21298 41300 21308
rect 41356 20914 41412 21308
rect 41356 20862 41358 20914
rect 41410 20862 41412 20914
rect 41356 20850 41412 20862
rect 41580 20692 41636 23548
rect 41916 23604 41972 25116
rect 41916 23538 41972 23548
rect 42140 24050 42196 25452
rect 42252 24948 42308 26852
rect 42364 26404 42420 26414
rect 42364 26310 42420 26348
rect 42476 26180 42532 26190
rect 42588 26180 42644 27694
rect 42812 27188 42868 28366
rect 42812 27122 42868 27132
rect 43148 26964 43204 28476
rect 43260 28308 43316 28588
rect 43260 28242 43316 28252
rect 43036 26908 43204 26964
rect 42924 26852 43092 26908
rect 42812 26404 42868 26414
rect 42924 26404 42980 26852
rect 42812 26402 42980 26404
rect 42812 26350 42814 26402
rect 42866 26350 42980 26402
rect 42812 26348 42980 26350
rect 43260 26404 43316 26414
rect 42812 26338 42868 26348
rect 43260 26290 43316 26348
rect 43260 26238 43262 26290
rect 43314 26238 43316 26290
rect 43260 26226 43316 26238
rect 42476 26178 42644 26180
rect 42476 26126 42478 26178
rect 42530 26126 42644 26178
rect 42476 26124 42644 26126
rect 42476 26114 42532 26124
rect 42252 24892 42420 24948
rect 42252 24724 42308 24734
rect 42252 24630 42308 24668
rect 42364 24164 42420 24892
rect 42140 23998 42142 24050
rect 42194 23998 42196 24050
rect 41692 23044 41748 23054
rect 41692 22950 41748 22988
rect 41916 21924 41972 21934
rect 40908 18398 40910 18450
rect 40962 18398 40964 18450
rect 40908 17668 40964 18398
rect 40908 17602 40964 17612
rect 41020 19628 41188 19684
rect 41244 20636 41636 20692
rect 41692 21474 41748 21486
rect 41692 21422 41694 21474
rect 41746 21422 41748 21474
rect 41692 20692 41748 21422
rect 41804 21364 41860 21374
rect 41804 21270 41860 21308
rect 41916 20804 41972 21868
rect 42140 21812 42196 23998
rect 42252 24108 42420 24164
rect 43036 24610 43092 24622
rect 43036 24558 43038 24610
rect 43090 24558 43092 24610
rect 43036 24164 43092 24558
rect 43148 24164 43204 24174
rect 43036 24162 43204 24164
rect 43036 24110 43150 24162
rect 43202 24110 43204 24162
rect 43036 24108 43204 24110
rect 42252 22484 42308 24108
rect 43148 24098 43204 24108
rect 42700 23938 42756 23950
rect 42700 23886 42702 23938
rect 42754 23886 42756 23938
rect 42476 23716 42532 23726
rect 42476 23622 42532 23660
rect 42700 23604 42756 23886
rect 43148 23938 43204 23950
rect 43148 23886 43150 23938
rect 43202 23886 43204 23938
rect 43148 23828 43204 23886
rect 43372 23940 43428 29148
rect 43484 28756 43540 30158
rect 43484 28690 43540 28700
rect 43596 28980 43652 28990
rect 43596 28530 43652 28924
rect 43596 28478 43598 28530
rect 43650 28478 43652 28530
rect 43596 28466 43652 28478
rect 43708 28308 43764 30492
rect 43932 30324 43988 30492
rect 43484 28252 43764 28308
rect 43820 30212 43876 30222
rect 43484 25618 43540 28252
rect 43708 27188 43764 27198
rect 43708 26178 43764 27132
rect 43708 26126 43710 26178
rect 43762 26126 43764 26178
rect 43708 26114 43764 26126
rect 43484 25566 43486 25618
rect 43538 25566 43540 25618
rect 43484 25554 43540 25566
rect 43820 25620 43876 30156
rect 43932 30210 43988 30268
rect 44492 30212 44548 31276
rect 44828 31220 44884 31276
rect 45052 31220 45108 35084
rect 45276 34916 45332 34926
rect 45388 34916 45444 35196
rect 45724 35028 45780 36206
rect 45948 36260 46004 36270
rect 46004 36204 46116 36260
rect 45948 36166 46004 36204
rect 46060 35810 46116 36204
rect 46396 35924 46452 38332
rect 46620 36482 46676 42476
rect 46844 38164 46900 44828
rect 47068 43652 47124 43662
rect 46956 42196 47012 42206
rect 46956 40626 47012 42140
rect 47068 41410 47124 43596
rect 47292 41972 47348 45948
rect 47964 45890 48020 45902
rect 47964 45838 47966 45890
rect 48018 45838 48020 45890
rect 47404 45668 47460 45678
rect 47404 45574 47460 45612
rect 47404 45220 47460 45230
rect 47404 45126 47460 45164
rect 47740 45108 47796 45118
rect 47740 44210 47796 45052
rect 47740 44158 47742 44210
rect 47794 44158 47796 44210
rect 47740 44146 47796 44158
rect 47404 43428 47460 43438
rect 47404 43334 47460 43372
rect 47852 42532 47908 42542
rect 47740 42530 47908 42532
rect 47740 42478 47854 42530
rect 47906 42478 47908 42530
rect 47740 42476 47908 42478
rect 47404 41972 47460 41982
rect 47292 41970 47460 41972
rect 47292 41918 47406 41970
rect 47458 41918 47460 41970
rect 47292 41916 47460 41918
rect 47404 41906 47460 41916
rect 47516 41972 47572 41982
rect 47068 41358 47070 41410
rect 47122 41358 47124 41410
rect 47068 41346 47124 41358
rect 46956 40574 46958 40626
rect 47010 40574 47012 40626
rect 46956 40562 47012 40574
rect 47516 40628 47572 41916
rect 47628 40628 47684 40638
rect 47516 40626 47684 40628
rect 47516 40574 47630 40626
rect 47682 40574 47684 40626
rect 47516 40572 47684 40574
rect 47628 40562 47684 40572
rect 47404 40516 47460 40526
rect 47180 40514 47460 40516
rect 47180 40462 47406 40514
rect 47458 40462 47460 40514
rect 47180 40460 47460 40462
rect 47068 40404 47124 40414
rect 47068 40310 47124 40348
rect 47180 40180 47236 40460
rect 47404 40450 47460 40460
rect 46956 40124 47236 40180
rect 47516 40402 47572 40414
rect 47516 40350 47518 40402
rect 47570 40350 47572 40402
rect 46956 38388 47012 40124
rect 47404 39506 47460 39518
rect 47404 39454 47406 39506
rect 47458 39454 47460 39506
rect 47404 39172 47460 39454
rect 47404 39106 47460 39116
rect 46956 38322 47012 38332
rect 47404 38722 47460 38734
rect 47404 38670 47406 38722
rect 47458 38670 47460 38722
rect 47404 38164 47460 38670
rect 46844 38108 47012 38164
rect 46844 37940 46900 37950
rect 46732 37828 46788 37838
rect 46732 37734 46788 37772
rect 46844 36706 46900 37884
rect 46844 36654 46846 36706
rect 46898 36654 46900 36706
rect 46844 36642 46900 36654
rect 46620 36430 46622 36482
rect 46674 36430 46676 36482
rect 46620 36418 46676 36430
rect 46396 35858 46452 35868
rect 46060 35758 46062 35810
rect 46114 35758 46116 35810
rect 46060 35746 46116 35758
rect 45276 34914 45444 34916
rect 45276 34862 45278 34914
rect 45330 34862 45444 34914
rect 45276 34860 45444 34862
rect 45612 34972 45780 35028
rect 45276 34692 45332 34860
rect 45164 34132 45220 34142
rect 45276 34132 45332 34636
rect 45164 34130 45332 34132
rect 45164 34078 45166 34130
rect 45218 34078 45332 34130
rect 45164 34076 45332 34078
rect 45164 33124 45220 34076
rect 45388 33124 45444 33134
rect 45164 33122 45444 33124
rect 45164 33070 45390 33122
rect 45442 33070 45444 33122
rect 45164 33068 45444 33070
rect 45388 32564 45444 33068
rect 45276 32562 45444 32564
rect 45276 32510 45390 32562
rect 45442 32510 45444 32562
rect 45276 32508 45444 32510
rect 45164 31892 45220 31902
rect 45164 31666 45220 31836
rect 45276 31780 45332 32508
rect 45388 32498 45444 32508
rect 45612 32004 45668 34972
rect 45724 34804 45780 34814
rect 46060 34804 46116 34814
rect 45724 34354 45780 34748
rect 45724 34302 45726 34354
rect 45778 34302 45780 34354
rect 45724 33348 45780 34302
rect 45836 34802 46116 34804
rect 45836 34750 46062 34802
rect 46114 34750 46116 34802
rect 45836 34748 46116 34750
rect 45836 34354 45892 34748
rect 46060 34738 46116 34748
rect 45836 34302 45838 34354
rect 45890 34302 45892 34354
rect 45836 34290 45892 34302
rect 45948 34132 46004 34142
rect 46284 34132 46340 34142
rect 45948 34130 46340 34132
rect 45948 34078 45950 34130
rect 46002 34078 46286 34130
rect 46338 34078 46340 34130
rect 45948 34076 46340 34078
rect 45948 34066 46004 34076
rect 46284 34066 46340 34076
rect 46620 34018 46676 34030
rect 46620 33966 46622 34018
rect 46674 33966 46676 34018
rect 45836 33348 45892 33358
rect 45724 33346 45892 33348
rect 45724 33294 45838 33346
rect 45890 33294 45892 33346
rect 45724 33292 45892 33294
rect 45724 32004 45780 32014
rect 45612 32002 45780 32004
rect 45612 31950 45726 32002
rect 45778 31950 45780 32002
rect 45612 31948 45780 31950
rect 45724 31938 45780 31948
rect 45836 32004 45892 33292
rect 46172 33236 46228 33246
rect 46172 33142 46228 33180
rect 46060 33122 46116 33134
rect 46508 33124 46564 33134
rect 46060 33070 46062 33122
rect 46114 33070 46116 33122
rect 46060 32674 46116 33070
rect 46060 32622 46062 32674
rect 46114 32622 46116 32674
rect 46060 32610 46116 32622
rect 46284 33122 46564 33124
rect 46284 33070 46510 33122
rect 46562 33070 46564 33122
rect 46284 33068 46564 33070
rect 45836 31948 46116 32004
rect 45836 31892 45892 31948
rect 45836 31826 45892 31836
rect 45276 31714 45332 31724
rect 45948 31778 46004 31790
rect 45948 31726 45950 31778
rect 46002 31726 46004 31778
rect 45164 31614 45166 31666
rect 45218 31614 45220 31666
rect 45164 31602 45220 31614
rect 45612 31668 45668 31678
rect 45612 31574 45668 31612
rect 44828 31164 45108 31220
rect 45612 31444 45668 31454
rect 44716 31108 44772 31118
rect 44716 31106 44996 31108
rect 44716 31054 44718 31106
rect 44770 31054 44996 31106
rect 44716 31052 44996 31054
rect 44716 31042 44772 31052
rect 43932 30158 43934 30210
rect 43986 30158 43988 30210
rect 43932 30146 43988 30158
rect 44044 30156 44548 30212
rect 44828 30882 44884 30894
rect 44828 30830 44830 30882
rect 44882 30830 44884 30882
rect 44044 29316 44100 30156
rect 44828 30100 44884 30830
rect 44940 30212 44996 31052
rect 45612 31106 45668 31388
rect 45948 31108 46004 31726
rect 45612 31054 45614 31106
rect 45666 31054 45668 31106
rect 45612 31042 45668 31054
rect 45836 31106 46004 31108
rect 45836 31054 45950 31106
rect 46002 31054 46004 31106
rect 45836 31052 46004 31054
rect 45052 30996 45108 31006
rect 45052 30902 45108 30940
rect 45276 30994 45332 31006
rect 45276 30942 45278 30994
rect 45330 30942 45332 30994
rect 44940 30146 44996 30156
rect 45164 30324 45220 30334
rect 45164 30210 45220 30268
rect 45276 30322 45332 30942
rect 45276 30270 45278 30322
rect 45330 30270 45332 30322
rect 45276 30258 45332 30270
rect 45836 30996 45892 31052
rect 45948 31042 46004 31052
rect 45164 30158 45166 30210
rect 45218 30158 45220 30210
rect 45164 30146 45220 30158
rect 45612 30212 45668 30222
rect 45612 30118 45668 30156
rect 44156 30044 44884 30100
rect 45052 30098 45108 30110
rect 45052 30046 45054 30098
rect 45106 30046 45108 30098
rect 44156 29538 44212 30044
rect 44156 29486 44158 29538
rect 44210 29486 44212 29538
rect 44156 29474 44212 29486
rect 45052 29988 45108 30046
rect 44492 29316 44548 29326
rect 44044 29260 44212 29316
rect 44044 28868 44100 28878
rect 43932 28756 43988 28766
rect 43932 28662 43988 28700
rect 44044 28642 44100 28812
rect 44044 28590 44046 28642
rect 44098 28590 44100 28642
rect 44044 28578 44100 28590
rect 43932 25620 43988 25630
rect 43820 25618 43988 25620
rect 43820 25566 43934 25618
rect 43986 25566 43988 25618
rect 43820 25564 43988 25566
rect 43932 25554 43988 25564
rect 43484 24500 43540 24510
rect 43484 24162 43540 24444
rect 43484 24110 43486 24162
rect 43538 24110 43540 24162
rect 43484 24098 43540 24110
rect 43372 23884 43540 23940
rect 43148 23762 43204 23772
rect 42700 23538 42756 23548
rect 42812 23716 42868 23726
rect 42252 22148 42308 22428
rect 42252 22082 42308 22092
rect 42252 21812 42308 21822
rect 42140 21810 42644 21812
rect 42140 21758 42254 21810
rect 42306 21758 42644 21810
rect 42140 21756 42644 21758
rect 42252 21746 42308 21756
rect 42476 20914 42532 20926
rect 42476 20862 42478 20914
rect 42530 20862 42532 20914
rect 42028 20804 42084 20814
rect 41916 20802 42084 20804
rect 41916 20750 42030 20802
rect 42082 20750 42084 20802
rect 41916 20748 42084 20750
rect 40684 17556 40740 17566
rect 40684 17554 40852 17556
rect 40684 17502 40686 17554
rect 40738 17502 40852 17554
rect 40684 17500 40852 17502
rect 40684 17490 40740 17500
rect 40796 14308 40852 17500
rect 40908 16884 40964 16894
rect 40908 16790 40964 16828
rect 41020 15428 41076 19628
rect 41020 15362 41076 15372
rect 41132 18452 41188 18462
rect 41132 15538 41188 18396
rect 41244 15988 41300 20636
rect 41692 20626 41748 20636
rect 41804 20020 41860 20030
rect 42028 20020 42084 20748
rect 42476 20130 42532 20862
rect 42588 20690 42644 21756
rect 42812 21588 42868 23660
rect 43148 22820 43204 22830
rect 43148 22370 43204 22764
rect 43148 22318 43150 22370
rect 43202 22318 43204 22370
rect 43148 22306 43204 22318
rect 43372 22596 43428 22606
rect 43372 22370 43428 22540
rect 43372 22318 43374 22370
rect 43426 22318 43428 22370
rect 43372 22306 43428 22318
rect 42588 20638 42590 20690
rect 42642 20638 42644 20690
rect 42588 20626 42644 20638
rect 42700 21532 42868 21588
rect 43260 21586 43316 21598
rect 43260 21534 43262 21586
rect 43314 21534 43316 21586
rect 42476 20078 42478 20130
rect 42530 20078 42532 20130
rect 42476 20066 42532 20078
rect 41804 20018 42084 20020
rect 41804 19966 41806 20018
rect 41858 19966 42084 20018
rect 41804 19964 42084 19966
rect 41580 18340 41636 18350
rect 41804 18340 41860 19964
rect 42364 19122 42420 19134
rect 42364 19070 42366 19122
rect 42418 19070 42420 19122
rect 42028 18340 42084 18350
rect 41804 18284 42028 18340
rect 41356 16210 41412 16222
rect 41356 16158 41358 16210
rect 41410 16158 41412 16210
rect 41356 16100 41412 16158
rect 41580 16100 41636 18284
rect 41916 17668 41972 17678
rect 41916 17574 41972 17612
rect 42028 16884 42084 18284
rect 42364 17780 42420 19070
rect 42700 18004 42756 21532
rect 42812 21364 42868 21374
rect 42812 21026 42868 21308
rect 42812 20974 42814 21026
rect 42866 20974 42868 21026
rect 42812 20962 42868 20974
rect 43036 19236 43092 19246
rect 43260 19236 43316 21534
rect 43036 19234 43316 19236
rect 43036 19182 43038 19234
rect 43090 19182 43316 19234
rect 43036 19180 43316 19182
rect 42924 19012 42980 19022
rect 42924 18004 42980 18956
rect 43036 18340 43092 19180
rect 43484 19124 43540 23884
rect 44156 23156 44212 29260
rect 44492 28084 44548 29260
rect 44716 28868 44772 28878
rect 44268 27188 44324 27198
rect 44268 27094 44324 27132
rect 44380 25620 44436 25630
rect 44492 25620 44548 28028
rect 44604 28812 44716 28868
rect 44604 26908 44660 28812
rect 44716 28802 44772 28812
rect 44940 28644 44996 28654
rect 45052 28644 45108 29932
rect 45388 29988 45444 29998
rect 45388 29986 45556 29988
rect 45388 29934 45390 29986
rect 45442 29934 45556 29986
rect 45388 29932 45556 29934
rect 45388 29922 45444 29932
rect 44996 28588 45108 28644
rect 45388 29540 45444 29550
rect 45388 28642 45444 29484
rect 45500 29428 45556 29932
rect 45836 29428 45892 30940
rect 46060 30434 46116 31948
rect 46172 31780 46228 31790
rect 46284 31780 46340 33068
rect 46508 33058 46564 33068
rect 46620 33124 46676 33966
rect 46844 33572 46900 33582
rect 46620 31892 46676 33068
rect 46172 31778 46340 31780
rect 46172 31726 46174 31778
rect 46226 31726 46340 31778
rect 46172 31724 46340 31726
rect 46396 31836 46676 31892
rect 46732 33570 46900 33572
rect 46732 33518 46846 33570
rect 46898 33518 46900 33570
rect 46732 33516 46900 33518
rect 46732 33348 46788 33516
rect 46844 33506 46900 33516
rect 46172 31714 46228 31724
rect 46172 31556 46228 31566
rect 46172 31218 46228 31500
rect 46396 31332 46452 31836
rect 46732 31778 46788 33292
rect 46956 33236 47012 38108
rect 47404 38098 47460 38108
rect 47516 37940 47572 40350
rect 47628 40404 47684 40414
rect 47628 38276 47684 40348
rect 47740 38668 47796 42476
rect 47852 42466 47908 42476
rect 47964 41860 48020 45838
rect 48188 45106 48244 45118
rect 48188 45054 48190 45106
rect 48242 45054 48244 45106
rect 48076 44212 48132 44222
rect 48076 44118 48132 44156
rect 48188 43540 48244 45054
rect 47964 41794 48020 41804
rect 48076 43538 48244 43540
rect 48076 43486 48190 43538
rect 48242 43486 48244 43538
rect 48076 43484 48244 43486
rect 48076 41970 48132 43484
rect 48188 43474 48244 43484
rect 48188 42644 48244 42654
rect 48188 42550 48244 42588
rect 48412 42644 48468 47068
rect 48412 42578 48468 42588
rect 48076 41918 48078 41970
rect 48130 41918 48132 41970
rect 47852 40516 47908 40526
rect 47852 40422 47908 40460
rect 48076 39618 48132 41918
rect 48076 39566 48078 39618
rect 48130 39566 48132 39618
rect 48076 38834 48132 39566
rect 48076 38782 48078 38834
rect 48130 38782 48132 38834
rect 47740 38612 47908 38668
rect 47628 38220 47796 38276
rect 47628 38052 47684 38062
rect 47628 37958 47684 37996
rect 47068 37884 47572 37940
rect 47068 37378 47124 37884
rect 47740 37716 47796 38220
rect 47068 37326 47070 37378
rect 47122 37326 47124 37378
rect 47068 37314 47124 37326
rect 47628 37660 47796 37716
rect 47404 36932 47460 36942
rect 47404 36482 47460 36876
rect 47628 36594 47684 37660
rect 47740 37492 47796 37502
rect 47740 37266 47796 37436
rect 47740 37214 47742 37266
rect 47794 37214 47796 37266
rect 47740 37044 47796 37214
rect 47740 36978 47796 36988
rect 47628 36542 47630 36594
rect 47682 36542 47684 36594
rect 47628 36530 47684 36542
rect 47404 36430 47406 36482
rect 47458 36430 47460 36482
rect 47404 36418 47460 36430
rect 47852 36372 47908 38612
rect 48076 37716 48132 38782
rect 48188 37826 48244 37838
rect 48188 37774 48190 37826
rect 48242 37774 48244 37826
rect 48188 37716 48244 37774
rect 48188 37660 48356 37716
rect 48076 37650 48132 37660
rect 48300 37268 48356 37660
rect 48300 37202 48356 37212
rect 47852 36316 48468 36372
rect 48188 35588 48244 35598
rect 48188 35494 48244 35532
rect 47180 35028 47236 35038
rect 47180 34130 47236 34972
rect 48188 35028 48244 35038
rect 48188 34934 48244 34972
rect 47852 34692 47908 34702
rect 47852 34354 47908 34636
rect 47852 34302 47854 34354
rect 47906 34302 47908 34354
rect 47852 34290 47908 34302
rect 47180 34078 47182 34130
rect 47234 34078 47236 34130
rect 47180 33460 47236 34078
rect 47180 33404 47684 33460
rect 46732 31726 46734 31778
rect 46786 31726 46788 31778
rect 46732 31714 46788 31726
rect 46844 33180 47012 33236
rect 47068 33348 47124 33358
rect 47180 33348 47236 33404
rect 47068 33346 47236 33348
rect 47068 33294 47070 33346
rect 47122 33294 47236 33346
rect 47068 33292 47236 33294
rect 47628 33346 47684 33404
rect 47628 33294 47630 33346
rect 47682 33294 47684 33346
rect 46172 31166 46174 31218
rect 46226 31166 46228 31218
rect 46172 31154 46228 31166
rect 46284 31276 46452 31332
rect 46508 31666 46564 31678
rect 46508 31614 46510 31666
rect 46562 31614 46564 31666
rect 46060 30382 46062 30434
rect 46114 30382 46116 30434
rect 46060 30370 46116 30382
rect 46172 30996 46228 31006
rect 46060 30212 46116 30222
rect 45500 29372 45836 29428
rect 45836 29362 45892 29372
rect 45948 30098 46004 30110
rect 45948 30046 45950 30098
rect 46002 30046 46004 30098
rect 45948 28756 46004 30046
rect 46060 29540 46116 30156
rect 46060 29474 46116 29484
rect 46172 28868 46228 30940
rect 46284 30436 46340 31276
rect 46396 31108 46452 31118
rect 46396 31014 46452 31052
rect 46508 30994 46564 31614
rect 46620 31444 46676 31454
rect 46676 31388 46788 31444
rect 46620 31378 46676 31388
rect 46508 30942 46510 30994
rect 46562 30942 46564 30994
rect 46396 30436 46452 30446
rect 46284 30380 46396 30436
rect 46396 30342 46452 30380
rect 46508 30324 46564 30942
rect 46508 30258 46564 30268
rect 46284 30212 46340 30222
rect 46732 30212 46788 31388
rect 46844 30436 46900 33180
rect 47068 33124 47124 33292
rect 47628 33282 47684 33294
rect 47852 33348 47908 33358
rect 47908 33292 48244 33348
rect 47852 33254 47908 33292
rect 47404 33234 47460 33246
rect 47404 33182 47406 33234
rect 47458 33182 47460 33234
rect 46956 33068 47124 33124
rect 47180 33124 47236 33134
rect 47404 33124 47460 33182
rect 47516 33236 47572 33246
rect 47516 33142 47572 33180
rect 47236 33068 47460 33124
rect 46956 31666 47012 33068
rect 47180 33058 47236 33068
rect 48188 32450 48244 33292
rect 48188 32398 48190 32450
rect 48242 32398 48244 32450
rect 48188 32386 48244 32398
rect 48076 32340 48132 32350
rect 46956 31614 46958 31666
rect 47010 31614 47012 31666
rect 46956 31602 47012 31614
rect 47628 31778 47684 31790
rect 47628 31726 47630 31778
rect 47682 31726 47684 31778
rect 47404 31108 47460 31118
rect 47404 31014 47460 31052
rect 46956 30882 47012 30894
rect 46956 30830 46958 30882
rect 47010 30830 47012 30882
rect 46956 30772 47012 30830
rect 46956 30706 47012 30716
rect 47628 30660 47684 31726
rect 48076 31780 48132 32284
rect 48076 31778 48356 31780
rect 48076 31726 48078 31778
rect 48130 31726 48356 31778
rect 48076 31724 48356 31726
rect 48076 31714 48132 31724
rect 48300 31218 48356 31724
rect 48300 31166 48302 31218
rect 48354 31166 48356 31218
rect 48300 31154 48356 31166
rect 47628 30594 47684 30604
rect 47628 30436 47684 30446
rect 46844 30380 47012 30436
rect 46844 30212 46900 30222
rect 46284 30210 46452 30212
rect 46284 30158 46286 30210
rect 46338 30158 46452 30210
rect 46284 30156 46452 30158
rect 46732 30210 46900 30212
rect 46732 30158 46846 30210
rect 46898 30158 46900 30210
rect 46732 30156 46900 30158
rect 46284 30146 46340 30156
rect 46396 29988 46452 30156
rect 46844 30146 46900 30156
rect 46396 29932 46900 29988
rect 46844 29650 46900 29932
rect 46956 29764 47012 30380
rect 47068 30212 47124 30222
rect 47068 30118 47124 30156
rect 47628 30210 47684 30380
rect 47628 30158 47630 30210
rect 47682 30158 47684 30210
rect 47628 30146 47684 30158
rect 47180 30100 47236 30110
rect 47180 30098 47348 30100
rect 47180 30046 47182 30098
rect 47234 30046 47348 30098
rect 47180 30044 47348 30046
rect 47180 30034 47236 30044
rect 46956 29708 47236 29764
rect 46844 29598 46846 29650
rect 46898 29598 46900 29650
rect 46844 29586 46900 29598
rect 46284 29540 46340 29550
rect 46284 29314 46340 29484
rect 46620 29540 46676 29550
rect 46620 29426 46676 29484
rect 46620 29374 46622 29426
rect 46674 29374 46676 29426
rect 46620 29362 46676 29374
rect 47068 29428 47124 29438
rect 47068 29334 47124 29372
rect 46284 29262 46286 29314
rect 46338 29262 46340 29314
rect 46284 29250 46340 29262
rect 46172 28802 46228 28812
rect 46060 28756 46116 28766
rect 45948 28754 46116 28756
rect 45948 28702 46062 28754
rect 46114 28702 46116 28754
rect 45948 28700 46116 28702
rect 46060 28690 46116 28700
rect 45388 28590 45390 28642
rect 45442 28590 45444 28642
rect 44940 28550 44996 28588
rect 44716 27746 44772 27758
rect 44716 27694 44718 27746
rect 44770 27694 44772 27746
rect 44716 27300 44772 27694
rect 45276 27636 45332 27646
rect 44716 27244 45108 27300
rect 44940 26962 44996 26974
rect 44940 26910 44942 26962
rect 44994 26910 44996 26962
rect 44940 26908 44996 26910
rect 44604 26852 44996 26908
rect 44380 25618 44548 25620
rect 44380 25566 44382 25618
rect 44434 25566 44548 25618
rect 44380 25564 44548 25566
rect 44380 25554 44436 25564
rect 44380 23828 44436 23838
rect 44380 23378 44436 23772
rect 44828 23716 44884 26852
rect 45052 26404 45108 27244
rect 45052 26338 45108 26348
rect 44940 25620 44996 25630
rect 44940 25394 44996 25564
rect 45052 25508 45108 25518
rect 45052 25414 45108 25452
rect 45164 25506 45220 25518
rect 45164 25454 45166 25506
rect 45218 25454 45220 25506
rect 44940 25342 44942 25394
rect 44994 25342 44996 25394
rect 44940 25330 44996 25342
rect 45164 25396 45220 25454
rect 45276 25396 45332 27580
rect 45164 25340 45276 25396
rect 45276 25330 45332 25340
rect 45388 27074 45444 28590
rect 47180 28532 47236 29708
rect 47292 29426 47348 30044
rect 48076 29988 48132 29998
rect 48076 29894 48132 29932
rect 47292 29374 47294 29426
rect 47346 29374 47348 29426
rect 47292 29204 47348 29374
rect 47852 29316 47908 29326
rect 48188 29316 48244 29326
rect 47852 29314 48020 29316
rect 47852 29262 47854 29314
rect 47906 29262 48020 29314
rect 47852 29260 48020 29262
rect 47852 29250 47908 29260
rect 47404 29204 47460 29214
rect 47292 29202 47460 29204
rect 47292 29150 47406 29202
rect 47458 29150 47460 29202
rect 47292 29148 47460 29150
rect 47404 29138 47460 29148
rect 47180 28476 47572 28532
rect 47516 28082 47572 28476
rect 47516 28030 47518 28082
rect 47570 28030 47572 28082
rect 45836 27860 45892 27870
rect 45836 27766 45892 27804
rect 46396 27858 46452 27870
rect 46396 27806 46398 27858
rect 46450 27806 46452 27858
rect 45500 27636 45556 27646
rect 45500 27542 45556 27580
rect 45612 27634 45668 27646
rect 45612 27582 45614 27634
rect 45666 27582 45668 27634
rect 45388 27022 45390 27074
rect 45442 27022 45444 27074
rect 45164 24724 45220 24734
rect 45164 24610 45220 24668
rect 45164 24558 45166 24610
rect 45218 24558 45220 24610
rect 45052 24052 45108 24062
rect 45052 23958 45108 23996
rect 44828 23650 44884 23660
rect 44380 23326 44382 23378
rect 44434 23326 44436 23378
rect 44380 23314 44436 23326
rect 44940 23268 44996 23278
rect 44940 23174 44996 23212
rect 44156 23090 44212 23100
rect 45164 23154 45220 24558
rect 45388 23938 45444 27022
rect 45388 23886 45390 23938
rect 45442 23886 45444 23938
rect 45388 23874 45444 23886
rect 45500 27412 45556 27422
rect 45500 23380 45556 27356
rect 45612 26908 45668 27582
rect 45948 27636 46004 27646
rect 45948 27634 46116 27636
rect 45948 27582 45950 27634
rect 46002 27582 46116 27634
rect 45948 27580 46116 27582
rect 45948 27570 46004 27580
rect 46060 27186 46116 27580
rect 46060 27134 46062 27186
rect 46114 27134 46116 27186
rect 46060 27122 46116 27134
rect 45612 26852 46004 26908
rect 45836 26740 45892 26750
rect 45612 26404 45668 26414
rect 45612 25506 45668 26348
rect 45612 25454 45614 25506
rect 45666 25454 45668 25506
rect 45612 25442 45668 25454
rect 45836 26292 45892 26684
rect 45836 25732 45892 26236
rect 45948 26068 46004 26852
rect 46396 26740 46452 27806
rect 46396 26674 46452 26684
rect 46508 27858 46564 27870
rect 46508 27806 46510 27858
rect 46562 27806 46564 27858
rect 46508 27188 46564 27806
rect 46508 26404 46564 27132
rect 46620 27858 46676 27870
rect 46620 27806 46622 27858
rect 46674 27806 46676 27858
rect 46620 26908 46676 27806
rect 47516 27860 47572 28030
rect 47068 27636 47124 27646
rect 47068 27542 47124 27580
rect 47068 27188 47124 27198
rect 47068 26908 47124 27132
rect 47516 26908 47572 27804
rect 47852 27970 47908 27982
rect 47852 27918 47854 27970
rect 47906 27918 47908 27970
rect 47852 27412 47908 27918
rect 47964 27860 48020 29260
rect 48188 29222 48244 29260
rect 48076 29202 48132 29214
rect 48076 29150 48078 29202
rect 48130 29150 48132 29202
rect 48076 28756 48132 29150
rect 48188 28756 48244 28766
rect 48076 28754 48244 28756
rect 48076 28702 48190 28754
rect 48242 28702 48244 28754
rect 48076 28700 48244 28702
rect 48188 28690 48244 28700
rect 48188 27860 48244 27870
rect 47964 27858 48244 27860
rect 47964 27806 48190 27858
rect 48242 27806 48244 27858
rect 47964 27804 48244 27806
rect 47852 27346 47908 27356
rect 48188 27412 48244 27804
rect 48188 27346 48244 27356
rect 48188 27188 48244 27198
rect 48188 27094 48244 27132
rect 46620 26852 47124 26908
rect 46732 26514 46788 26526
rect 46732 26462 46734 26514
rect 46786 26462 46788 26514
rect 46172 26348 46676 26404
rect 46172 26290 46228 26348
rect 46172 26238 46174 26290
rect 46226 26238 46228 26290
rect 46172 26226 46228 26238
rect 45948 26012 46452 26068
rect 45836 25394 45892 25676
rect 46396 25618 46452 26012
rect 46396 25566 46398 25618
rect 46450 25566 46452 25618
rect 46396 25554 46452 25566
rect 46508 25732 46564 25742
rect 46508 25506 46564 25676
rect 46508 25454 46510 25506
rect 46562 25454 46564 25506
rect 46508 25442 46564 25454
rect 45836 25342 45838 25394
rect 45890 25342 45892 25394
rect 45836 25330 45892 25342
rect 46284 25394 46340 25406
rect 46284 25342 46286 25394
rect 46338 25342 46340 25394
rect 46060 25284 46116 25294
rect 46284 25284 46340 25342
rect 46620 25284 46676 26348
rect 46284 25228 46676 25284
rect 45948 24724 46004 24734
rect 45612 24500 45668 24510
rect 45612 24406 45668 24444
rect 45388 23324 45556 23380
rect 45948 23380 46004 24668
rect 46060 24050 46116 25228
rect 46732 25172 46788 26462
rect 47068 26404 47124 26852
rect 46844 26402 47124 26404
rect 46844 26350 47070 26402
rect 47122 26350 47124 26402
rect 46844 26348 47124 26350
rect 46844 25506 46900 26348
rect 47068 26338 47124 26348
rect 47404 26852 47572 26908
rect 47404 25844 47460 26852
rect 48188 26292 48244 26302
rect 47404 25778 47460 25788
rect 47516 26290 48244 26292
rect 47516 26238 48190 26290
rect 48242 26238 48244 26290
rect 47516 26236 48244 26238
rect 47292 25620 47348 25630
rect 46844 25454 46846 25506
rect 46898 25454 46900 25506
rect 46844 25442 46900 25454
rect 46956 25618 47348 25620
rect 46956 25566 47294 25618
rect 47346 25566 47348 25618
rect 46956 25564 47348 25566
rect 46732 25106 46788 25116
rect 46956 24948 47012 25564
rect 47292 25554 47348 25564
rect 47516 25620 47572 26236
rect 47628 25844 47684 25854
rect 47628 25730 47684 25788
rect 47628 25678 47630 25730
rect 47682 25678 47684 25730
rect 47628 25666 47684 25678
rect 47404 25508 47460 25518
rect 47404 25414 47460 25452
rect 46060 23998 46062 24050
rect 46114 23998 46116 24050
rect 46060 23986 46116 23998
rect 46396 24946 47012 24948
rect 46396 24894 46958 24946
rect 47010 24894 47012 24946
rect 46396 24892 47012 24894
rect 46396 24610 46452 24892
rect 46956 24882 47012 24892
rect 47180 25396 47236 25406
rect 47180 24724 47236 25340
rect 47292 25284 47348 25294
rect 47292 25190 47348 25228
rect 47292 24724 47348 24734
rect 47180 24722 47348 24724
rect 47180 24670 47294 24722
rect 47346 24670 47348 24722
rect 47180 24668 47348 24670
rect 47292 24658 47348 24668
rect 47516 24722 47572 25564
rect 47516 24670 47518 24722
rect 47570 24670 47572 24722
rect 47516 24658 47572 24670
rect 47628 25172 47684 25182
rect 46396 24558 46398 24610
rect 46450 24558 46452 24610
rect 46060 23380 46116 23390
rect 45948 23378 46116 23380
rect 45948 23326 46062 23378
rect 46114 23326 46116 23378
rect 45948 23324 46116 23326
rect 45164 23102 45166 23154
rect 45218 23102 45220 23154
rect 45164 23090 45220 23102
rect 45276 23156 45332 23166
rect 43820 23042 43876 23054
rect 43820 22990 43822 23042
rect 43874 22990 43876 23042
rect 43820 22820 43876 22990
rect 44268 23044 44324 23054
rect 44268 22950 44324 22988
rect 45052 23042 45108 23054
rect 45052 22990 45054 23042
rect 45106 22990 45108 23042
rect 44156 22932 44212 22942
rect 43820 22754 43876 22764
rect 43932 22930 44212 22932
rect 43932 22878 44158 22930
rect 44210 22878 44212 22930
rect 43932 22876 44212 22878
rect 43932 22596 43988 22876
rect 44156 22866 44212 22876
rect 44156 22596 44212 22606
rect 43596 22540 43988 22596
rect 44044 22540 44156 22596
rect 43596 22482 43652 22540
rect 43596 22430 43598 22482
rect 43650 22430 43652 22482
rect 43596 22418 43652 22430
rect 43932 22372 43988 22382
rect 44044 22372 44100 22540
rect 44156 22530 44212 22540
rect 43932 22370 44100 22372
rect 43932 22318 43934 22370
rect 43986 22318 44100 22370
rect 43932 22316 44100 22318
rect 43932 22306 43988 22316
rect 44268 22260 44324 22270
rect 44828 22260 44884 22270
rect 44268 22258 44884 22260
rect 44268 22206 44270 22258
rect 44322 22206 44830 22258
rect 44882 22206 44884 22258
rect 44268 22204 44884 22206
rect 44268 22194 44324 22204
rect 44828 22194 44884 22204
rect 45052 22258 45108 22990
rect 45052 22206 45054 22258
rect 45106 22206 45108 22258
rect 45052 22194 45108 22206
rect 44044 22148 44100 22158
rect 44044 22054 44100 22092
rect 44940 22146 44996 22158
rect 44940 22094 44942 22146
rect 44994 22094 44996 22146
rect 44940 21812 44996 22094
rect 45276 22036 45332 23100
rect 44044 21756 44996 21812
rect 45052 21980 45332 22036
rect 44044 21698 44100 21756
rect 44044 21646 44046 21698
rect 44098 21646 44100 21698
rect 44044 21634 44100 21646
rect 44044 21476 44100 21486
rect 43932 21364 43988 21374
rect 43932 20020 43988 21308
rect 43932 19458 43988 19964
rect 43932 19406 43934 19458
rect 43986 19406 43988 19458
rect 43932 19394 43988 19406
rect 43708 19348 43764 19358
rect 43708 19254 43764 19292
rect 43036 18274 43092 18284
rect 43260 19068 43540 19124
rect 42924 17948 43092 18004
rect 42700 17938 42756 17948
rect 42924 17780 42980 17790
rect 42364 17778 42980 17780
rect 42364 17726 42926 17778
rect 42978 17726 42980 17778
rect 42364 17724 42980 17726
rect 42924 17714 42980 17724
rect 43036 17780 43092 17948
rect 43036 17666 43092 17724
rect 43036 17614 43038 17666
rect 43090 17614 43092 17666
rect 43036 17602 43092 17614
rect 42028 16818 42084 16828
rect 42812 17554 42868 17566
rect 42812 17502 42814 17554
rect 42866 17502 42868 17554
rect 41692 16770 41748 16782
rect 41692 16718 41694 16770
rect 41746 16718 41748 16770
rect 41692 16212 41748 16718
rect 41804 16212 41860 16222
rect 42700 16212 42756 16222
rect 41692 16210 41860 16212
rect 41692 16158 41806 16210
rect 41858 16158 41860 16210
rect 41692 16156 41860 16158
rect 41804 16146 41860 16156
rect 42364 16210 42756 16212
rect 42364 16158 42702 16210
rect 42754 16158 42756 16210
rect 42364 16156 42756 16158
rect 41356 16044 41524 16100
rect 41580 16044 41748 16100
rect 41244 15932 41412 15988
rect 41132 15486 41134 15538
rect 41186 15486 41188 15538
rect 40908 15314 40964 15326
rect 40908 15262 40910 15314
rect 40962 15262 40964 15314
rect 40908 14532 40964 15262
rect 41132 15148 41188 15486
rect 41244 15764 41300 15774
rect 41244 15426 41300 15708
rect 41244 15374 41246 15426
rect 41298 15374 41300 15426
rect 41244 15362 41300 15374
rect 41356 15428 41412 15932
rect 41468 15652 41524 16044
rect 41692 15986 41748 16044
rect 42364 16098 42420 16156
rect 42700 16146 42756 16156
rect 42364 16046 42366 16098
rect 42418 16046 42420 16098
rect 42364 16034 42420 16046
rect 42588 15988 42644 15998
rect 42812 15988 42868 17502
rect 43148 17556 43204 17566
rect 43036 16548 43092 16558
rect 42924 16100 42980 16110
rect 42924 16006 42980 16044
rect 41692 15934 41694 15986
rect 41746 15934 41748 15986
rect 41692 15922 41748 15934
rect 42476 15986 42868 15988
rect 42476 15934 42590 15986
rect 42642 15934 42868 15986
rect 42476 15932 42868 15934
rect 41916 15876 41972 15886
rect 41916 15782 41972 15820
rect 42476 15876 42532 15932
rect 42588 15922 42644 15932
rect 41468 15596 41860 15652
rect 41580 15428 41636 15438
rect 41356 15426 41636 15428
rect 41356 15374 41582 15426
rect 41634 15374 41636 15426
rect 41356 15372 41636 15374
rect 41580 15362 41636 15372
rect 41692 15428 41748 15438
rect 41692 15148 41748 15372
rect 41804 15314 41860 15596
rect 42476 15538 42532 15820
rect 42476 15486 42478 15538
rect 42530 15486 42532 15538
rect 42476 15474 42532 15486
rect 41804 15262 41806 15314
rect 41858 15262 41860 15314
rect 41804 15250 41860 15262
rect 42812 15316 42868 15326
rect 41132 15092 41412 15148
rect 41356 14642 41412 15092
rect 41356 14590 41358 14642
rect 41410 14590 41412 14642
rect 41356 14578 41412 14590
rect 41580 15092 41748 15148
rect 42140 15204 42196 15242
rect 42812 15222 42868 15260
rect 42140 15138 42196 15148
rect 40908 14466 40964 14476
rect 40908 14308 40964 14318
rect 40796 14252 40908 14308
rect 40572 14018 40628 14028
rect 40908 13524 40964 14252
rect 41020 14084 41076 14094
rect 41020 13970 41076 14028
rect 41020 13918 41022 13970
rect 41074 13918 41076 13970
rect 41020 13906 41076 13918
rect 41580 13970 41636 15092
rect 41580 13918 41582 13970
rect 41634 13918 41636 13970
rect 41580 13906 41636 13918
rect 40908 13458 40964 13468
rect 41692 13634 41748 13646
rect 41692 13582 41694 13634
rect 41746 13582 41748 13634
rect 41020 13300 41076 13310
rect 40684 13076 40740 13086
rect 40684 12982 40740 13020
rect 41020 13076 41076 13244
rect 41692 13076 41748 13582
rect 41020 13074 41300 13076
rect 41020 13022 41022 13074
rect 41074 13022 41300 13074
rect 41020 13020 41300 13022
rect 41020 13010 41076 13020
rect 40460 12898 40516 12908
rect 40348 12628 40404 12638
rect 40348 12402 40404 12572
rect 40348 12350 40350 12402
rect 40402 12350 40404 12402
rect 40348 12338 40404 12350
rect 39788 12178 40180 12180
rect 39788 12126 39790 12178
rect 39842 12126 40180 12178
rect 39788 12124 40180 12126
rect 41244 12178 41300 13020
rect 41692 13010 41748 13020
rect 41804 13522 41860 13534
rect 41804 13470 41806 13522
rect 41858 13470 41860 13522
rect 41244 12126 41246 12178
rect 41298 12126 41300 12178
rect 39788 12114 39844 12124
rect 41244 12114 41300 12126
rect 41468 12628 41524 12638
rect 41132 12068 41188 12078
rect 39676 11900 39844 11956
rect 39564 9662 39566 9714
rect 39618 9662 39620 9714
rect 39564 9650 39620 9662
rect 39676 10610 39732 10622
rect 39676 10558 39678 10610
rect 39730 10558 39732 10610
rect 39676 10500 39732 10558
rect 38892 9324 39172 9380
rect 39676 9602 39732 10444
rect 39788 9828 39844 11900
rect 40572 11732 40628 11742
rect 40572 11506 40628 11676
rect 41132 11732 41188 12012
rect 41132 11666 41188 11676
rect 40572 11454 40574 11506
rect 40626 11454 40628 11506
rect 40572 11442 40628 11454
rect 41468 11508 41524 12572
rect 41804 12292 41860 13470
rect 42812 13412 42868 13422
rect 42812 12964 42868 13356
rect 42812 12404 42868 12908
rect 43036 12852 43092 16492
rect 43148 16098 43204 17500
rect 43148 16046 43150 16098
rect 43202 16046 43204 16098
rect 43148 15540 43204 16046
rect 43148 15474 43204 15484
rect 43148 15314 43204 15326
rect 43148 15262 43150 15314
rect 43202 15262 43204 15314
rect 43148 15204 43204 15262
rect 43148 15138 43204 15148
rect 43260 13972 43316 19068
rect 43820 18452 43876 18490
rect 43820 18386 43876 18396
rect 43820 18228 43876 18238
rect 43372 18226 43876 18228
rect 43372 18174 43822 18226
rect 43874 18174 43876 18226
rect 43372 18172 43876 18174
rect 43372 17890 43428 18172
rect 43820 18162 43876 18172
rect 44044 18004 44100 21420
rect 44380 20916 44436 20926
rect 44380 20822 44436 20860
rect 45052 20914 45108 21980
rect 45388 21812 45444 23324
rect 45836 23266 45892 23278
rect 45836 23214 45838 23266
rect 45890 23214 45892 23266
rect 45276 21756 45444 21812
rect 45500 23156 45556 23166
rect 45836 23156 45892 23214
rect 45500 23154 45892 23156
rect 45500 23102 45502 23154
rect 45554 23102 45892 23154
rect 45500 23100 45892 23102
rect 45500 22370 45556 23100
rect 45948 23044 46004 23324
rect 46060 23314 46116 23324
rect 46396 23268 46452 24558
rect 47180 23268 47236 23278
rect 46396 23154 46452 23212
rect 46956 23212 47180 23268
rect 46732 23156 46788 23166
rect 46396 23102 46398 23154
rect 46450 23102 46452 23154
rect 46396 23090 46452 23102
rect 46620 23100 46732 23156
rect 45836 22988 46004 23044
rect 45724 22930 45780 22942
rect 45724 22878 45726 22930
rect 45778 22878 45780 22930
rect 45724 22596 45780 22878
rect 45724 22530 45780 22540
rect 45500 22318 45502 22370
rect 45554 22318 45556 22370
rect 45276 21252 45332 21756
rect 45276 21186 45332 21196
rect 45388 21588 45444 21598
rect 45388 21028 45444 21532
rect 45500 21476 45556 22318
rect 45724 22372 45780 22382
rect 45836 22372 45892 22988
rect 45948 22820 46004 22830
rect 45948 22594 46004 22764
rect 45948 22542 45950 22594
rect 46002 22542 46004 22594
rect 45948 22530 46004 22542
rect 46620 22594 46676 23100
rect 46732 23062 46788 23100
rect 46956 22820 47012 23212
rect 47180 23174 47236 23212
rect 47516 23268 47572 23278
rect 47404 23044 47460 23054
rect 47404 22950 47460 22988
rect 46620 22542 46622 22594
rect 46674 22542 46676 22594
rect 45724 22370 45892 22372
rect 45724 22318 45726 22370
rect 45778 22318 45892 22370
rect 45724 22316 45892 22318
rect 46620 22372 46676 22542
rect 45724 22306 45780 22316
rect 46396 22146 46452 22158
rect 46396 22094 46398 22146
rect 46450 22094 46452 22146
rect 46396 21700 46452 22094
rect 46620 21810 46676 22316
rect 46844 22764 47012 22820
rect 46844 22258 46900 22764
rect 46844 22206 46846 22258
rect 46898 22206 46900 22258
rect 46844 22194 46900 22206
rect 46956 22482 47012 22494
rect 46956 22430 46958 22482
rect 47010 22430 47012 22482
rect 46620 21758 46622 21810
rect 46674 21758 46676 21810
rect 46620 21746 46676 21758
rect 46396 21634 46452 21644
rect 46956 21586 47012 22430
rect 47180 22372 47236 22382
rect 47180 22278 47236 22316
rect 47516 22370 47572 23212
rect 47628 23156 47684 25116
rect 47964 24724 48020 24734
rect 47852 24498 47908 24510
rect 47852 24446 47854 24498
rect 47906 24446 47908 24498
rect 47852 23268 47908 24446
rect 47964 24052 48020 24668
rect 48076 24052 48132 26236
rect 48188 26226 48244 26236
rect 48188 25844 48244 25854
rect 48188 25618 48244 25788
rect 48188 25566 48190 25618
rect 48242 25566 48244 25618
rect 48188 25554 48244 25566
rect 48412 24724 48468 36316
rect 48412 24658 48468 24668
rect 48188 24052 48244 24062
rect 48076 24050 48244 24052
rect 48076 23998 48190 24050
rect 48242 23998 48244 24050
rect 48076 23996 48244 23998
rect 47964 23986 48020 23996
rect 48188 23986 48244 23996
rect 47852 23202 47908 23212
rect 47964 23266 48020 23278
rect 47964 23214 47966 23266
rect 48018 23214 48020 23266
rect 47628 23154 47796 23156
rect 47628 23102 47630 23154
rect 47682 23102 47796 23154
rect 47628 23100 47796 23102
rect 47628 23090 47684 23100
rect 47516 22318 47518 22370
rect 47570 22318 47572 22370
rect 47516 22306 47572 22318
rect 47740 22370 47796 23100
rect 47740 22318 47742 22370
rect 47794 22318 47796 22370
rect 47740 22306 47796 22318
rect 47516 22146 47572 22158
rect 47516 22094 47518 22146
rect 47570 22094 47572 22146
rect 46956 21534 46958 21586
rect 47010 21534 47012 21586
rect 46172 21476 46228 21486
rect 45500 21474 46228 21476
rect 45500 21422 46174 21474
rect 46226 21422 46228 21474
rect 45500 21420 46228 21422
rect 46172 21410 46228 21420
rect 45388 20972 45668 21028
rect 45052 20862 45054 20914
rect 45106 20862 45108 20914
rect 45052 20244 45108 20862
rect 45052 20178 45108 20188
rect 45388 20802 45444 20814
rect 45388 20750 45390 20802
rect 45442 20750 45444 20802
rect 45052 20020 45108 20030
rect 45052 19926 45108 19964
rect 45276 20018 45332 20030
rect 45276 19966 45278 20018
rect 45330 19966 45332 20018
rect 44604 19908 44660 19918
rect 44604 19348 44660 19852
rect 45276 19908 45332 19966
rect 45276 19842 45332 19852
rect 45052 19796 45108 19806
rect 45052 19794 45220 19796
rect 45052 19742 45054 19794
rect 45106 19742 45220 19794
rect 45052 19740 45220 19742
rect 45052 19730 45108 19740
rect 44604 19282 44660 19292
rect 44268 19012 44324 19022
rect 44268 19010 44772 19012
rect 44268 18958 44270 19010
rect 44322 18958 44772 19010
rect 44268 18956 44772 18958
rect 44268 18946 44324 18956
rect 44492 18562 44548 18574
rect 44492 18510 44494 18562
rect 44546 18510 44548 18562
rect 43372 17838 43374 17890
rect 43426 17838 43428 17890
rect 43372 17826 43428 17838
rect 43932 17948 44100 18004
rect 44156 18228 44212 18238
rect 44492 18228 44548 18510
rect 44716 18564 44772 18956
rect 45052 19010 45108 19022
rect 45052 18958 45054 19010
rect 45106 18958 45108 19010
rect 45052 18900 45108 18958
rect 45164 18900 45220 19740
rect 45388 19234 45444 20750
rect 45388 19182 45390 19234
rect 45442 19182 45444 19234
rect 45164 18844 45332 18900
rect 45052 18834 45108 18844
rect 45164 18674 45220 18686
rect 45164 18622 45166 18674
rect 45218 18622 45220 18674
rect 45164 18564 45220 18622
rect 44716 18508 45220 18564
rect 44716 18450 44772 18508
rect 45276 18452 45332 18844
rect 44716 18398 44718 18450
rect 44770 18398 44772 18450
rect 44716 18386 44772 18398
rect 45164 18396 45332 18452
rect 44156 18226 44548 18228
rect 44156 18174 44158 18226
rect 44210 18174 44548 18226
rect 44156 18172 44548 18174
rect 43372 17666 43428 17678
rect 43596 17668 43652 17678
rect 43372 17614 43374 17666
rect 43426 17614 43428 17666
rect 43372 17556 43428 17614
rect 43372 17490 43428 17500
rect 43484 17612 43596 17668
rect 43484 16098 43540 17612
rect 43596 17602 43652 17612
rect 43820 16772 43876 16782
rect 43484 16046 43486 16098
rect 43538 16046 43540 16098
rect 43484 16034 43540 16046
rect 43708 16770 43876 16772
rect 43708 16718 43822 16770
rect 43874 16718 43876 16770
rect 43708 16716 43876 16718
rect 43708 16100 43764 16716
rect 43820 16706 43876 16716
rect 43932 16772 43988 17948
rect 44044 17780 44100 17790
rect 44044 17686 44100 17724
rect 44156 17108 44212 18172
rect 45164 17780 45220 18396
rect 45388 18340 45444 19182
rect 45500 18564 45556 18574
rect 45500 18470 45556 18508
rect 45052 17724 45220 17780
rect 45276 18284 45444 18340
rect 44716 17668 44772 17678
rect 44716 17574 44772 17612
rect 44940 17442 44996 17454
rect 44940 17390 44942 17442
rect 44994 17390 44996 17442
rect 44156 17052 44436 17108
rect 43932 16706 43988 16716
rect 44156 16884 44212 16894
rect 43708 15986 43764 16044
rect 43820 16100 43876 16110
rect 44044 16100 44100 16110
rect 43820 16098 44044 16100
rect 43820 16046 43822 16098
rect 43874 16046 44044 16098
rect 43820 16044 44044 16046
rect 43820 16034 43876 16044
rect 43708 15934 43710 15986
rect 43762 15934 43764 15986
rect 43708 15922 43764 15934
rect 43484 15540 43540 15550
rect 43484 15446 43540 15484
rect 43932 15540 43988 15550
rect 43932 15446 43988 15484
rect 43708 14532 43764 14542
rect 43484 14418 43540 14430
rect 43484 14366 43486 14418
rect 43538 14366 43540 14418
rect 43484 13972 43540 14366
rect 43596 13972 43652 13982
rect 43484 13970 43652 13972
rect 43484 13918 43598 13970
rect 43650 13918 43652 13970
rect 43484 13916 43652 13918
rect 43260 13906 43316 13916
rect 43596 13906 43652 13916
rect 43484 13746 43540 13758
rect 43484 13694 43486 13746
rect 43538 13694 43540 13746
rect 43148 13076 43204 13086
rect 43148 12982 43204 13020
rect 43036 12786 43092 12796
rect 42588 12402 42868 12404
rect 42588 12350 42814 12402
rect 42866 12350 42868 12402
rect 42588 12348 42868 12350
rect 41916 12292 41972 12302
rect 41804 12290 41972 12292
rect 41804 12238 41918 12290
rect 41970 12238 41972 12290
rect 41804 12236 41972 12238
rect 41916 12226 41972 12236
rect 42364 12068 42420 12078
rect 42364 11974 42420 12012
rect 41468 11414 41524 11452
rect 42364 11508 42420 11518
rect 40236 11396 40292 11406
rect 40236 11302 40292 11340
rect 41132 11396 41188 11406
rect 41132 11302 41188 11340
rect 42028 11396 42084 11406
rect 42028 11302 42084 11340
rect 42364 11394 42420 11452
rect 42364 11342 42366 11394
rect 42418 11342 42420 11394
rect 42364 11330 42420 11342
rect 41020 11284 41076 11294
rect 40012 10836 40068 10846
rect 40012 10834 40292 10836
rect 40012 10782 40014 10834
rect 40066 10782 40292 10834
rect 40012 10780 40292 10782
rect 40012 10770 40068 10780
rect 40012 10612 40068 10622
rect 40012 10518 40068 10556
rect 40124 9940 40180 9950
rect 40012 9828 40068 9838
rect 39788 9826 40068 9828
rect 39788 9774 40014 9826
rect 40066 9774 40068 9826
rect 39788 9772 40068 9774
rect 40012 9762 40068 9772
rect 39676 9550 39678 9602
rect 39730 9550 39732 9602
rect 38556 9102 38558 9154
rect 38610 9102 38612 9154
rect 38556 9090 38612 9102
rect 38780 9266 38836 9278
rect 38780 9214 38782 9266
rect 38834 9214 38836 9266
rect 38444 8306 38500 8316
rect 38780 8260 38836 9214
rect 38892 9154 38948 9324
rect 39340 9268 39396 9278
rect 38892 9102 38894 9154
rect 38946 9102 38948 9154
rect 38892 9090 38948 9102
rect 39116 9212 39340 9268
rect 39116 9154 39172 9212
rect 39340 9202 39396 9212
rect 39116 9102 39118 9154
rect 39170 9102 39172 9154
rect 39116 9090 39172 9102
rect 39676 9042 39732 9550
rect 39676 8990 39678 9042
rect 39730 8990 39732 9042
rect 39676 8978 39732 8990
rect 39900 9268 39956 9278
rect 38892 8260 38948 8270
rect 39564 8260 39620 8270
rect 38780 8258 39620 8260
rect 38780 8206 38894 8258
rect 38946 8206 39566 8258
rect 39618 8206 39620 8258
rect 38780 8204 39620 8206
rect 38892 8194 38948 8204
rect 39564 8194 39620 8204
rect 39788 8258 39844 8270
rect 39788 8206 39790 8258
rect 39842 8206 39844 8258
rect 38444 8034 38500 8046
rect 38444 7982 38446 8034
rect 38498 7982 38500 8034
rect 38444 7924 38500 7982
rect 38668 8036 38724 8046
rect 38668 7942 38724 7980
rect 38780 8036 38836 8046
rect 38780 8034 39060 8036
rect 38780 7982 38782 8034
rect 38834 7982 39060 8034
rect 38780 7980 39060 7982
rect 38780 7970 38836 7980
rect 38556 7924 38612 7934
rect 38444 7868 38556 7924
rect 38556 7858 38612 7868
rect 38220 7756 38500 7812
rect 38108 7382 38164 7420
rect 37884 7364 37940 7374
rect 37212 6850 37268 6860
rect 37324 7196 37604 7252
rect 37772 7252 37828 7262
rect 37100 6638 37102 6690
rect 37154 6638 37156 6690
rect 37100 6626 37156 6638
rect 35980 6578 36036 6590
rect 35980 6526 35982 6578
rect 36034 6526 36036 6578
rect 35980 6132 36036 6526
rect 35980 6066 36036 6076
rect 36092 6466 36148 6478
rect 36092 6414 36094 6466
rect 36146 6414 36148 6466
rect 35756 5906 35924 5908
rect 35756 5854 35758 5906
rect 35810 5854 35924 5906
rect 35756 5852 35924 5854
rect 35756 5842 35812 5852
rect 35308 5740 35700 5796
rect 34972 5684 35028 5694
rect 35028 5628 35140 5684
rect 34972 5618 35028 5628
rect 34636 5404 34916 5460
rect 34636 5236 34692 5246
rect 34636 5142 34692 5180
rect 34748 5124 34804 5134
rect 34748 5030 34804 5068
rect 34860 4452 34916 5404
rect 35084 5234 35140 5628
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35084 5182 35086 5234
rect 35138 5182 35140 5234
rect 35084 5170 35140 5182
rect 35644 5234 35700 5740
rect 35868 5684 35924 5694
rect 35868 5590 35924 5628
rect 35644 5182 35646 5234
rect 35698 5182 35700 5234
rect 35644 5170 35700 5182
rect 35980 5236 36036 5246
rect 36092 5236 36148 6414
rect 36204 6244 36260 6254
rect 36204 6130 36260 6188
rect 36204 6078 36206 6130
rect 36258 6078 36260 6130
rect 36204 6066 36260 6078
rect 36428 6132 36484 6142
rect 36428 6018 36484 6076
rect 36428 5966 36430 6018
rect 36482 5966 36484 6018
rect 36428 5954 36484 5966
rect 37212 6132 37268 6142
rect 36652 5906 36708 5918
rect 36652 5854 36654 5906
rect 36706 5854 36708 5906
rect 36652 5572 36708 5854
rect 36764 5796 36820 5806
rect 36764 5794 37156 5796
rect 36764 5742 36766 5794
rect 36818 5742 37156 5794
rect 36764 5740 37156 5742
rect 36764 5730 36820 5740
rect 36764 5572 36820 5582
rect 36652 5516 36764 5572
rect 36764 5506 36820 5516
rect 35980 5234 36148 5236
rect 35980 5182 35982 5234
rect 36034 5182 36148 5234
rect 35980 5180 36148 5182
rect 37100 5234 37156 5740
rect 37100 5182 37102 5234
rect 37154 5182 37156 5234
rect 35980 5170 36036 5180
rect 37100 5170 37156 5182
rect 36988 5124 37044 5134
rect 36764 5122 37044 5124
rect 36764 5070 36990 5122
rect 37042 5070 37044 5122
rect 36764 5068 37044 5070
rect 35980 5012 36036 5022
rect 34860 4386 34916 4396
rect 35196 4898 35252 4910
rect 35196 4846 35198 4898
rect 35250 4846 35252 4898
rect 35196 4450 35252 4846
rect 35196 4398 35198 4450
rect 35250 4398 35252 4450
rect 35196 4386 35252 4398
rect 35980 4338 36036 4956
rect 36092 4900 36148 4910
rect 36092 4806 36148 4844
rect 35980 4286 35982 4338
rect 36034 4286 36036 4338
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 35532 3668 35588 3678
rect 35980 3668 36036 4286
rect 36316 4228 36372 4238
rect 36316 4134 36372 4172
rect 35532 3666 36036 3668
rect 35532 3614 35534 3666
rect 35586 3614 36036 3666
rect 35532 3612 36036 3614
rect 35532 3602 35588 3612
rect 35980 3554 36036 3612
rect 36764 3666 36820 5068
rect 36988 5058 37044 5068
rect 37212 5012 37268 6076
rect 37324 5572 37380 7196
rect 37772 7158 37828 7196
rect 37772 6804 37828 6814
rect 37772 6578 37828 6748
rect 37772 6526 37774 6578
rect 37826 6526 37828 6578
rect 37772 6514 37828 6526
rect 37436 6468 37492 6478
rect 37492 6412 37716 6468
rect 37436 6374 37492 6412
rect 37660 6130 37716 6412
rect 37660 6078 37662 6130
rect 37714 6078 37716 6130
rect 37660 6066 37716 6078
rect 37324 5506 37380 5516
rect 37212 4946 37268 4956
rect 36764 3614 36766 3666
rect 36818 3614 36820 3666
rect 36764 3602 36820 3614
rect 35980 3502 35982 3554
rect 36034 3502 36036 3554
rect 35980 3490 36036 3502
rect 37884 3556 37940 7308
rect 38332 7364 38388 7374
rect 38332 7270 38388 7308
rect 38220 7252 38276 7262
rect 38108 6916 38164 6926
rect 38108 6822 38164 6860
rect 38220 6914 38276 7196
rect 38220 6862 38222 6914
rect 38274 6862 38276 6914
rect 38220 6850 38276 6862
rect 38444 6356 38500 7756
rect 38892 7700 38948 7710
rect 38668 7476 38724 7486
rect 38668 7382 38724 7420
rect 38780 7362 38836 7374
rect 38780 7310 38782 7362
rect 38834 7310 38836 7362
rect 38780 6916 38836 7310
rect 38892 7364 38948 7644
rect 39004 7364 39060 7980
rect 39228 8034 39284 8046
rect 39228 7982 39230 8034
rect 39282 7982 39284 8034
rect 39228 7700 39284 7982
rect 39788 8036 39844 8206
rect 39676 7924 39732 7934
rect 39284 7644 39620 7700
rect 39228 7634 39284 7644
rect 39116 7588 39172 7598
rect 39116 7494 39172 7532
rect 39004 7308 39508 7364
rect 38892 7298 38948 7308
rect 38780 6850 38836 6860
rect 39340 7028 39396 7038
rect 38892 6804 38948 6814
rect 38780 6692 38836 6702
rect 38892 6692 38948 6748
rect 39116 6804 39172 6814
rect 39116 6802 39284 6804
rect 39116 6750 39118 6802
rect 39170 6750 39284 6802
rect 39116 6748 39284 6750
rect 39116 6738 39172 6748
rect 38780 6690 38948 6692
rect 38780 6638 38782 6690
rect 38834 6638 38948 6690
rect 38780 6636 38948 6638
rect 38780 6626 38836 6636
rect 38556 6580 38612 6590
rect 38556 6486 38612 6524
rect 39004 6578 39060 6590
rect 39004 6526 39006 6578
rect 39058 6526 39060 6578
rect 39004 6356 39060 6526
rect 38444 6300 39060 6356
rect 38780 5572 38836 5582
rect 38444 4900 38500 4910
rect 38444 4450 38500 4844
rect 38444 4398 38446 4450
rect 38498 4398 38500 4450
rect 38444 4386 38500 4398
rect 38780 3668 38836 5516
rect 39004 5460 39060 6300
rect 39228 5460 39284 6748
rect 39340 6130 39396 6972
rect 39452 6914 39508 7308
rect 39452 6862 39454 6914
rect 39506 6862 39508 6914
rect 39452 6850 39508 6862
rect 39564 6914 39620 7644
rect 39564 6862 39566 6914
rect 39618 6862 39620 6914
rect 39564 6850 39620 6862
rect 39676 7474 39732 7868
rect 39676 7422 39678 7474
rect 39730 7422 39732 7474
rect 39340 6078 39342 6130
rect 39394 6078 39396 6130
rect 39340 6066 39396 6078
rect 39564 6468 39620 6478
rect 39564 6018 39620 6412
rect 39676 6244 39732 7422
rect 39788 7476 39844 7980
rect 39900 7700 39956 9212
rect 40012 9266 40068 9278
rect 40012 9214 40014 9266
rect 40066 9214 40068 9266
rect 40012 8148 40068 9214
rect 40124 9154 40180 9884
rect 40124 9102 40126 9154
rect 40178 9102 40180 9154
rect 40124 9090 40180 9102
rect 40012 8082 40068 8092
rect 40124 8372 40180 8382
rect 40236 8372 40292 10780
rect 41020 10722 41076 11228
rect 42476 11170 42532 11182
rect 42476 11118 42478 11170
rect 42530 11118 42532 11170
rect 42476 10836 42532 11118
rect 41020 10670 41022 10722
rect 41074 10670 41076 10722
rect 41020 10658 41076 10670
rect 42364 10780 42532 10836
rect 40348 10610 40404 10622
rect 40348 10558 40350 10610
rect 40402 10558 40404 10610
rect 40348 9828 40404 10558
rect 40908 10610 40964 10622
rect 41804 10612 41860 10622
rect 40908 10558 40910 10610
rect 40962 10558 40964 10610
rect 40908 10500 40964 10558
rect 41692 10610 41860 10612
rect 41692 10558 41806 10610
rect 41858 10558 41860 10610
rect 41692 10556 41860 10558
rect 40908 10434 40964 10444
rect 41020 10498 41076 10510
rect 41020 10446 41022 10498
rect 41074 10446 41076 10498
rect 41020 9940 41076 10446
rect 40348 9762 40404 9772
rect 40908 9884 41076 9940
rect 41692 10052 41748 10556
rect 41804 10546 41860 10556
rect 42364 10052 42420 10780
rect 42476 10612 42532 10622
rect 42588 10612 42644 12348
rect 42812 12338 42868 12348
rect 43484 11844 43540 13694
rect 43708 13746 43764 14476
rect 43932 14532 43988 14542
rect 43932 13748 43988 14476
rect 43708 13694 43710 13746
rect 43762 13694 43764 13746
rect 43708 13682 43764 13694
rect 43820 13746 43988 13748
rect 43820 13694 43934 13746
rect 43986 13694 43988 13746
rect 43820 13692 43988 13694
rect 43820 13188 43876 13692
rect 43932 13682 43988 13692
rect 43484 11778 43540 11788
rect 43708 13132 43876 13188
rect 43036 11508 43092 11518
rect 43036 11414 43092 11452
rect 43484 11508 43540 11518
rect 43484 11414 43540 11452
rect 42476 10610 42644 10612
rect 42476 10558 42478 10610
rect 42530 10558 42644 10610
rect 42476 10556 42644 10558
rect 42700 11170 42756 11182
rect 42700 11118 42702 11170
rect 42754 11118 42756 11170
rect 42476 10546 42532 10556
rect 42476 10052 42532 10062
rect 42364 9996 42476 10052
rect 40460 9156 40516 9166
rect 40908 9156 40964 9884
rect 41020 9716 41076 9726
rect 41020 9622 41076 9660
rect 40348 9044 40404 9054
rect 40460 9044 40516 9100
rect 40348 9042 40516 9044
rect 40348 8990 40350 9042
rect 40402 8990 40516 9042
rect 40348 8988 40516 8990
rect 40348 8978 40404 8988
rect 40236 8316 40404 8372
rect 39900 7644 40068 7700
rect 40012 7476 40068 7644
rect 40124 7698 40180 8316
rect 40236 8036 40292 8046
rect 40236 7942 40292 7980
rect 40124 7646 40126 7698
rect 40178 7646 40180 7698
rect 40124 7634 40180 7646
rect 40236 7700 40292 7710
rect 40236 7606 40292 7644
rect 40348 7698 40404 8316
rect 40348 7646 40350 7698
rect 40402 7646 40404 7698
rect 40348 7588 40404 7646
rect 40348 7522 40404 7532
rect 40460 7476 40516 8988
rect 40796 9154 40964 9156
rect 40796 9102 40910 9154
rect 40962 9102 40964 9154
rect 40796 9100 40964 9102
rect 40796 8372 40852 9100
rect 40908 9090 40964 9100
rect 41020 9156 41076 9166
rect 41020 9154 41188 9156
rect 41020 9102 41022 9154
rect 41074 9102 41188 9154
rect 41020 9100 41188 9102
rect 41020 9090 41076 9100
rect 40796 8306 40852 8316
rect 40908 8258 40964 8270
rect 40908 8206 40910 8258
rect 40962 8206 40964 8258
rect 40908 7700 40964 8206
rect 41020 8260 41076 8270
rect 41020 7924 41076 8204
rect 41020 7858 41076 7868
rect 41132 7700 41188 9100
rect 41244 9042 41300 9054
rect 41244 8990 41246 9042
rect 41298 8990 41300 9042
rect 41244 8260 41300 8990
rect 41692 8930 41748 9996
rect 42476 9986 42532 9996
rect 41692 8878 41694 8930
rect 41746 8878 41748 8930
rect 41692 8866 41748 8878
rect 41916 9828 41972 9838
rect 41244 8194 41300 8204
rect 41356 8484 41412 8494
rect 41356 8148 41412 8428
rect 41916 8260 41972 9772
rect 42140 9828 42196 9838
rect 42364 9828 42420 9838
rect 42140 9826 42420 9828
rect 42140 9774 42142 9826
rect 42194 9774 42366 9826
rect 42418 9774 42420 9826
rect 42140 9772 42420 9774
rect 42140 9762 42196 9772
rect 42364 9762 42420 9772
rect 42476 8932 42532 8942
rect 42252 8372 42308 8382
rect 42140 8260 42196 8270
rect 41916 8258 42084 8260
rect 41916 8206 41918 8258
rect 41970 8206 42084 8258
rect 41916 8204 42084 8206
rect 41916 8194 41972 8204
rect 41356 8146 41524 8148
rect 41356 8094 41358 8146
rect 41410 8094 41524 8146
rect 41356 8092 41524 8094
rect 41356 8082 41412 8092
rect 40908 7634 40964 7644
rect 41020 7644 41188 7700
rect 41244 7700 41300 7710
rect 40908 7476 40964 7486
rect 40012 7420 40292 7476
rect 40460 7474 40964 7476
rect 40460 7422 40910 7474
rect 40962 7422 40964 7474
rect 40460 7420 40964 7422
rect 39788 7410 39844 7420
rect 40124 7140 40180 7150
rect 40124 6804 40180 7084
rect 40124 6690 40180 6748
rect 40124 6638 40126 6690
rect 40178 6638 40180 6690
rect 40124 6626 40180 6638
rect 40236 6692 40292 7420
rect 40348 6692 40404 6702
rect 40236 6690 40404 6692
rect 40236 6638 40350 6690
rect 40402 6638 40404 6690
rect 40236 6636 40404 6638
rect 39788 6580 39844 6590
rect 39788 6486 39844 6524
rect 40236 6468 40292 6478
rect 40236 6374 40292 6412
rect 40348 6244 40404 6636
rect 39676 6188 40292 6244
rect 40236 6130 40292 6188
rect 40348 6178 40404 6188
rect 40236 6078 40238 6130
rect 40290 6078 40292 6130
rect 40236 6066 40292 6078
rect 39564 5966 39566 6018
rect 39618 5966 39620 6018
rect 39564 5954 39620 5966
rect 40796 5796 40852 7420
rect 40908 7410 40964 7420
rect 41020 7252 41076 7644
rect 41244 7586 41300 7644
rect 41244 7534 41246 7586
rect 41298 7534 41300 7586
rect 40908 7196 41076 7252
rect 41132 7474 41188 7486
rect 41132 7422 41134 7474
rect 41186 7422 41188 7474
rect 40908 6466 40964 7196
rect 40908 6414 40910 6466
rect 40962 6414 40964 6466
rect 40908 6356 40964 6414
rect 40908 6290 40964 6300
rect 41020 6020 41076 6030
rect 41020 5906 41076 5964
rect 41020 5854 41022 5906
rect 41074 5854 41076 5906
rect 40908 5796 40964 5806
rect 40796 5740 40908 5796
rect 40908 5730 40964 5740
rect 39676 5684 39732 5694
rect 39676 5682 40068 5684
rect 39676 5630 39678 5682
rect 39730 5630 40068 5682
rect 39676 5628 40068 5630
rect 39676 5618 39732 5628
rect 39788 5460 39844 5470
rect 39228 5404 39620 5460
rect 39004 5394 39060 5404
rect 39228 5124 39284 5134
rect 39116 5122 39284 5124
rect 39116 5070 39230 5122
rect 39282 5070 39284 5122
rect 39116 5068 39284 5070
rect 38892 5012 38948 5022
rect 39116 5012 39172 5068
rect 39228 5058 39284 5068
rect 38948 4956 39172 5012
rect 38892 4918 38948 4956
rect 39116 4564 39172 4956
rect 39116 4338 39172 4508
rect 39564 4450 39620 5404
rect 39564 4398 39566 4450
rect 39618 4398 39620 4450
rect 39564 4386 39620 4398
rect 39116 4286 39118 4338
rect 39170 4286 39172 4338
rect 39116 4274 39172 4286
rect 39676 4116 39732 4126
rect 39676 4022 39732 4060
rect 38892 3668 38948 3678
rect 38780 3666 38948 3668
rect 38780 3614 38894 3666
rect 38946 3614 38948 3666
rect 38780 3612 38948 3614
rect 38892 3602 38948 3612
rect 39788 3666 39844 5404
rect 40012 5234 40068 5628
rect 40012 5182 40014 5234
rect 40066 5182 40068 5234
rect 40012 5170 40068 5182
rect 40124 4564 40180 4574
rect 40124 4470 40180 4508
rect 41020 4564 41076 5854
rect 41020 4498 41076 4508
rect 41132 4450 41188 7422
rect 41244 7140 41300 7534
rect 41244 7074 41300 7084
rect 41468 7698 41524 8092
rect 41468 7646 41470 7698
rect 41522 7646 41524 7698
rect 41468 7028 41524 7646
rect 41580 8146 41636 8158
rect 41580 8094 41582 8146
rect 41634 8094 41636 8146
rect 41580 7700 41636 8094
rect 41580 7634 41636 7644
rect 41692 8034 41748 8046
rect 41692 7982 41694 8034
rect 41746 7982 41748 8034
rect 41468 6962 41524 6972
rect 41356 6690 41412 6702
rect 41356 6638 41358 6690
rect 41410 6638 41412 6690
rect 41356 6020 41412 6638
rect 41692 6468 41748 7982
rect 41916 8036 41972 8046
rect 41804 7476 41860 7486
rect 41804 7382 41860 7420
rect 41916 7474 41972 7980
rect 41916 7422 41918 7474
rect 41970 7422 41972 7474
rect 41916 7410 41972 7422
rect 42028 7252 42084 8204
rect 42140 8166 42196 8204
rect 42252 7474 42308 8316
rect 42476 8034 42532 8876
rect 42588 8260 42644 8270
rect 42700 8260 42756 11118
rect 43148 10724 43204 10734
rect 43148 10630 43204 10668
rect 42812 10052 42868 10062
rect 42812 9958 42868 9996
rect 43036 9828 43092 9838
rect 43036 9734 43092 9772
rect 43260 9826 43316 9838
rect 43260 9774 43262 9826
rect 43314 9774 43316 9826
rect 43260 9156 43316 9774
rect 43484 9714 43540 9726
rect 43484 9662 43486 9714
rect 43538 9662 43540 9714
rect 43484 9268 43540 9662
rect 43484 9202 43540 9212
rect 43260 9090 43316 9100
rect 42588 8258 42756 8260
rect 42588 8206 42590 8258
rect 42642 8206 42756 8258
rect 42588 8204 42756 8206
rect 42812 8596 42868 8606
rect 42812 8260 42868 8540
rect 42588 8194 42644 8204
rect 42812 8166 42868 8204
rect 43148 8148 43204 8158
rect 43148 8054 43204 8092
rect 42476 7982 42478 8034
rect 42530 7982 42532 8034
rect 42476 7970 42532 7982
rect 43260 8036 43316 8046
rect 43260 7942 43316 7980
rect 43372 8034 43428 8046
rect 43372 7982 43374 8034
rect 43426 7982 43428 8034
rect 42812 7924 42868 7934
rect 42812 7698 42868 7868
rect 43372 7924 43428 7982
rect 43372 7858 43428 7868
rect 43708 7700 43764 13132
rect 44044 13076 44100 16044
rect 44156 14530 44212 16828
rect 44156 14478 44158 14530
rect 44210 14478 44212 14530
rect 44156 14466 44212 14478
rect 44268 15426 44324 15438
rect 44268 15374 44270 15426
rect 44322 15374 44324 15426
rect 44268 14532 44324 15374
rect 44380 15316 44436 17052
rect 44940 16994 44996 17390
rect 44940 16942 44942 16994
rect 44994 16942 44996 16994
rect 44940 16930 44996 16942
rect 45052 16100 45108 17724
rect 45164 17556 45220 17566
rect 45164 17462 45220 17500
rect 45276 16884 45332 18284
rect 45612 17780 45668 20972
rect 46060 20692 46116 20702
rect 46060 20690 46676 20692
rect 46060 20638 46062 20690
rect 46114 20638 46676 20690
rect 46060 20636 46676 20638
rect 46060 20626 46116 20636
rect 46396 20244 46452 20254
rect 46396 20150 46452 20188
rect 45836 20020 45892 20030
rect 45836 18564 45892 19964
rect 46508 20018 46564 20030
rect 46508 19966 46510 20018
rect 46562 19966 46564 20018
rect 46060 19122 46116 19134
rect 46508 19124 46564 19966
rect 46620 19460 46676 20636
rect 46732 20130 46788 20142
rect 46732 20078 46734 20130
rect 46786 20078 46788 20130
rect 46732 19572 46788 20078
rect 46956 20132 47012 21534
rect 47180 21700 47236 21710
rect 47180 21588 47236 21644
rect 47516 21698 47572 22094
rect 47516 21646 47518 21698
rect 47570 21646 47572 21698
rect 47516 21634 47572 21646
rect 47852 21700 47908 21710
rect 47852 21606 47908 21644
rect 47180 21586 47348 21588
rect 47180 21534 47182 21586
rect 47234 21534 47348 21586
rect 47180 21532 47348 21534
rect 47180 21522 47236 21532
rect 47068 21476 47124 21486
rect 47068 21382 47124 21420
rect 47292 20242 47348 21532
rect 47964 21476 48020 23214
rect 48076 23044 48132 23054
rect 48132 22988 48356 23044
rect 48076 22978 48132 22988
rect 47292 20190 47294 20242
rect 47346 20190 47348 20242
rect 47292 20178 47348 20190
rect 47516 21420 48020 21476
rect 48076 22260 48132 22270
rect 48076 21586 48132 22204
rect 48076 21534 48078 21586
rect 48130 21534 48132 21586
rect 47180 20132 47236 20142
rect 46956 20130 47236 20132
rect 46956 20078 47182 20130
rect 47234 20078 47236 20130
rect 46956 20076 47236 20078
rect 47180 20066 47236 20076
rect 47516 20130 47572 21420
rect 48076 20916 48132 21534
rect 48076 20850 48132 20860
rect 48188 20914 48244 20926
rect 48188 20862 48190 20914
rect 48242 20862 48244 20914
rect 48188 20188 48244 20862
rect 47516 20078 47518 20130
rect 47570 20078 47572 20130
rect 47516 20066 47572 20078
rect 47628 20132 48244 20188
rect 46844 20020 46900 20030
rect 46844 19926 46900 19964
rect 47068 19796 47124 19806
rect 46732 19516 47012 19572
rect 46620 19404 46900 19460
rect 46060 19070 46062 19122
rect 46114 19070 46116 19122
rect 46060 18676 46116 19070
rect 46284 19068 46564 19124
rect 46172 18676 46228 18686
rect 46060 18674 46228 18676
rect 46060 18622 46174 18674
rect 46226 18622 46228 18674
rect 46060 18620 46228 18622
rect 46172 18610 46228 18620
rect 45836 18116 45892 18508
rect 45948 18450 46004 18462
rect 45948 18398 45950 18450
rect 46002 18398 46004 18450
rect 45948 18340 46004 18398
rect 46172 18452 46228 18462
rect 46284 18452 46340 19068
rect 46172 18450 46340 18452
rect 46172 18398 46174 18450
rect 46226 18398 46340 18450
rect 46172 18396 46340 18398
rect 46396 18450 46452 18462
rect 46396 18398 46398 18450
rect 46450 18398 46452 18450
rect 46172 18386 46228 18396
rect 46004 18284 46116 18340
rect 45948 18274 46004 18284
rect 45836 18060 46004 18116
rect 45500 17724 45668 17780
rect 45388 17668 45444 17678
rect 45388 17574 45444 17612
rect 45500 17332 45556 17724
rect 45612 17556 45668 17566
rect 45612 17462 45668 17500
rect 45948 17554 46004 18060
rect 45948 17502 45950 17554
rect 46002 17502 46004 17554
rect 45836 17442 45892 17454
rect 45836 17390 45838 17442
rect 45890 17390 45892 17442
rect 45500 17276 45668 17332
rect 45332 16828 45444 16884
rect 45276 16818 45332 16828
rect 45052 15538 45108 16044
rect 45388 16098 45444 16828
rect 45388 16046 45390 16098
rect 45442 16046 45444 16098
rect 45388 16034 45444 16046
rect 45052 15486 45054 15538
rect 45106 15486 45108 15538
rect 45052 15474 45108 15486
rect 45388 15426 45444 15438
rect 45388 15374 45390 15426
rect 45442 15374 45444 15426
rect 44380 15250 44436 15260
rect 44716 15316 44772 15326
rect 44268 14466 44324 14476
rect 44044 13020 44324 13076
rect 43820 12964 43876 12974
rect 43876 12908 44212 12964
rect 43820 12870 43876 12908
rect 44156 12404 44212 12908
rect 44156 12310 44212 12348
rect 44268 11284 44324 13020
rect 44716 12740 44772 15260
rect 45388 15316 45444 15374
rect 45388 15250 45444 15260
rect 45500 15204 45556 15214
rect 45276 14530 45332 14542
rect 45276 14478 45278 14530
rect 45330 14478 45332 14530
rect 44940 14308 44996 14318
rect 45276 14308 45332 14478
rect 44940 14306 45332 14308
rect 44940 14254 44942 14306
rect 44994 14254 45332 14306
rect 44940 14252 45332 14254
rect 44828 12740 44884 12750
rect 44716 12738 44884 12740
rect 44716 12686 44830 12738
rect 44882 12686 44884 12738
rect 44716 12684 44884 12686
rect 44044 11228 44324 11284
rect 44380 11844 44436 11854
rect 44044 9826 44100 11228
rect 44044 9774 44046 9826
rect 44098 9774 44100 9826
rect 43820 8932 43876 8942
rect 43820 8838 43876 8876
rect 43820 8258 43876 8270
rect 43820 8206 43822 8258
rect 43874 8206 43876 8258
rect 43820 8036 43876 8206
rect 44044 8036 44100 9774
rect 44268 11060 44324 11070
rect 44268 9714 44324 11004
rect 44268 9662 44270 9714
rect 44322 9662 44324 9714
rect 44268 9650 44324 9662
rect 44156 8260 44212 8270
rect 44156 8166 44212 8204
rect 44044 7980 44324 8036
rect 43820 7970 43876 7980
rect 42812 7646 42814 7698
rect 42866 7646 42868 7698
rect 42812 7634 42868 7646
rect 43596 7644 43764 7700
rect 43820 7700 43876 7710
rect 44156 7700 44212 7710
rect 43820 7698 44156 7700
rect 43820 7646 43822 7698
rect 43874 7646 44156 7698
rect 43820 7644 44156 7646
rect 42252 7422 42254 7474
rect 42306 7422 42308 7474
rect 42252 7410 42308 7422
rect 42476 7588 42532 7598
rect 42476 7474 42532 7532
rect 42476 7422 42478 7474
rect 42530 7422 42532 7474
rect 42476 7410 42532 7422
rect 41692 6402 41748 6412
rect 41916 7196 42084 7252
rect 43260 7362 43316 7374
rect 43260 7310 43262 7362
rect 43314 7310 43316 7362
rect 41356 5954 41412 5964
rect 41804 5796 41860 5806
rect 41244 5794 41860 5796
rect 41244 5742 41806 5794
rect 41858 5742 41860 5794
rect 41244 5740 41860 5742
rect 41244 4562 41300 5740
rect 41804 5730 41860 5740
rect 41916 5572 41972 7196
rect 43260 7028 43316 7310
rect 43596 7252 43652 7644
rect 43820 7634 43876 7644
rect 43708 7476 43764 7486
rect 43708 7382 43764 7420
rect 43596 7196 43764 7252
rect 43260 6962 43316 6972
rect 42140 6580 42196 6590
rect 42140 6486 42196 6524
rect 42476 6468 42532 6478
rect 41244 4510 41246 4562
rect 41298 4510 41300 4562
rect 41244 4498 41300 4510
rect 41804 5516 41972 5572
rect 42140 6244 42196 6254
rect 41132 4398 41134 4450
rect 41186 4398 41188 4450
rect 41132 4386 41188 4398
rect 41580 4228 41636 4238
rect 41804 4228 41860 5516
rect 42140 5234 42196 6188
rect 42140 5182 42142 5234
rect 42194 5182 42196 5234
rect 42140 5170 42196 5182
rect 42476 5234 42532 6412
rect 43708 6356 43764 7196
rect 43932 6916 43988 7644
rect 44156 7634 44212 7644
rect 44268 7698 44324 7980
rect 44268 7646 44270 7698
rect 44322 7646 44324 7698
rect 44268 7634 44324 7646
rect 44044 7476 44100 7486
rect 44044 7474 44212 7476
rect 44044 7422 44046 7474
rect 44098 7422 44212 7474
rect 44044 7420 44212 7422
rect 44044 7410 44100 7420
rect 44156 7028 44212 7420
rect 44380 7252 44436 11788
rect 44492 9604 44548 9614
rect 44492 9042 44548 9548
rect 44716 9268 44772 12684
rect 44828 12674 44884 12684
rect 44940 12404 44996 14252
rect 45500 13858 45556 15148
rect 45612 14756 45668 17276
rect 45836 16772 45892 17390
rect 45836 16706 45892 16716
rect 45948 15428 46004 17502
rect 46060 17108 46116 18284
rect 46396 17890 46452 18398
rect 46396 17838 46398 17890
rect 46450 17838 46452 17890
rect 46396 17826 46452 17838
rect 46732 18450 46788 18462
rect 46732 18398 46734 18450
rect 46786 18398 46788 18450
rect 46732 17666 46788 18398
rect 46844 18450 46900 19404
rect 46844 18398 46846 18450
rect 46898 18398 46900 18450
rect 46844 18386 46900 18398
rect 46956 19348 47012 19516
rect 46732 17614 46734 17666
rect 46786 17614 46788 17666
rect 46732 17602 46788 17614
rect 46284 17556 46340 17566
rect 46060 17052 46228 17108
rect 46060 16884 46116 16894
rect 46060 16210 46116 16828
rect 46060 16158 46062 16210
rect 46114 16158 46116 16210
rect 46060 16146 46116 16158
rect 45948 15362 46004 15372
rect 46172 15538 46228 17052
rect 46172 15486 46174 15538
rect 46226 15486 46228 15538
rect 45836 15314 45892 15326
rect 45836 15262 45838 15314
rect 45890 15262 45892 15314
rect 45836 15204 45892 15262
rect 45836 15138 45892 15148
rect 46172 15148 46228 15486
rect 46284 15316 46340 17500
rect 46956 17554 47012 19292
rect 47068 18562 47124 19740
rect 47068 18510 47070 18562
rect 47122 18510 47124 18562
rect 47068 18498 47124 18510
rect 47180 18450 47236 18462
rect 47180 18398 47182 18450
rect 47234 18398 47236 18450
rect 47180 18340 47236 18398
rect 47180 18274 47236 18284
rect 46956 17502 46958 17554
rect 47010 17502 47012 17554
rect 46956 17490 47012 17502
rect 47068 17556 47124 17566
rect 47068 17462 47124 17500
rect 47516 17556 47572 17566
rect 47516 17462 47572 17500
rect 46396 17442 46452 17454
rect 46396 17390 46398 17442
rect 46450 17390 46452 17442
rect 46396 16772 46452 17390
rect 47292 16884 47348 16894
rect 47180 16882 47348 16884
rect 47180 16830 47294 16882
rect 47346 16830 47348 16882
rect 47180 16828 47348 16830
rect 47068 16772 47124 16782
rect 46452 16770 47124 16772
rect 46452 16718 47070 16770
rect 47122 16718 47124 16770
rect 46452 16716 47124 16718
rect 46396 16678 46452 16716
rect 47068 16706 47124 16716
rect 46956 16548 47012 16558
rect 46956 15538 47012 16492
rect 46956 15486 46958 15538
rect 47010 15486 47012 15538
rect 46956 15474 47012 15486
rect 47180 15538 47236 16828
rect 47292 16818 47348 16828
rect 47516 16884 47572 16894
rect 47516 16790 47572 16828
rect 47628 16548 47684 20132
rect 47852 20130 47908 20132
rect 47852 20078 47854 20130
rect 47906 20078 47908 20130
rect 47852 20066 47908 20078
rect 47740 20020 47796 20030
rect 47740 19926 47796 19964
rect 47852 19796 47908 19806
rect 47852 19702 47908 19740
rect 48188 19348 48244 19358
rect 48188 19254 48244 19292
rect 47852 18562 47908 18574
rect 47852 18510 47854 18562
rect 47906 18510 47908 18562
rect 47852 17778 47908 18510
rect 48076 18452 48132 18462
rect 47852 17726 47854 17778
rect 47906 17726 47908 17778
rect 47852 17714 47908 17726
rect 47964 18340 48020 18350
rect 47964 16994 48020 18284
rect 48076 17556 48132 18396
rect 48076 17490 48132 17500
rect 47964 16942 47966 16994
rect 48018 16942 48020 16994
rect 47964 16930 48020 16942
rect 47628 16482 47684 16492
rect 47740 16882 47796 16894
rect 47740 16830 47742 16882
rect 47794 16830 47796 16882
rect 47180 15486 47182 15538
rect 47234 15486 47236 15538
rect 47180 15474 47236 15486
rect 47740 15538 47796 16830
rect 48188 16210 48244 16222
rect 48188 16158 48190 16210
rect 48242 16158 48244 16210
rect 48076 15540 48132 15550
rect 48188 15540 48244 16158
rect 47740 15486 47742 15538
rect 47794 15486 47796 15538
rect 47740 15474 47796 15486
rect 47852 15538 48244 15540
rect 47852 15486 48078 15538
rect 48130 15486 48244 15538
rect 47852 15484 48244 15486
rect 47404 15428 47460 15438
rect 47404 15334 47460 15372
rect 47516 15426 47572 15438
rect 47516 15374 47518 15426
rect 47570 15374 47572 15426
rect 46284 15250 46340 15260
rect 46844 15316 46900 15326
rect 47516 15316 47572 15374
rect 47852 15316 47908 15484
rect 48076 15474 48132 15484
rect 47516 15260 47908 15316
rect 47964 15316 48020 15326
rect 46844 15222 46900 15260
rect 47964 15222 48020 15260
rect 46172 15092 46676 15148
rect 48076 15092 48132 15102
rect 45612 14690 45668 14700
rect 46060 14420 46116 14430
rect 46060 14326 46116 14364
rect 45500 13806 45502 13858
rect 45554 13806 45556 13858
rect 45500 13794 45556 13806
rect 45836 13860 45892 13870
rect 45836 13858 46564 13860
rect 45836 13806 45838 13858
rect 45890 13806 46564 13858
rect 45836 13804 46564 13806
rect 45164 12738 45220 12750
rect 45724 12740 45780 12750
rect 45164 12686 45166 12738
rect 45218 12686 45220 12738
rect 44996 12348 45108 12404
rect 44940 12310 44996 12348
rect 44828 11282 44884 11294
rect 44828 11230 44830 11282
rect 44882 11230 44884 11282
rect 44828 11060 44884 11230
rect 44940 11284 44996 11294
rect 44940 11190 44996 11228
rect 44828 10994 44884 11004
rect 44940 9604 44996 9614
rect 45052 9604 45108 12348
rect 45164 11396 45220 12686
rect 45388 12738 45780 12740
rect 45388 12686 45726 12738
rect 45778 12686 45780 12738
rect 45388 12684 45780 12686
rect 45276 12404 45332 12414
rect 45276 12178 45332 12348
rect 45276 12126 45278 12178
rect 45330 12126 45332 12178
rect 45276 12114 45332 12126
rect 45164 11330 45220 11340
rect 45388 11394 45444 12684
rect 45724 12674 45780 12684
rect 45388 11342 45390 11394
rect 45442 11342 45444 11394
rect 45388 11330 45444 11342
rect 45724 11620 45780 11630
rect 45724 11394 45780 11564
rect 45724 11342 45726 11394
rect 45778 11342 45780 11394
rect 45724 11330 45780 11342
rect 45836 11620 45892 13804
rect 46508 12962 46564 13804
rect 46620 13858 46676 15092
rect 47404 15090 48132 15092
rect 47404 15038 48078 15090
rect 48130 15038 48132 15090
rect 47404 15036 48132 15038
rect 46956 14420 47012 14430
rect 46956 13970 47012 14364
rect 46956 13918 46958 13970
rect 47010 13918 47012 13970
rect 46956 13906 47012 13918
rect 46620 13806 46622 13858
rect 46674 13806 46676 13858
rect 46620 13794 46676 13806
rect 46956 13748 47012 13758
rect 46956 13654 47012 13692
rect 47292 13748 47348 13758
rect 47404 13748 47460 15036
rect 48076 15026 48132 15036
rect 48188 14642 48244 14654
rect 48188 14590 48190 14642
rect 48242 14590 48244 14642
rect 47628 13972 47684 13982
rect 48188 13972 48244 14590
rect 47628 13970 48244 13972
rect 47628 13918 47630 13970
rect 47682 13918 48244 13970
rect 47628 13916 48244 13918
rect 47628 13906 47684 13916
rect 47292 13746 47460 13748
rect 47292 13694 47294 13746
rect 47346 13694 47460 13746
rect 47292 13692 47460 13694
rect 47516 13748 47572 13758
rect 47852 13748 47908 13758
rect 47516 13746 47796 13748
rect 47516 13694 47518 13746
rect 47570 13694 47796 13746
rect 47516 13692 47796 13694
rect 47292 13682 47348 13692
rect 47516 13682 47572 13692
rect 46508 12910 46510 12962
rect 46562 12910 46564 12962
rect 46508 12898 46564 12910
rect 46844 12964 46900 12974
rect 46844 12962 47012 12964
rect 46844 12910 46846 12962
rect 46898 12910 47012 12962
rect 46844 12908 47012 12910
rect 46844 12898 46900 12908
rect 46060 12852 46116 12862
rect 46060 12850 46340 12852
rect 46060 12798 46062 12850
rect 46114 12798 46340 12850
rect 46060 12796 46340 12798
rect 46060 12786 46116 12796
rect 45948 12738 46004 12750
rect 45948 12686 45950 12738
rect 46002 12686 46004 12738
rect 45948 12068 46004 12686
rect 46284 12628 46340 12796
rect 46844 12740 46900 12750
rect 46284 12562 46340 12572
rect 46396 12738 46900 12740
rect 46396 12686 46846 12738
rect 46898 12686 46900 12738
rect 46396 12684 46900 12686
rect 46396 12404 46452 12684
rect 46844 12674 46900 12684
rect 46060 12348 46452 12404
rect 46844 12516 46900 12526
rect 46060 12290 46116 12348
rect 46060 12238 46062 12290
rect 46114 12238 46116 12290
rect 46060 12226 46116 12238
rect 45948 12002 46004 12012
rect 46732 12180 46788 12190
rect 46396 11620 46452 11630
rect 45836 11564 46340 11620
rect 45836 11394 45892 11564
rect 45836 11342 45838 11394
rect 45890 11342 45892 11394
rect 45836 11330 45892 11342
rect 45276 11284 45332 11294
rect 45164 11172 45220 11182
rect 45164 11078 45220 11116
rect 45276 10498 45332 11228
rect 45500 11170 45556 11182
rect 45500 11118 45502 11170
rect 45554 11118 45556 11170
rect 45500 10724 45556 11118
rect 45500 10658 45556 10668
rect 46060 11172 46116 11182
rect 46060 10610 46116 11116
rect 46284 11060 46340 11564
rect 46396 11526 46452 11564
rect 46508 11396 46564 11406
rect 46508 11302 46564 11340
rect 46396 11284 46452 11294
rect 46396 11190 46452 11228
rect 46732 11060 46788 12124
rect 46844 11284 46900 12460
rect 46956 11396 47012 12908
rect 47180 12962 47236 12974
rect 47180 12910 47182 12962
rect 47234 12910 47236 12962
rect 46956 11340 47124 11396
rect 46844 11190 46900 11228
rect 46956 11170 47012 11182
rect 46956 11118 46958 11170
rect 47010 11118 47012 11170
rect 46956 11060 47012 11118
rect 47068 11172 47124 11340
rect 47180 11394 47236 12910
rect 47628 12738 47684 12750
rect 47628 12686 47630 12738
rect 47682 12686 47684 12738
rect 47628 12628 47684 12686
rect 47628 12562 47684 12572
rect 47180 11342 47182 11394
rect 47234 11342 47236 11394
rect 47180 11330 47236 11342
rect 47516 12068 47572 12078
rect 47516 11282 47572 12012
rect 47516 11230 47518 11282
rect 47570 11230 47572 11282
rect 47516 11218 47572 11230
rect 47628 11396 47684 11406
rect 47740 11396 47796 13692
rect 47852 13654 47908 13692
rect 47852 12852 47908 12862
rect 47852 12758 47908 12796
rect 47852 12180 47908 12190
rect 47964 12180 48020 13916
rect 48188 12738 48244 12750
rect 48188 12686 48190 12738
rect 48242 12686 48244 12738
rect 48188 12628 48244 12686
rect 48188 12562 48244 12572
rect 47908 12124 48020 12180
rect 47852 12114 47908 12124
rect 48188 12068 48244 12078
rect 48188 11974 48244 12012
rect 48300 11508 48356 22988
rect 48300 11442 48356 11452
rect 47684 11340 47796 11396
rect 47292 11172 47348 11182
rect 47068 11170 47348 11172
rect 47068 11118 47294 11170
rect 47346 11118 47348 11170
rect 47068 11116 47348 11118
rect 47292 11106 47348 11116
rect 46284 11004 46452 11060
rect 46732 11004 47012 11060
rect 46060 10558 46062 10610
rect 46114 10558 46116 10610
rect 46060 10546 46116 10558
rect 45276 10446 45278 10498
rect 45330 10446 45332 10498
rect 45276 10434 45332 10446
rect 46284 10498 46340 10510
rect 46284 10446 46286 10498
rect 46338 10446 46340 10498
rect 46284 10052 46340 10446
rect 46060 9996 46340 10052
rect 46396 10500 46452 11004
rect 46956 10836 47012 10846
rect 47628 10836 47684 11340
rect 46620 10834 47012 10836
rect 46620 10782 46958 10834
rect 47010 10782 47012 10834
rect 46620 10780 47012 10782
rect 46508 10724 46564 10734
rect 46620 10724 46676 10780
rect 46956 10770 47012 10780
rect 47292 10780 47684 10836
rect 46508 10722 46676 10724
rect 46508 10670 46510 10722
rect 46562 10670 46676 10722
rect 46508 10668 46676 10670
rect 47180 10722 47236 10734
rect 47180 10670 47182 10722
rect 47234 10670 47236 10722
rect 46508 10658 46564 10668
rect 46732 10610 46788 10622
rect 46732 10558 46734 10610
rect 46786 10558 46788 10610
rect 46732 10500 46788 10558
rect 46396 10444 46788 10500
rect 46956 10612 47012 10622
rect 46060 9938 46116 9996
rect 46060 9886 46062 9938
rect 46114 9886 46116 9938
rect 46060 9874 46116 9886
rect 45276 9826 45332 9838
rect 45276 9774 45278 9826
rect 45330 9774 45332 9826
rect 45276 9604 45332 9774
rect 44996 9548 45332 9604
rect 44940 9510 44996 9548
rect 44940 9268 44996 9278
rect 44716 9266 44996 9268
rect 44716 9214 44942 9266
rect 44994 9214 44996 9266
rect 44716 9212 44996 9214
rect 44940 9202 44996 9212
rect 44492 8990 44494 9042
rect 44546 8990 44548 9042
rect 44492 8260 44548 8990
rect 44492 7588 44548 8204
rect 45276 9154 45332 9166
rect 45276 9102 45278 9154
rect 45330 9102 45332 9154
rect 44940 8036 44996 8046
rect 44940 7942 44996 7980
rect 45052 7700 45108 7710
rect 45052 7606 45108 7644
rect 44492 7522 44548 7532
rect 44604 7586 44660 7598
rect 44604 7534 44606 7586
rect 44658 7534 44660 7586
rect 44604 7476 44660 7534
rect 45164 7476 45220 7486
rect 44604 7474 45220 7476
rect 44604 7422 45166 7474
rect 45218 7422 45220 7474
rect 44604 7420 45220 7422
rect 45052 7252 45108 7262
rect 44380 7250 45108 7252
rect 44380 7198 45054 7250
rect 45106 7198 45108 7250
rect 44380 7196 45108 7198
rect 45052 7186 45108 7196
rect 44156 6972 45108 7028
rect 43932 6860 44324 6916
rect 44268 6802 44324 6860
rect 44268 6750 44270 6802
rect 44322 6750 44324 6802
rect 44268 6738 44324 6750
rect 44716 6690 44772 6702
rect 44716 6638 44718 6690
rect 44770 6638 44772 6690
rect 43708 6290 43764 6300
rect 44380 6468 44436 6478
rect 44380 6018 44436 6412
rect 44716 6130 44772 6638
rect 45052 6690 45108 6972
rect 45052 6638 45054 6690
rect 45106 6638 45108 6690
rect 45052 6626 45108 6638
rect 44940 6580 44996 6590
rect 44940 6486 44996 6524
rect 45164 6580 45220 7420
rect 45276 7476 45332 9102
rect 46396 9154 46452 10444
rect 46956 10164 47012 10556
rect 46956 10108 47124 10164
rect 46732 9268 46788 9278
rect 46396 9102 46398 9154
rect 46450 9102 46452 9154
rect 46396 9090 46452 9102
rect 46508 9266 46788 9268
rect 46508 9214 46734 9266
rect 46786 9214 46788 9266
rect 46508 9212 46788 9214
rect 47068 9268 47124 10108
rect 47180 9380 47236 10670
rect 47292 10722 47348 10780
rect 47292 10670 47294 10722
rect 47346 10670 47348 10722
rect 47292 10658 47348 10670
rect 48188 9938 48244 9950
rect 48188 9886 48190 9938
rect 48242 9886 48244 9938
rect 48188 9380 48244 9886
rect 47180 9324 48244 9380
rect 47068 9212 47348 9268
rect 45724 8932 45780 8942
rect 45612 8930 45780 8932
rect 45612 8878 45726 8930
rect 45778 8878 45780 8930
rect 45612 8876 45780 8878
rect 45388 8260 45444 8270
rect 45612 8260 45668 8876
rect 45724 8866 45780 8876
rect 46508 8484 46564 9212
rect 46732 9202 46788 9212
rect 47292 9154 47348 9212
rect 47404 9266 47460 9324
rect 47404 9214 47406 9266
rect 47458 9214 47460 9266
rect 47404 9202 47460 9214
rect 47292 9102 47294 9154
rect 47346 9102 47348 9154
rect 47292 9090 47348 9102
rect 46060 8428 46564 8484
rect 46620 9042 46676 9054
rect 46620 8990 46622 9042
rect 46674 8990 46676 9042
rect 46060 8370 46116 8428
rect 46060 8318 46062 8370
rect 46114 8318 46116 8370
rect 46060 8306 46116 8318
rect 45444 8204 45668 8260
rect 45388 8166 45444 8204
rect 45612 7698 45668 8204
rect 45612 7646 45614 7698
rect 45666 7646 45668 7698
rect 45612 7634 45668 7646
rect 46620 7698 46676 8990
rect 47068 9042 47124 9054
rect 47068 8990 47070 9042
rect 47122 8990 47124 9042
rect 47068 8820 47124 8990
rect 47852 9044 47908 9054
rect 47852 8950 47908 8988
rect 47964 8930 48020 8942
rect 47964 8878 47966 8930
rect 48018 8878 48020 8930
rect 47404 8820 47460 8830
rect 47068 8818 47460 8820
rect 47068 8766 47406 8818
rect 47458 8766 47460 8818
rect 47068 8764 47460 8766
rect 47404 8754 47460 8764
rect 47404 8372 47460 8382
rect 46620 7646 46622 7698
rect 46674 7646 46676 7698
rect 46620 7634 46676 7646
rect 46844 7700 46900 7710
rect 47404 7700 47460 8316
rect 46844 7698 47460 7700
rect 46844 7646 46846 7698
rect 46898 7646 47406 7698
rect 47458 7646 47460 7698
rect 46844 7644 47460 7646
rect 46844 7634 46900 7644
rect 47404 7634 47460 7644
rect 47852 7700 47908 7710
rect 47964 7700 48020 8878
rect 48188 8372 48244 8382
rect 48188 8278 48244 8316
rect 47852 7698 48020 7700
rect 47852 7646 47854 7698
rect 47906 7646 48020 7698
rect 47852 7644 48020 7646
rect 48188 7700 48244 7710
rect 47852 7634 47908 7644
rect 48188 7588 48244 7644
rect 48188 7586 48356 7588
rect 48188 7534 48190 7586
rect 48242 7534 48356 7586
rect 48188 7532 48356 7534
rect 48188 7522 48244 7532
rect 45276 7410 45332 7420
rect 46956 7476 47012 7486
rect 47292 7476 47348 7486
rect 46956 7382 47012 7420
rect 47180 7474 47348 7476
rect 47180 7422 47294 7474
rect 47346 7422 47348 7474
rect 47180 7420 47348 7422
rect 46956 6692 47012 6702
rect 46956 6598 47012 6636
rect 45164 6514 45220 6524
rect 45388 6578 45444 6590
rect 45388 6526 45390 6578
rect 45442 6526 45444 6578
rect 45388 6356 45444 6526
rect 46060 6580 46116 6590
rect 46060 6486 46116 6524
rect 46620 6578 46676 6590
rect 46620 6526 46622 6578
rect 46674 6526 46676 6578
rect 46172 6468 46228 6478
rect 46172 6374 46228 6412
rect 46396 6466 46452 6478
rect 46396 6414 46398 6466
rect 46450 6414 46452 6466
rect 45388 6290 45444 6300
rect 44716 6078 44718 6130
rect 44770 6078 44772 6130
rect 44716 6066 44772 6078
rect 44380 5966 44382 6018
rect 44434 5966 44436 6018
rect 44380 5954 44436 5966
rect 44492 6018 44548 6030
rect 44492 5966 44494 6018
rect 44546 5966 44548 6018
rect 43932 5796 43988 5806
rect 43932 5702 43988 5740
rect 42476 5182 42478 5234
rect 42530 5182 42532 5234
rect 42476 5170 42532 5182
rect 44492 5012 44548 5966
rect 46060 6020 46116 6030
rect 46060 5926 46116 5964
rect 44492 4946 44548 4956
rect 45276 5906 45332 5918
rect 45276 5854 45278 5906
rect 45330 5854 45332 5906
rect 45276 5236 45332 5854
rect 45388 5236 45444 5246
rect 45276 5234 45444 5236
rect 45276 5182 45390 5234
rect 45442 5182 45444 5234
rect 45276 5180 45444 5182
rect 42588 4900 42644 4910
rect 42588 4806 42644 4844
rect 43036 4898 43092 4910
rect 43036 4846 43038 4898
rect 43090 4846 43092 4898
rect 41580 4226 41860 4228
rect 41580 4174 41582 4226
rect 41634 4174 41860 4226
rect 41580 4172 41860 4174
rect 42588 4564 42644 4574
rect 43036 4564 43092 4846
rect 42644 4508 43092 4564
rect 43708 4900 43764 4910
rect 41580 4162 41636 4172
rect 39788 3614 39790 3666
rect 39842 3614 39844 3666
rect 39788 3602 39844 3614
rect 41916 4116 41972 4126
rect 41916 3666 41972 4060
rect 41916 3614 41918 3666
rect 41970 3614 41972 3666
rect 41916 3602 41972 3614
rect 42588 3668 42644 4508
rect 43708 4450 43764 4844
rect 43708 4398 43710 4450
rect 43762 4398 43764 4450
rect 43708 4386 43764 4398
rect 44156 4900 44212 4910
rect 44156 4340 44212 4844
rect 44940 4900 44996 4910
rect 44940 4564 44996 4844
rect 44940 4562 45108 4564
rect 44940 4510 44942 4562
rect 44994 4510 45108 4562
rect 44940 4508 45108 4510
rect 44940 4498 44996 4508
rect 44380 4340 44436 4350
rect 44156 4338 44436 4340
rect 44156 4286 44382 4338
rect 44434 4286 44436 4338
rect 44156 4284 44436 4286
rect 37884 3490 37940 3500
rect 42588 3554 42644 3612
rect 43820 3668 43876 3678
rect 44156 3668 44212 4284
rect 44380 4274 44436 4284
rect 45052 4340 45108 4508
rect 45276 4340 45332 5180
rect 45388 5170 45444 5180
rect 46396 5124 46452 6414
rect 46620 6356 46676 6526
rect 47180 6580 47236 7420
rect 47292 7410 47348 7420
rect 47516 7476 47572 7486
rect 47404 7252 47460 7262
rect 47292 7250 47460 7252
rect 47292 7198 47406 7250
rect 47458 7198 47460 7250
rect 47292 7196 47460 7198
rect 47292 6690 47348 7196
rect 47404 7186 47460 7196
rect 47292 6638 47294 6690
rect 47346 6638 47348 6690
rect 47292 6626 47348 6638
rect 47180 6514 47236 6524
rect 47516 6578 47572 7420
rect 48300 6802 48356 7532
rect 48300 6750 48302 6802
rect 48354 6750 48356 6802
rect 48300 6738 48356 6750
rect 47852 6692 47908 6702
rect 47852 6598 47908 6636
rect 47516 6526 47518 6578
rect 47570 6526 47572 6578
rect 46620 6290 46676 6300
rect 46956 6466 47012 6478
rect 46956 6414 46958 6466
rect 47010 6414 47012 6466
rect 46956 6020 47012 6414
rect 46956 5954 47012 5964
rect 47068 6356 47124 6366
rect 46508 5124 46564 5134
rect 46396 5122 46564 5124
rect 46396 5070 46510 5122
rect 46562 5070 46564 5122
rect 46396 5068 46564 5070
rect 46508 5058 46564 5068
rect 46956 5124 47012 5134
rect 46956 5030 47012 5068
rect 47068 5122 47124 6300
rect 47068 5070 47070 5122
rect 47122 5070 47124 5122
rect 47068 5058 47124 5070
rect 47516 5122 47572 6526
rect 47628 6468 47684 6478
rect 47628 6374 47684 6412
rect 48188 6468 48244 6478
rect 48188 5794 48244 6412
rect 48188 5742 48190 5794
rect 48242 5742 48244 5794
rect 48188 5730 48244 5742
rect 47516 5070 47518 5122
rect 47570 5070 47572 5122
rect 47516 5058 47572 5070
rect 47852 5124 47908 5134
rect 47852 5030 47908 5068
rect 47628 5012 47684 5022
rect 47628 4918 47684 4956
rect 48188 5012 48244 5022
rect 46732 4900 46788 4910
rect 46060 4898 46788 4900
rect 46060 4846 46734 4898
rect 46786 4846 46788 4898
rect 46060 4844 46788 4846
rect 46060 4450 46116 4844
rect 46732 4834 46788 4844
rect 46060 4398 46062 4450
rect 46114 4398 46116 4450
rect 46060 4386 46116 4398
rect 45052 4338 45332 4340
rect 45052 4286 45278 4338
rect 45330 4286 45332 4338
rect 45052 4284 45332 4286
rect 43876 3612 44212 3668
rect 45052 3666 45108 4284
rect 45276 4274 45332 4284
rect 48188 4226 48244 4956
rect 48188 4174 48190 4226
rect 48242 4174 48244 4226
rect 48188 4162 48244 4174
rect 45052 3614 45054 3666
rect 45106 3614 45108 3666
rect 43820 3574 43876 3612
rect 45052 3602 45108 3614
rect 42588 3502 42590 3554
rect 42642 3502 42644 3554
rect 42588 3490 42644 3502
rect 47628 3556 47684 3566
rect 46956 3444 47012 3482
rect 47628 3462 47684 3500
rect 46956 3378 47012 3388
rect 48076 3444 48132 3454
rect 48188 3444 48244 3482
rect 48132 3442 48244 3444
rect 48132 3390 48190 3442
rect 48242 3390 48244 3442
rect 48132 3388 48244 3390
rect 48076 3378 48132 3388
rect 48188 2772 48244 3388
rect 48188 2706 48244 2716
rect 34468 2604 34580 2660
rect 34412 2594 34468 2604
rect 32284 2258 32340 2268
rect 30380 1474 30436 1484
rect 25788 1250 25844 1260
<< via2 >>
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 5628 45612 5684 45668
rect 7980 45388 8036 45444
rect 8540 45388 8596 45444
rect 3276 44380 3332 44436
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4732 44434 4788 44436
rect 4732 44382 4734 44434
rect 4734 44382 4786 44434
rect 4786 44382 4788 44434
rect 4732 44380 4788 44382
rect 3500 43708 3556 43764
rect 3276 43596 3332 43652
rect 1932 43260 1988 43316
rect 4844 43650 4900 43652
rect 4844 43598 4846 43650
rect 4846 43598 4898 43650
rect 4898 43598 4900 43650
rect 4844 43596 4900 43598
rect 3388 42812 3444 42868
rect 1708 42476 1764 42532
rect 1708 41468 1764 41524
rect 1372 41356 1428 41412
rect 1932 39340 1988 39396
rect 1484 37436 1540 37492
rect 1708 34636 1764 34692
rect 1820 34748 1876 34804
rect 2268 42476 2324 42532
rect 3500 42588 3556 42644
rect 3612 43260 3668 43316
rect 3164 42476 3220 42532
rect 2828 42364 2884 42420
rect 2380 40348 2436 40404
rect 2604 40514 2660 40516
rect 2604 40462 2606 40514
rect 2606 40462 2658 40514
rect 2658 40462 2660 40514
rect 2604 40460 2660 40462
rect 3388 40514 3444 40516
rect 3388 40462 3390 40514
rect 3390 40462 3442 40514
rect 3442 40462 3444 40514
rect 3388 40460 3444 40462
rect 3164 40402 3220 40404
rect 3164 40350 3166 40402
rect 3166 40350 3218 40402
rect 3218 40350 3220 40402
rect 3164 40348 3220 40350
rect 3724 42866 3780 42868
rect 3724 42814 3726 42866
rect 3726 42814 3778 42866
rect 3778 42814 3780 42866
rect 3724 42812 3780 42814
rect 4508 43260 4564 43316
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4844 42924 4900 42980
rect 3612 39340 3668 39396
rect 4732 42588 4788 42644
rect 6188 44434 6244 44436
rect 6188 44382 6190 44434
rect 6190 44382 6242 44434
rect 6242 44382 6244 44434
rect 6188 44380 6244 44382
rect 7756 44322 7812 44324
rect 7756 44270 7758 44322
rect 7758 44270 7810 44322
rect 7810 44270 7812 44322
rect 7756 44268 7812 44270
rect 7756 44044 7812 44100
rect 7308 43762 7364 43764
rect 7308 43710 7310 43762
rect 7310 43710 7362 43762
rect 7362 43710 7364 43762
rect 7308 43708 7364 43710
rect 5740 43426 5796 43428
rect 5740 43374 5742 43426
rect 5742 43374 5794 43426
rect 5794 43374 5796 43426
rect 5740 43372 5796 43374
rect 6300 42978 6356 42980
rect 6300 42926 6302 42978
rect 6302 42926 6354 42978
rect 6354 42926 6356 42978
rect 6300 42924 6356 42926
rect 6636 42924 6692 42980
rect 8428 44268 8484 44324
rect 8204 44156 8260 44212
rect 8092 43708 8148 43764
rect 6748 43372 6804 43428
rect 5740 42642 5796 42644
rect 5740 42590 5742 42642
rect 5742 42590 5794 42642
rect 5794 42590 5796 42642
rect 5740 42588 5796 42590
rect 6300 42530 6356 42532
rect 6300 42478 6302 42530
rect 6302 42478 6354 42530
rect 6354 42478 6356 42530
rect 6300 42476 6356 42478
rect 6748 42588 6804 42644
rect 7196 42476 7252 42532
rect 6412 42364 6468 42420
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 3836 41244 3892 41300
rect 4620 41298 4676 41300
rect 4620 41246 4622 41298
rect 4622 41246 4674 41298
rect 4674 41246 4676 41298
rect 4620 41244 4676 41246
rect 4732 40908 4788 40964
rect 5740 42028 5796 42084
rect 7308 41804 7364 41860
rect 7644 42476 7700 42532
rect 9436 45666 9492 45668
rect 9436 45614 9438 45666
rect 9438 45614 9490 45666
rect 9490 45614 9492 45666
rect 9436 45612 9492 45614
rect 9548 45388 9604 45444
rect 13020 45724 13076 45780
rect 11340 45666 11396 45668
rect 11340 45614 11342 45666
rect 11342 45614 11394 45666
rect 11394 45614 11396 45666
rect 11340 45612 11396 45614
rect 10892 45388 10948 45444
rect 13916 45778 13972 45780
rect 13916 45726 13918 45778
rect 13918 45726 13970 45778
rect 13970 45726 13972 45778
rect 13916 45724 13972 45726
rect 14588 45724 14644 45780
rect 13132 45612 13188 45668
rect 14028 45276 14084 45332
rect 9660 44322 9716 44324
rect 9660 44270 9662 44322
rect 9662 44270 9714 44322
rect 9714 44270 9716 44322
rect 9660 44268 9716 44270
rect 9548 44210 9604 44212
rect 9548 44158 9550 44210
rect 9550 44158 9602 44210
rect 9602 44158 9604 44210
rect 9548 44156 9604 44158
rect 8652 42700 8708 42756
rect 8764 42028 8820 42084
rect 8540 41916 8596 41972
rect 8092 41692 8148 41748
rect 9660 43148 9716 43204
rect 9660 42700 9716 42756
rect 10892 44044 10948 44100
rect 12684 44044 12740 44100
rect 12684 43820 12740 43876
rect 13020 43762 13076 43764
rect 13020 43710 13022 43762
rect 13022 43710 13074 43762
rect 13074 43710 13076 43762
rect 13020 43708 13076 43710
rect 14588 45052 14644 45108
rect 13356 43820 13412 43876
rect 12460 43650 12516 43652
rect 12460 43598 12462 43650
rect 12462 43598 12514 43650
rect 12514 43598 12516 43650
rect 12460 43596 12516 43598
rect 10108 43148 10164 43204
rect 10780 43148 10836 43204
rect 10332 42588 10388 42644
rect 9548 42140 9604 42196
rect 9436 41804 9492 41860
rect 5852 40962 5908 40964
rect 5852 40910 5854 40962
rect 5854 40910 5906 40962
rect 5906 40910 5908 40962
rect 5852 40908 5908 40910
rect 7084 40908 7140 40964
rect 3836 40460 3892 40516
rect 3164 38834 3220 38836
rect 3164 38782 3166 38834
rect 3166 38782 3218 38834
rect 3218 38782 3220 38834
rect 3164 38780 3220 38782
rect 3388 38722 3444 38724
rect 3388 38670 3390 38722
rect 3390 38670 3442 38722
rect 3442 38670 3444 38722
rect 3388 38668 3444 38670
rect 2156 38220 2212 38276
rect 3164 38162 3220 38164
rect 3164 38110 3166 38162
rect 3166 38110 3218 38162
rect 3218 38110 3220 38162
rect 3164 38108 3220 38110
rect 3388 38108 3444 38164
rect 2492 37154 2548 37156
rect 2492 37102 2494 37154
rect 2494 37102 2546 37154
rect 2546 37102 2548 37154
rect 2492 37100 2548 37102
rect 2156 36988 2212 37044
rect 1932 34412 1988 34468
rect 2492 36204 2548 36260
rect 2268 35084 2324 35140
rect 1708 33234 1764 33236
rect 1708 33182 1710 33234
rect 1710 33182 1762 33234
rect 1762 33182 1764 33234
rect 1708 33180 1764 33182
rect 1932 33964 1988 34020
rect 2716 35084 2772 35140
rect 2828 34188 2884 34244
rect 2380 33628 2436 33684
rect 2044 33122 2100 33124
rect 2044 33070 2046 33122
rect 2046 33070 2098 33122
rect 2098 33070 2100 33122
rect 2044 33068 2100 33070
rect 2268 32956 2324 33012
rect 1708 31836 1764 31892
rect 2044 32172 2100 32228
rect 2268 32060 2324 32116
rect 2492 31948 2548 32004
rect 1932 30322 1988 30324
rect 1932 30270 1934 30322
rect 1934 30270 1986 30322
rect 1986 30270 1988 30322
rect 1932 30268 1988 30270
rect 2156 31164 2212 31220
rect 2380 31554 2436 31556
rect 2380 31502 2382 31554
rect 2382 31502 2434 31554
rect 2434 31502 2436 31554
rect 2380 31500 2436 31502
rect 1820 29820 1876 29876
rect 2044 30098 2100 30100
rect 2044 30046 2046 30098
rect 2046 30046 2098 30098
rect 2098 30046 2100 30098
rect 2044 30044 2100 30046
rect 1932 29036 1988 29092
rect 1820 28476 1876 28532
rect 1484 26684 1540 26740
rect 1596 28252 1652 28308
rect 2156 28700 2212 28756
rect 1820 28028 1876 28084
rect 1708 26236 1764 26292
rect 1484 25116 1540 25172
rect 1372 22092 1428 22148
rect 1596 24892 1652 24948
rect 1484 21980 1540 22036
rect 1148 21308 1204 21364
rect 1036 19852 1092 19908
rect 1260 18844 1316 18900
rect 1484 17164 1540 17220
rect 2380 29036 2436 29092
rect 3052 34748 3108 34804
rect 2940 33516 2996 33572
rect 3388 34636 3444 34692
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 4172 38834 4228 38836
rect 4172 38782 4174 38834
rect 4174 38782 4226 38834
rect 4226 38782 4228 38834
rect 4172 38780 4228 38782
rect 5068 39394 5124 39396
rect 5068 39342 5070 39394
rect 5070 39342 5122 39394
rect 5122 39342 5124 39394
rect 5068 39340 5124 39342
rect 4508 38780 4564 38836
rect 4844 38780 4900 38836
rect 4396 38668 4452 38724
rect 4956 38668 5012 38724
rect 5628 39340 5684 39396
rect 6860 38892 6916 38948
rect 5180 38556 5236 38612
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 5852 38444 5908 38500
rect 5068 38162 5124 38164
rect 5068 38110 5070 38162
rect 5070 38110 5122 38162
rect 5122 38110 5124 38162
rect 5068 38108 5124 38110
rect 3500 37436 3556 37492
rect 3276 33516 3332 33572
rect 3948 36428 4004 36484
rect 4284 37212 4340 37268
rect 4732 37772 4788 37828
rect 5292 37772 5348 37828
rect 4732 37436 4788 37492
rect 5180 37436 5236 37492
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4396 36482 4452 36484
rect 4396 36430 4398 36482
rect 4398 36430 4450 36482
rect 4450 36430 4452 36482
rect 4396 36428 4452 36430
rect 4844 36316 4900 36372
rect 5516 37772 5572 37828
rect 6972 39004 7028 39060
rect 8316 41186 8372 41188
rect 8316 41134 8318 41186
rect 8318 41134 8370 41186
rect 8370 41134 8372 41186
rect 8316 41132 8372 41134
rect 7756 40908 7812 40964
rect 7532 40124 7588 40180
rect 7532 38780 7588 38836
rect 6636 38444 6692 38500
rect 5516 37266 5572 37268
rect 5516 37214 5518 37266
rect 5518 37214 5570 37266
rect 5570 37214 5572 37266
rect 5516 37212 5572 37214
rect 5852 37212 5908 37268
rect 5292 36988 5348 37044
rect 5180 36876 5236 36932
rect 5404 36876 5460 36932
rect 5292 36764 5348 36820
rect 5068 36428 5124 36484
rect 5068 36092 5124 36148
rect 5964 37154 6020 37156
rect 5964 37102 5966 37154
rect 5966 37102 6018 37154
rect 6018 37102 6020 37154
rect 5964 37100 6020 37102
rect 7084 38050 7140 38052
rect 7084 37998 7086 38050
rect 7086 37998 7138 38050
rect 7138 37998 7140 38050
rect 7084 37996 7140 37998
rect 7644 38444 7700 38500
rect 6860 37212 6916 37268
rect 6188 36988 6244 37044
rect 6188 36428 6244 36484
rect 5852 36370 5908 36372
rect 5852 36318 5854 36370
rect 5854 36318 5906 36370
rect 5906 36318 5908 36370
rect 5852 36316 5908 36318
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 3724 35084 3780 35140
rect 5740 35308 5796 35364
rect 5180 34860 5236 34916
rect 4172 34802 4228 34804
rect 4172 34750 4174 34802
rect 4174 34750 4226 34802
rect 4226 34750 4228 34802
rect 4172 34748 4228 34750
rect 4620 34690 4676 34692
rect 4620 34638 4622 34690
rect 4622 34638 4674 34690
rect 4674 34638 4676 34690
rect 4620 34636 4676 34638
rect 5180 34690 5236 34692
rect 5180 34638 5182 34690
rect 5182 34638 5234 34690
rect 5234 34638 5236 34690
rect 5180 34636 5236 34638
rect 5068 34188 5124 34244
rect 4844 34076 4900 34132
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 5628 34914 5684 34916
rect 5628 34862 5630 34914
rect 5630 34862 5682 34914
rect 5682 34862 5684 34914
rect 5628 34860 5684 34862
rect 6412 36258 6468 36260
rect 6412 36206 6414 36258
rect 6414 36206 6466 36258
rect 6466 36206 6468 36258
rect 6412 36204 6468 36206
rect 6300 35756 6356 35812
rect 7196 36482 7252 36484
rect 7196 36430 7198 36482
rect 7198 36430 7250 36482
rect 7250 36430 7252 36482
rect 7196 36428 7252 36430
rect 6524 35868 6580 35924
rect 6636 36316 6692 36372
rect 7420 36370 7476 36372
rect 7420 36318 7422 36370
rect 7422 36318 7474 36370
rect 7474 36318 7476 36370
rect 7420 36316 7476 36318
rect 7644 37490 7700 37492
rect 7644 37438 7646 37490
rect 7646 37438 7698 37490
rect 7698 37438 7700 37490
rect 7644 37436 7700 37438
rect 7532 36204 7588 36260
rect 7644 35922 7700 35924
rect 7644 35870 7646 35922
rect 7646 35870 7698 35922
rect 7698 35870 7700 35922
rect 7644 35868 7700 35870
rect 7084 35810 7140 35812
rect 7084 35758 7086 35810
rect 7086 35758 7138 35810
rect 7138 35758 7140 35810
rect 7084 35756 7140 35758
rect 8316 40796 8372 40852
rect 8428 39340 8484 39396
rect 8092 39058 8148 39060
rect 8092 39006 8094 39058
rect 8094 39006 8146 39058
rect 8146 39006 8148 39058
rect 8092 39004 8148 39006
rect 8316 38946 8372 38948
rect 8316 38894 8318 38946
rect 8318 38894 8370 38946
rect 8370 38894 8372 38946
rect 8316 38892 8372 38894
rect 8204 38834 8260 38836
rect 8204 38782 8206 38834
rect 8206 38782 8258 38834
rect 8258 38782 8260 38834
rect 8204 38780 8260 38782
rect 8988 39452 9044 39508
rect 8540 39004 8596 39060
rect 8652 38892 8708 38948
rect 6524 35308 6580 35364
rect 6076 34412 6132 34468
rect 5628 34130 5684 34132
rect 5628 34078 5630 34130
rect 5630 34078 5682 34130
rect 5682 34078 5684 34130
rect 5628 34076 5684 34078
rect 3164 32844 3220 32900
rect 3052 32674 3108 32676
rect 3052 32622 3054 32674
rect 3054 32622 3106 32674
rect 3106 32622 3108 32674
rect 3052 32620 3108 32622
rect 2828 32562 2884 32564
rect 2828 32510 2830 32562
rect 2830 32510 2882 32562
rect 2882 32510 2884 32562
rect 2828 32508 2884 32510
rect 3164 31948 3220 32004
rect 2828 31778 2884 31780
rect 2828 31726 2830 31778
rect 2830 31726 2882 31778
rect 2882 31726 2884 31778
rect 2828 31724 2884 31726
rect 3164 31612 3220 31668
rect 3388 32060 3444 32116
rect 3276 31388 3332 31444
rect 3388 31276 3444 31332
rect 2940 30210 2996 30212
rect 2940 30158 2942 30210
rect 2942 30158 2994 30210
rect 2994 30158 2996 30210
rect 2940 30156 2996 30158
rect 3836 32956 3892 33012
rect 4172 32956 4228 33012
rect 3836 32674 3892 32676
rect 3836 32622 3838 32674
rect 3838 32622 3890 32674
rect 3890 32622 3892 32674
rect 3836 32620 3892 32622
rect 3948 32396 4004 32452
rect 3612 31724 3668 31780
rect 3948 32060 4004 32116
rect 3724 31666 3780 31668
rect 3724 31614 3726 31666
rect 3726 31614 3778 31666
rect 3778 31614 3780 31666
rect 3724 31612 3780 31614
rect 3836 31554 3892 31556
rect 3836 31502 3838 31554
rect 3838 31502 3890 31554
rect 3890 31502 3892 31554
rect 3836 31500 3892 31502
rect 4060 31164 4116 31220
rect 4956 32732 5012 32788
rect 5068 32620 5124 32676
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4844 31948 4900 32004
rect 4508 31500 4564 31556
rect 4732 31554 4788 31556
rect 4732 31502 4734 31554
rect 4734 31502 4786 31554
rect 4786 31502 4788 31554
rect 4732 31500 4788 31502
rect 4508 31276 4564 31332
rect 4396 31052 4452 31108
rect 3724 30268 3780 30324
rect 2492 28812 2548 28868
rect 2604 28476 2660 28532
rect 4060 30098 4116 30100
rect 4060 30046 4062 30098
rect 4062 30046 4114 30098
rect 4114 30046 4116 30098
rect 4060 30044 4116 30046
rect 2604 28028 2660 28084
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4956 31612 5012 31668
rect 5068 31388 5124 31444
rect 5628 33516 5684 33572
rect 5628 32844 5684 32900
rect 6076 33852 6132 33908
rect 6412 33516 6468 33572
rect 6636 33852 6692 33908
rect 5964 32620 6020 32676
rect 5964 31724 6020 31780
rect 5852 31666 5908 31668
rect 5852 31614 5854 31666
rect 5854 31614 5906 31666
rect 5906 31614 5908 31666
rect 5852 31612 5908 31614
rect 6076 31612 6132 31668
rect 5292 31388 5348 31444
rect 6076 31164 6132 31220
rect 5180 30994 5236 30996
rect 5180 30942 5182 30994
rect 5182 30942 5234 30994
rect 5234 30942 5236 30994
rect 5180 30940 5236 30942
rect 4284 30156 4340 30212
rect 4956 30322 5012 30324
rect 4956 30270 4958 30322
rect 4958 30270 5010 30322
rect 5010 30270 5012 30322
rect 4956 30268 5012 30270
rect 4844 30156 4900 30212
rect 4732 29148 4788 29204
rect 3500 27804 3556 27860
rect 2156 25564 2212 25620
rect 2156 25116 2212 25172
rect 1708 19346 1764 19348
rect 1708 19294 1710 19346
rect 1710 19294 1762 19346
rect 1762 19294 1764 19346
rect 1708 19292 1764 19294
rect 2044 21644 2100 21700
rect 1932 21474 1988 21476
rect 1932 21422 1934 21474
rect 1934 21422 1986 21474
rect 1986 21422 1988 21474
rect 1932 21420 1988 21422
rect 2716 24722 2772 24724
rect 2716 24670 2718 24722
rect 2718 24670 2770 24722
rect 2770 24670 2772 24722
rect 2716 24668 2772 24670
rect 2940 24834 2996 24836
rect 2940 24782 2942 24834
rect 2942 24782 2994 24834
rect 2994 24782 2996 24834
rect 2940 24780 2996 24782
rect 2604 23884 2660 23940
rect 2492 23436 2548 23492
rect 2380 23324 2436 23380
rect 2268 21420 2324 21476
rect 2156 19906 2212 19908
rect 2156 19854 2158 19906
rect 2158 19854 2210 19906
rect 2210 19854 2212 19906
rect 2156 19852 2212 19854
rect 1820 18060 1876 18116
rect 1932 19404 1988 19460
rect 2044 18450 2100 18452
rect 2044 18398 2046 18450
rect 2046 18398 2098 18450
rect 2098 18398 2100 18450
rect 2044 18396 2100 18398
rect 1036 15148 1092 15204
rect 1372 14364 1428 14420
rect 1484 13916 1540 13972
rect 2380 18956 2436 19012
rect 2268 16882 2324 16884
rect 2268 16830 2270 16882
rect 2270 16830 2322 16882
rect 2322 16830 2324 16882
rect 2268 16828 2324 16830
rect 2492 18450 2548 18452
rect 2492 18398 2494 18450
rect 2494 18398 2546 18450
rect 2546 18398 2548 18450
rect 2492 18396 2548 18398
rect 2828 24108 2884 24164
rect 3388 24722 3444 24724
rect 3388 24670 3390 24722
rect 3390 24670 3442 24722
rect 3442 24670 3444 24722
rect 3388 24668 3444 24670
rect 3164 24108 3220 24164
rect 3052 23996 3108 24052
rect 4844 29260 4900 29316
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4508 28866 4564 28868
rect 4508 28814 4510 28866
rect 4510 28814 4562 28866
rect 4562 28814 4564 28866
rect 4508 28812 4564 28814
rect 4172 27804 4228 27860
rect 4284 28588 4340 28644
rect 3164 23660 3220 23716
rect 4508 28476 4564 28532
rect 4844 27916 4900 27972
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 3836 24834 3892 24836
rect 3836 24782 3838 24834
rect 3838 24782 3890 24834
rect 3890 24782 3892 24834
rect 3836 24780 3892 24782
rect 3612 23324 3668 23380
rect 3724 24668 3780 24724
rect 2716 20860 2772 20916
rect 2716 18732 2772 18788
rect 3276 20972 3332 21028
rect 3948 23436 4004 23492
rect 3948 22482 4004 22484
rect 3948 22430 3950 22482
rect 3950 22430 4002 22482
rect 4002 22430 4004 22482
rect 3948 22428 4004 22430
rect 4844 26460 4900 26516
rect 4620 26290 4676 26292
rect 4620 26238 4622 26290
rect 4622 26238 4674 26290
rect 4674 26238 4676 26290
rect 4620 26236 4676 26238
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4620 25618 4676 25620
rect 4620 25566 4622 25618
rect 4622 25566 4674 25618
rect 4674 25566 4676 25618
rect 4620 25564 4676 25566
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4284 24108 4340 24164
rect 5292 29538 5348 29540
rect 5292 29486 5294 29538
rect 5294 29486 5346 29538
rect 5346 29486 5348 29538
rect 5292 29484 5348 29486
rect 5068 29148 5124 29204
rect 5068 28476 5124 28532
rect 6076 30268 6132 30324
rect 5852 30156 5908 30212
rect 5628 29202 5684 29204
rect 5628 29150 5630 29202
rect 5630 29150 5682 29202
rect 5682 29150 5684 29202
rect 5628 29148 5684 29150
rect 5516 28140 5572 28196
rect 5180 27580 5236 27636
rect 5068 27132 5124 27188
rect 5404 27020 5460 27076
rect 5516 26908 5572 26964
rect 5852 28924 5908 28980
rect 6412 31612 6468 31668
rect 6524 31164 6580 31220
rect 6524 30994 6580 30996
rect 6524 30942 6526 30994
rect 6526 30942 6578 30994
rect 6578 30942 6580 30994
rect 6524 30940 6580 30942
rect 6524 30716 6580 30772
rect 6076 29426 6132 29428
rect 6076 29374 6078 29426
rect 6078 29374 6130 29426
rect 6130 29374 6132 29426
rect 6076 29372 6132 29374
rect 6076 28642 6132 28644
rect 6076 28590 6078 28642
rect 6078 28590 6130 28642
rect 6130 28590 6132 28642
rect 6076 28588 6132 28590
rect 7196 34860 7252 34916
rect 7420 34524 7476 34580
rect 7980 37996 8036 38052
rect 8764 37772 8820 37828
rect 8428 37324 8484 37380
rect 8204 36482 8260 36484
rect 8204 36430 8206 36482
rect 8206 36430 8258 36482
rect 8258 36430 8260 36482
rect 8204 36428 8260 36430
rect 8092 36092 8148 36148
rect 8204 36204 8260 36260
rect 9660 41916 9716 41972
rect 10108 41692 10164 41748
rect 10220 41132 10276 41188
rect 9772 40962 9828 40964
rect 9772 40910 9774 40962
rect 9774 40910 9826 40962
rect 9826 40910 9828 40962
rect 9772 40908 9828 40910
rect 10668 41298 10724 41300
rect 10668 41246 10670 41298
rect 10670 41246 10722 41298
rect 10722 41246 10724 41298
rect 10668 41244 10724 41246
rect 13916 43650 13972 43652
rect 13916 43598 13918 43650
rect 13918 43598 13970 43650
rect 13970 43598 13972 43650
rect 13916 43596 13972 43598
rect 11788 43036 11844 43092
rect 10668 40796 10724 40852
rect 10108 40460 10164 40516
rect 11676 42140 11732 42196
rect 11564 41356 11620 41412
rect 11676 40908 11732 40964
rect 12796 42588 12852 42644
rect 12124 42530 12180 42532
rect 12124 42478 12126 42530
rect 12126 42478 12178 42530
rect 12178 42478 12180 42530
rect 12124 42476 12180 42478
rect 12012 41244 12068 41300
rect 12348 41132 12404 41188
rect 12460 41356 12516 41412
rect 11564 40796 11620 40852
rect 12236 40962 12292 40964
rect 12236 40910 12238 40962
rect 12238 40910 12290 40962
rect 12290 40910 12292 40962
rect 12236 40908 12292 40910
rect 12684 41244 12740 41300
rect 14140 43484 14196 43540
rect 13580 43036 13636 43092
rect 13580 42530 13636 42532
rect 13580 42478 13582 42530
rect 13582 42478 13634 42530
rect 13634 42478 13636 42530
rect 13580 42476 13636 42478
rect 13468 41746 13524 41748
rect 13468 41694 13470 41746
rect 13470 41694 13522 41746
rect 13522 41694 13524 41746
rect 13468 41692 13524 41694
rect 13468 41186 13524 41188
rect 13468 41134 13470 41186
rect 13470 41134 13522 41186
rect 13522 41134 13524 41186
rect 13468 41132 13524 41134
rect 13916 42700 13972 42756
rect 14140 42588 14196 42644
rect 15372 44546 15428 44548
rect 15372 44494 15374 44546
rect 15374 44494 15426 44546
rect 15426 44494 15428 44546
rect 15372 44492 15428 44494
rect 20860 46060 20916 46116
rect 22092 46114 22148 46116
rect 22092 46062 22094 46114
rect 22094 46062 22146 46114
rect 22146 46062 22148 46114
rect 22092 46060 22148 46062
rect 22428 46060 22484 46116
rect 16940 45778 16996 45780
rect 16940 45726 16942 45778
rect 16942 45726 16994 45778
rect 16994 45726 16996 45778
rect 16940 45724 16996 45726
rect 17500 45106 17556 45108
rect 17500 45054 17502 45106
rect 17502 45054 17554 45106
rect 17554 45054 17556 45106
rect 17500 45052 17556 45054
rect 16156 44492 16212 44548
rect 16828 44044 16884 44100
rect 14700 43650 14756 43652
rect 14700 43598 14702 43650
rect 14702 43598 14754 43650
rect 14754 43598 14756 43650
rect 14700 43596 14756 43598
rect 15372 43650 15428 43652
rect 15372 43598 15374 43650
rect 15374 43598 15426 43650
rect 15426 43598 15428 43650
rect 15372 43596 15428 43598
rect 15260 43538 15316 43540
rect 15260 43486 15262 43538
rect 15262 43486 15314 43538
rect 15314 43486 15316 43538
rect 15260 43484 15316 43486
rect 14924 43426 14980 43428
rect 14924 43374 14926 43426
rect 14926 43374 14978 43426
rect 14978 43374 14980 43426
rect 14924 43372 14980 43374
rect 15484 43260 15540 43316
rect 14588 42754 14644 42756
rect 14588 42702 14590 42754
rect 14590 42702 14642 42754
rect 14642 42702 14644 42754
rect 14588 42700 14644 42702
rect 15484 42700 15540 42756
rect 16156 43538 16212 43540
rect 16156 43486 16158 43538
rect 16158 43486 16210 43538
rect 16210 43486 16212 43538
rect 16156 43484 16212 43486
rect 16268 43426 16324 43428
rect 16268 43374 16270 43426
rect 16270 43374 16322 43426
rect 16322 43374 16324 43426
rect 16268 43372 16324 43374
rect 16380 43260 16436 43316
rect 16940 43260 16996 43316
rect 15708 42924 15764 42980
rect 12684 40684 12740 40740
rect 10892 40514 10948 40516
rect 10892 40462 10894 40514
rect 10894 40462 10946 40514
rect 10946 40462 10948 40514
rect 10892 40460 10948 40462
rect 9884 40348 9940 40404
rect 9772 40178 9828 40180
rect 9772 40126 9774 40178
rect 9774 40126 9826 40178
rect 9826 40126 9828 40178
rect 9772 40124 9828 40126
rect 9660 39730 9716 39732
rect 9660 39678 9662 39730
rect 9662 39678 9714 39730
rect 9714 39678 9716 39730
rect 9660 39676 9716 39678
rect 9996 40124 10052 40180
rect 12012 40514 12068 40516
rect 12012 40462 12014 40514
rect 12014 40462 12066 40514
rect 12066 40462 12068 40514
rect 12012 40460 12068 40462
rect 11004 40348 11060 40404
rect 9548 39452 9604 39508
rect 9324 39340 9380 39396
rect 9212 39004 9268 39060
rect 8988 37324 9044 37380
rect 9100 37548 9156 37604
rect 8876 36764 8932 36820
rect 9660 38946 9716 38948
rect 9660 38894 9662 38946
rect 9662 38894 9714 38946
rect 9714 38894 9716 38946
rect 9660 38892 9716 38894
rect 9548 38668 9604 38724
rect 10780 39676 10836 39732
rect 10332 39506 10388 39508
rect 10332 39454 10334 39506
rect 10334 39454 10386 39506
rect 10386 39454 10388 39506
rect 10332 39452 10388 39454
rect 9884 39340 9940 39396
rect 10108 38780 10164 38836
rect 9324 37826 9380 37828
rect 9324 37774 9326 37826
rect 9326 37774 9378 37826
rect 9378 37774 9380 37826
rect 9324 37772 9380 37774
rect 9548 37772 9604 37828
rect 9660 37548 9716 37604
rect 8764 36428 8820 36484
rect 8652 36204 8708 36260
rect 9212 36482 9268 36484
rect 9212 36430 9214 36482
rect 9214 36430 9266 36482
rect 9266 36430 9268 36482
rect 9212 36428 9268 36430
rect 8540 35420 8596 35476
rect 8204 34748 8260 34804
rect 7084 34076 7140 34132
rect 6972 32620 7028 32676
rect 7756 33964 7812 34020
rect 7420 33180 7476 33236
rect 7084 31724 7140 31780
rect 7196 31666 7252 31668
rect 7196 31614 7198 31666
rect 7198 31614 7250 31666
rect 7250 31614 7252 31666
rect 7196 31612 7252 31614
rect 6860 31500 6916 31556
rect 7196 31388 7252 31444
rect 6860 31052 6916 31108
rect 6636 30156 6692 30212
rect 6972 30940 7028 30996
rect 7084 30210 7140 30212
rect 7084 30158 7086 30210
rect 7086 30158 7138 30210
rect 7138 30158 7140 30210
rect 7084 30156 7140 30158
rect 8092 34130 8148 34132
rect 8092 34078 8094 34130
rect 8094 34078 8146 34130
rect 8146 34078 8148 34130
rect 8092 34076 8148 34078
rect 8316 33852 8372 33908
rect 7980 33458 8036 33460
rect 7980 33406 7982 33458
rect 7982 33406 8034 33458
rect 8034 33406 8036 33458
rect 7980 33404 8036 33406
rect 7420 31500 7476 31556
rect 7532 31276 7588 31332
rect 6636 29708 6692 29764
rect 6300 28700 6356 28756
rect 6524 28588 6580 28644
rect 6076 28140 6132 28196
rect 8540 34524 8596 34580
rect 8428 32172 8484 32228
rect 8540 32060 8596 32116
rect 7868 31164 7924 31220
rect 7084 28700 7140 28756
rect 6972 28418 7028 28420
rect 6972 28366 6974 28418
rect 6974 28366 7026 28418
rect 7026 28366 7028 28418
rect 6972 28364 7028 28366
rect 6748 27970 6804 27972
rect 6748 27918 6750 27970
rect 6750 27918 6802 27970
rect 6802 27918 6804 27970
rect 6748 27916 6804 27918
rect 6860 27132 6916 27188
rect 5068 25282 5124 25284
rect 5068 25230 5070 25282
rect 5070 25230 5122 25282
rect 5122 25230 5124 25282
rect 5068 25228 5124 25230
rect 6972 27074 7028 27076
rect 6972 27022 6974 27074
rect 6974 27022 7026 27074
rect 7026 27022 7028 27074
rect 6972 27020 7028 27022
rect 5964 26962 6020 26964
rect 5964 26910 5966 26962
rect 5966 26910 6018 26962
rect 6018 26910 6020 26962
rect 5964 26908 6020 26910
rect 5852 26236 5908 26292
rect 6076 26684 6132 26740
rect 6300 26402 6356 26404
rect 6300 26350 6302 26402
rect 6302 26350 6354 26402
rect 6354 26350 6356 26402
rect 6300 26348 6356 26350
rect 5740 26124 5796 26180
rect 5964 25394 6020 25396
rect 5964 25342 5966 25394
rect 5966 25342 6018 25394
rect 6018 25342 6020 25394
rect 5964 25340 6020 25342
rect 5516 25228 5572 25284
rect 5404 25004 5460 25060
rect 5068 24892 5124 24948
rect 5068 23996 5124 24052
rect 4508 23938 4564 23940
rect 4508 23886 4510 23938
rect 4510 23886 4562 23938
rect 4562 23886 4564 23938
rect 4508 23884 4564 23886
rect 4284 23772 4340 23828
rect 4844 23714 4900 23716
rect 4844 23662 4846 23714
rect 4846 23662 4898 23714
rect 4898 23662 4900 23714
rect 4844 23660 4900 23662
rect 4732 23324 4788 23380
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 3836 22146 3892 22148
rect 3836 22094 3838 22146
rect 3838 22094 3890 22146
rect 3890 22094 3892 22146
rect 3836 22092 3892 22094
rect 3836 19906 3892 19908
rect 3836 19854 3838 19906
rect 3838 19854 3890 19906
rect 3890 19854 3892 19906
rect 3836 19852 3892 19854
rect 2940 19292 2996 19348
rect 2828 18060 2884 18116
rect 2604 16882 2660 16884
rect 2604 16830 2606 16882
rect 2606 16830 2658 16882
rect 2658 16830 2660 16882
rect 2604 16828 2660 16830
rect 2940 17836 2996 17892
rect 3052 19740 3108 19796
rect 4396 21644 4452 21700
rect 3948 19404 4004 19460
rect 4060 19292 4116 19348
rect 4620 21532 4676 21588
rect 4732 21644 4788 21700
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4284 18396 4340 18452
rect 3836 18284 3892 18340
rect 3500 18060 3556 18116
rect 5180 21644 5236 21700
rect 5292 21586 5348 21588
rect 5292 21534 5294 21586
rect 5294 21534 5346 21586
rect 5346 21534 5348 21586
rect 5292 21532 5348 21534
rect 5292 20188 5348 20244
rect 5292 19740 5348 19796
rect 5628 24946 5684 24948
rect 5628 24894 5630 24946
rect 5630 24894 5682 24946
rect 5682 24894 5684 24946
rect 5628 24892 5684 24894
rect 5516 23772 5572 23828
rect 5628 23324 5684 23380
rect 7196 26460 7252 26516
rect 7308 28700 7364 28756
rect 8204 31724 8260 31780
rect 9772 37436 9828 37492
rect 9772 35922 9828 35924
rect 9772 35870 9774 35922
rect 9774 35870 9826 35922
rect 9826 35870 9828 35922
rect 9772 35868 9828 35870
rect 10556 38668 10612 38724
rect 11788 40402 11844 40404
rect 11788 40350 11790 40402
rect 11790 40350 11842 40402
rect 11842 40350 11844 40402
rect 11788 40348 11844 40350
rect 11900 40236 11956 40292
rect 11004 39452 11060 39508
rect 10892 39228 10948 39284
rect 11116 39058 11172 39060
rect 11116 39006 11118 39058
rect 11118 39006 11170 39058
rect 11170 39006 11172 39058
rect 11116 39004 11172 39006
rect 11004 38946 11060 38948
rect 11004 38894 11006 38946
rect 11006 38894 11058 38946
rect 11058 38894 11060 38946
rect 11004 38892 11060 38894
rect 11228 38892 11284 38948
rect 10780 38556 10836 38612
rect 10444 37938 10500 37940
rect 10444 37886 10446 37938
rect 10446 37886 10498 37938
rect 10498 37886 10500 37938
rect 10444 37884 10500 37886
rect 10220 37436 10276 37492
rect 10444 37212 10500 37268
rect 10444 36988 10500 37044
rect 10332 36764 10388 36820
rect 9996 35810 10052 35812
rect 9996 35758 9998 35810
rect 9998 35758 10050 35810
rect 10050 35758 10052 35810
rect 9996 35756 10052 35758
rect 9884 35026 9940 35028
rect 9884 34974 9886 35026
rect 9886 34974 9938 35026
rect 9938 34974 9940 35026
rect 9884 34972 9940 34974
rect 8876 33516 8932 33572
rect 9100 34690 9156 34692
rect 9100 34638 9102 34690
rect 9102 34638 9154 34690
rect 9154 34638 9156 34690
rect 9100 34636 9156 34638
rect 8988 33292 9044 33348
rect 9436 34524 9492 34580
rect 8764 33068 8820 33124
rect 8764 31948 8820 32004
rect 8876 31612 8932 31668
rect 9996 34860 10052 34916
rect 10668 37378 10724 37380
rect 10668 37326 10670 37378
rect 10670 37326 10722 37378
rect 10722 37326 10724 37378
rect 10668 37324 10724 37326
rect 11788 39340 11844 39396
rect 11452 38780 11508 38836
rect 11564 39004 11620 39060
rect 11564 38668 11620 38724
rect 11004 37826 11060 37828
rect 11004 37774 11006 37826
rect 11006 37774 11058 37826
rect 11058 37774 11060 37826
rect 11004 37772 11060 37774
rect 10668 35868 10724 35924
rect 10444 35308 10500 35364
rect 9772 34748 9828 34804
rect 10332 34802 10388 34804
rect 10332 34750 10334 34802
rect 10334 34750 10386 34802
rect 10386 34750 10388 34802
rect 10332 34748 10388 34750
rect 9772 33964 9828 34020
rect 10332 34130 10388 34132
rect 10332 34078 10334 34130
rect 10334 34078 10386 34130
rect 10386 34078 10388 34130
rect 10332 34076 10388 34078
rect 10108 34018 10164 34020
rect 10108 33966 10110 34018
rect 10110 33966 10162 34018
rect 10162 33966 10164 34018
rect 10108 33964 10164 33966
rect 9996 33404 10052 33460
rect 10332 33740 10388 33796
rect 9772 32060 9828 32116
rect 9436 31948 9492 32004
rect 8988 31836 9044 31892
rect 9436 31778 9492 31780
rect 9436 31726 9438 31778
rect 9438 31726 9490 31778
rect 9490 31726 9492 31778
rect 9436 31724 9492 31726
rect 8988 31052 9044 31108
rect 8204 30940 8260 30996
rect 8428 30770 8484 30772
rect 8428 30718 8430 30770
rect 8430 30718 8482 30770
rect 8482 30718 8484 30770
rect 8428 30716 8484 30718
rect 9660 31052 9716 31108
rect 9436 30716 9492 30772
rect 9212 30210 9268 30212
rect 9212 30158 9214 30210
rect 9214 30158 9266 30210
rect 9266 30158 9268 30210
rect 9212 30156 9268 30158
rect 8428 29538 8484 29540
rect 8428 29486 8430 29538
rect 8430 29486 8482 29538
rect 8482 29486 8484 29538
rect 8428 29484 8484 29486
rect 8540 29260 8596 29316
rect 8540 28812 8596 28868
rect 8092 28700 8148 28756
rect 7980 28140 8036 28196
rect 8316 28028 8372 28084
rect 7644 27916 7700 27972
rect 7532 27858 7588 27860
rect 7532 27806 7534 27858
rect 7534 27806 7586 27858
rect 7586 27806 7588 27858
rect 7532 27804 7588 27806
rect 7420 27746 7476 27748
rect 7420 27694 7422 27746
rect 7422 27694 7474 27746
rect 7474 27694 7476 27746
rect 7420 27692 7476 27694
rect 7532 27580 7588 27636
rect 7308 26348 7364 26404
rect 8428 27020 8484 27076
rect 8540 28364 8596 28420
rect 8652 27970 8708 27972
rect 8652 27918 8654 27970
rect 8654 27918 8706 27970
rect 8706 27918 8708 27970
rect 8652 27916 8708 27918
rect 6412 24892 6468 24948
rect 7084 26012 7140 26068
rect 6748 25452 6804 25508
rect 6188 24780 6244 24836
rect 7420 25228 7476 25284
rect 6972 24834 7028 24836
rect 6972 24782 6974 24834
rect 6974 24782 7026 24834
rect 7026 24782 7028 24834
rect 6972 24780 7028 24782
rect 6076 23884 6132 23940
rect 6412 23436 6468 23492
rect 6188 23154 6244 23156
rect 6188 23102 6190 23154
rect 6190 23102 6242 23154
rect 6242 23102 6244 23154
rect 6188 23100 6244 23102
rect 5852 21644 5908 21700
rect 5740 21308 5796 21364
rect 5740 20860 5796 20916
rect 5628 19346 5684 19348
rect 5628 19294 5630 19346
rect 5630 19294 5682 19346
rect 5682 19294 5684 19346
rect 5628 19292 5684 19294
rect 5516 18396 5572 18452
rect 4956 18060 5012 18116
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4396 17836 4452 17892
rect 3948 17612 4004 17668
rect 3276 17442 3332 17444
rect 3276 17390 3278 17442
rect 3278 17390 3330 17442
rect 3330 17390 3332 17442
rect 3276 17388 3332 17390
rect 3164 16994 3220 16996
rect 3164 16942 3166 16994
rect 3166 16942 3218 16994
rect 3218 16942 3220 16994
rect 3164 16940 3220 16942
rect 3164 16716 3220 16772
rect 3724 17164 3780 17220
rect 4844 17836 4900 17892
rect 4844 17612 4900 17668
rect 5180 17948 5236 18004
rect 5740 18172 5796 18228
rect 6748 20972 6804 21028
rect 6972 22428 7028 22484
rect 6300 20802 6356 20804
rect 6300 20750 6302 20802
rect 6302 20750 6354 20802
rect 6354 20750 6356 20802
rect 6300 20748 6356 20750
rect 6076 20636 6132 20692
rect 6524 20524 6580 20580
rect 6188 19404 6244 19460
rect 6076 19122 6132 19124
rect 6076 19070 6078 19122
rect 6078 19070 6130 19122
rect 6130 19070 6132 19122
rect 6076 19068 6132 19070
rect 6188 18956 6244 19012
rect 5964 18844 6020 18900
rect 5852 17948 5908 18004
rect 6412 18620 6468 18676
rect 7420 21756 7476 21812
rect 7420 20188 7476 20244
rect 7756 26908 7812 26964
rect 8876 29820 8932 29876
rect 8988 29372 9044 29428
rect 9548 30380 9604 30436
rect 9660 30210 9716 30212
rect 9660 30158 9662 30210
rect 9662 30158 9714 30210
rect 9714 30158 9716 30210
rect 9660 30156 9716 30158
rect 9884 31500 9940 31556
rect 9772 29820 9828 29876
rect 9884 29538 9940 29540
rect 9884 29486 9886 29538
rect 9886 29486 9938 29538
rect 9938 29486 9940 29538
rect 9884 29484 9940 29486
rect 9548 29426 9604 29428
rect 9548 29374 9550 29426
rect 9550 29374 9602 29426
rect 9602 29374 9604 29426
rect 9548 29372 9604 29374
rect 8988 28588 9044 28644
rect 9212 28700 9268 28756
rect 10332 31276 10388 31332
rect 10220 31164 10276 31220
rect 10332 30380 10388 30436
rect 10220 29708 10276 29764
rect 9884 28476 9940 28532
rect 9212 28140 9268 28196
rect 8204 26012 8260 26068
rect 8204 24722 8260 24724
rect 8204 24670 8206 24722
rect 8206 24670 8258 24722
rect 8258 24670 8260 24722
rect 8204 24668 8260 24670
rect 7756 20972 7812 21028
rect 7756 20636 7812 20692
rect 8316 23996 8372 24052
rect 8204 22876 8260 22932
rect 8540 25506 8596 25508
rect 8540 25454 8542 25506
rect 8542 25454 8594 25506
rect 8594 25454 8596 25506
rect 8540 25452 8596 25454
rect 8204 21644 8260 21700
rect 8092 20524 8148 20580
rect 8540 20972 8596 21028
rect 7980 20412 8036 20468
rect 7644 19404 7700 19460
rect 6300 18396 6356 18452
rect 6524 18060 6580 18116
rect 5516 17612 5572 17668
rect 5404 17500 5460 17556
rect 3612 16940 3668 16996
rect 3276 16156 3332 16212
rect 3500 16828 3556 16884
rect 2716 15874 2772 15876
rect 2716 15822 2718 15874
rect 2718 15822 2770 15874
rect 2770 15822 2772 15874
rect 2716 15820 2772 15822
rect 2268 13970 2324 13972
rect 2268 13918 2270 13970
rect 2270 13918 2322 13970
rect 2322 13918 2324 13970
rect 2268 13916 2324 13918
rect 2828 15036 2884 15092
rect 2716 14364 2772 14420
rect 3164 13692 3220 13748
rect 3276 13132 3332 13188
rect 1932 12460 1988 12516
rect 2268 11788 2324 11844
rect 2156 10498 2212 10500
rect 2156 10446 2158 10498
rect 2158 10446 2210 10498
rect 2210 10446 2212 10498
rect 2156 10444 2212 10446
rect 2044 9714 2100 9716
rect 2044 9662 2046 9714
rect 2046 9662 2098 9714
rect 2098 9662 2100 9714
rect 2044 9660 2100 9662
rect 2044 9042 2100 9044
rect 2044 8990 2046 9042
rect 2046 8990 2098 9042
rect 2098 8990 2100 9042
rect 2044 8988 2100 8990
rect 3836 16828 3892 16884
rect 4956 16828 5012 16884
rect 4060 16658 4116 16660
rect 4060 16606 4062 16658
rect 4062 16606 4114 16658
rect 4114 16606 4116 16658
rect 4060 16604 4116 16606
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4956 16492 5012 16548
rect 3948 15932 4004 15988
rect 4060 16268 4116 16324
rect 3500 15596 3556 15652
rect 3948 15484 4004 15540
rect 4396 16044 4452 16100
rect 4284 15986 4340 15988
rect 4284 15934 4286 15986
rect 4286 15934 4338 15986
rect 4338 15934 4340 15986
rect 4284 15932 4340 15934
rect 4844 15986 4900 15988
rect 4844 15934 4846 15986
rect 4846 15934 4898 15986
rect 4898 15934 4900 15986
rect 4844 15932 4900 15934
rect 4956 15874 5012 15876
rect 4956 15822 4958 15874
rect 4958 15822 5010 15874
rect 5010 15822 5012 15874
rect 4956 15820 5012 15822
rect 6300 17554 6356 17556
rect 6300 17502 6302 17554
rect 6302 17502 6354 17554
rect 6354 17502 6356 17554
rect 6300 17500 6356 17502
rect 5740 16828 5796 16884
rect 5628 15932 5684 15988
rect 4620 15484 4676 15540
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4172 14700 4228 14756
rect 4844 14588 4900 14644
rect 3500 13020 3556 13076
rect 3612 13580 3668 13636
rect 3052 12178 3108 12180
rect 3052 12126 3054 12178
rect 3054 12126 3106 12178
rect 3106 12126 3108 12178
rect 3052 12124 3108 12126
rect 2828 12066 2884 12068
rect 2828 12014 2830 12066
rect 2830 12014 2882 12066
rect 2882 12014 2884 12066
rect 2828 12012 2884 12014
rect 3052 11788 3108 11844
rect 2940 10780 2996 10836
rect 3052 10892 3108 10948
rect 2940 9266 2996 9268
rect 2940 9214 2942 9266
rect 2942 9214 2994 9266
rect 2994 9214 2996 9266
rect 2940 9212 2996 9214
rect 3500 11452 3556 11508
rect 4172 14252 4228 14308
rect 4060 13020 4116 13076
rect 3836 12290 3892 12292
rect 3836 12238 3838 12290
rect 3838 12238 3890 12290
rect 3890 12238 3892 12290
rect 3836 12236 3892 12238
rect 3948 12124 4004 12180
rect 4172 12738 4228 12740
rect 4172 12686 4174 12738
rect 4174 12686 4226 12738
rect 4226 12686 4228 12738
rect 4172 12684 4228 12686
rect 3388 9602 3444 9604
rect 3388 9550 3390 9602
rect 3390 9550 3442 9602
rect 3442 9550 3444 9602
rect 3388 9548 3444 9550
rect 3388 9324 3444 9380
rect 3836 9826 3892 9828
rect 3836 9774 3838 9826
rect 3838 9774 3890 9826
rect 3890 9774 3892 9826
rect 3836 9772 3892 9774
rect 4844 14418 4900 14420
rect 4844 14366 4846 14418
rect 4846 14366 4898 14418
rect 4898 14366 4900 14418
rect 4844 14364 4900 14366
rect 4620 13468 4676 13524
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 5292 15484 5348 15540
rect 5516 15426 5572 15428
rect 5516 15374 5518 15426
rect 5518 15374 5570 15426
rect 5570 15374 5572 15426
rect 5516 15372 5572 15374
rect 7084 18674 7140 18676
rect 7084 18622 7086 18674
rect 7086 18622 7138 18674
rect 7138 18622 7140 18674
rect 7084 18620 7140 18622
rect 6972 18396 7028 18452
rect 7196 18338 7252 18340
rect 7196 18286 7198 18338
rect 7198 18286 7250 18338
rect 7250 18286 7252 18338
rect 7196 18284 7252 18286
rect 6636 16882 6692 16884
rect 6636 16830 6638 16882
rect 6638 16830 6690 16882
rect 6690 16830 6692 16882
rect 6636 16828 6692 16830
rect 6076 16210 6132 16212
rect 6076 16158 6078 16210
rect 6078 16158 6130 16210
rect 6130 16158 6132 16210
rect 6076 16156 6132 16158
rect 6300 15986 6356 15988
rect 6300 15934 6302 15986
rect 6302 15934 6354 15986
rect 6354 15934 6356 15986
rect 6300 15932 6356 15934
rect 5068 14476 5124 14532
rect 5404 14924 5460 14980
rect 5292 14812 5348 14868
rect 5068 13692 5124 13748
rect 5292 13468 5348 13524
rect 5516 14700 5572 14756
rect 5404 14364 5460 14420
rect 4844 12572 4900 12628
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 5068 11564 5124 11620
rect 4508 11116 4564 11172
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 5292 10220 5348 10276
rect 4684 10164 4740 10166
rect 4060 9212 4116 9268
rect 4172 9324 4228 9380
rect 3276 8818 3332 8820
rect 3276 8766 3278 8818
rect 3278 8766 3330 8818
rect 3330 8766 3332 8818
rect 3276 8764 3332 8766
rect 2828 8034 2884 8036
rect 2828 7982 2830 8034
rect 2830 7982 2882 8034
rect 2882 7982 2884 8034
rect 2828 7980 2884 7982
rect 3164 7362 3220 7364
rect 3164 7310 3166 7362
rect 3166 7310 3218 7362
rect 3218 7310 3220 7362
rect 3164 7308 3220 7310
rect 2716 6860 2772 6916
rect 4060 8316 4116 8372
rect 3724 8258 3780 8260
rect 3724 8206 3726 8258
rect 3726 8206 3778 8258
rect 3778 8206 3780 8258
rect 3724 8204 3780 8206
rect 3388 6578 3444 6580
rect 3388 6526 3390 6578
rect 3390 6526 3442 6578
rect 3442 6526 3444 6578
rect 3388 6524 3444 6526
rect 3836 6690 3892 6692
rect 3836 6638 3838 6690
rect 3838 6638 3890 6690
rect 3890 6638 3892 6690
rect 3836 6636 3892 6638
rect 3836 5180 3892 5236
rect 5068 9436 5124 9492
rect 4284 9100 4340 9156
rect 5516 13468 5572 13524
rect 5740 14306 5796 14308
rect 5740 14254 5742 14306
rect 5742 14254 5794 14306
rect 5794 14254 5796 14306
rect 5740 14252 5796 14254
rect 6188 15874 6244 15876
rect 6188 15822 6190 15874
rect 6190 15822 6242 15874
rect 6242 15822 6244 15874
rect 6188 15820 6244 15822
rect 6412 15314 6468 15316
rect 6412 15262 6414 15314
rect 6414 15262 6466 15314
rect 6466 15262 6468 15314
rect 6412 15260 6468 15262
rect 6300 15148 6356 15204
rect 6300 14924 6356 14980
rect 6636 16044 6692 16100
rect 7196 17388 7252 17444
rect 7308 17276 7364 17332
rect 8092 19906 8148 19908
rect 8092 19854 8094 19906
rect 8094 19854 8146 19906
rect 8146 19854 8148 19906
rect 8092 19852 8148 19854
rect 7868 19516 7924 19572
rect 7756 19122 7812 19124
rect 7756 19070 7758 19122
rect 7758 19070 7810 19122
rect 7810 19070 7812 19122
rect 7756 19068 7812 19070
rect 7644 18396 7700 18452
rect 7532 17948 7588 18004
rect 7420 17164 7476 17220
rect 7196 16940 7252 16996
rect 6748 15932 6804 15988
rect 7196 16156 7252 16212
rect 6860 15820 6916 15876
rect 7308 16098 7364 16100
rect 7308 16046 7310 16098
rect 7310 16046 7362 16098
rect 7362 16046 7364 16098
rect 7308 16044 7364 16046
rect 7196 15202 7252 15204
rect 7196 15150 7198 15202
rect 7198 15150 7250 15202
rect 7250 15150 7252 15202
rect 7196 15148 7252 15150
rect 7420 15372 7476 15428
rect 6524 14812 6580 14868
rect 5964 14700 6020 14756
rect 6076 14588 6132 14644
rect 5964 14418 6020 14420
rect 5964 14366 5966 14418
rect 5966 14366 6018 14418
rect 6018 14366 6020 14418
rect 5964 14364 6020 14366
rect 6412 14364 6468 14420
rect 6636 14418 6692 14420
rect 6636 14366 6638 14418
rect 6638 14366 6690 14418
rect 6690 14366 6692 14418
rect 6636 14364 6692 14366
rect 6076 14252 6132 14308
rect 6524 14306 6580 14308
rect 6524 14254 6526 14306
rect 6526 14254 6578 14306
rect 6578 14254 6580 14306
rect 6524 14252 6580 14254
rect 6300 13468 6356 13524
rect 5852 13132 5908 13188
rect 6412 13244 6468 13300
rect 5628 10668 5684 10724
rect 5740 12460 5796 12516
rect 5516 9436 5572 9492
rect 6188 12236 6244 12292
rect 6412 12124 6468 12180
rect 5964 11900 6020 11956
rect 5852 11170 5908 11172
rect 5852 11118 5854 11170
rect 5854 11118 5906 11170
rect 5906 11118 5908 11170
rect 5852 11116 5908 11118
rect 6300 11394 6356 11396
rect 6300 11342 6302 11394
rect 6302 11342 6354 11394
rect 6354 11342 6356 11394
rect 6300 11340 6356 11342
rect 5964 9660 6020 9716
rect 6076 11004 6132 11060
rect 5740 9324 5796 9380
rect 5404 8988 5460 9044
rect 5516 9212 5572 9268
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4956 8876 5012 8932
rect 4620 7868 4676 7924
rect 4172 7586 4228 7588
rect 4172 7534 4174 7586
rect 4174 7534 4226 7586
rect 4226 7534 4228 7586
rect 4172 7532 4228 7534
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4284 6578 4340 6580
rect 4284 6526 4286 6578
rect 4286 6526 4338 6578
rect 4338 6526 4340 6578
rect 4284 6524 4340 6526
rect 5740 8146 5796 8148
rect 5740 8094 5742 8146
rect 5742 8094 5794 8146
rect 5794 8094 5796 8146
rect 5740 8092 5796 8094
rect 5628 7532 5684 7588
rect 5516 6524 5572 6580
rect 5852 6524 5908 6580
rect 5964 6972 6020 7028
rect 5180 6188 5236 6244
rect 4620 5794 4676 5796
rect 4620 5742 4622 5794
rect 4622 5742 4674 5794
rect 4674 5742 4676 5794
rect 4620 5740 4676 5742
rect 5628 5740 5684 5796
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 5740 5292 5796 5348
rect 4620 5234 4676 5236
rect 4620 5182 4622 5234
rect 4622 5182 4674 5234
rect 4674 5182 4676 5234
rect 4620 5180 4676 5182
rect 5068 5234 5124 5236
rect 5068 5182 5070 5234
rect 5070 5182 5122 5234
rect 5122 5182 5124 5234
rect 5068 5180 5124 5182
rect 6188 10444 6244 10500
rect 6972 13468 7028 13524
rect 7084 13020 7140 13076
rect 7084 12460 7140 12516
rect 6748 12402 6804 12404
rect 6748 12350 6750 12402
rect 6750 12350 6802 12402
rect 6802 12350 6804 12402
rect 6748 12348 6804 12350
rect 6860 11676 6916 11732
rect 6972 11564 7028 11620
rect 6748 11394 6804 11396
rect 6748 11342 6750 11394
rect 6750 11342 6802 11394
rect 6802 11342 6804 11394
rect 6748 11340 6804 11342
rect 7756 17554 7812 17556
rect 7756 17502 7758 17554
rect 7758 17502 7810 17554
rect 7810 17502 7812 17554
rect 7756 17500 7812 17502
rect 7644 17442 7700 17444
rect 7644 17390 7646 17442
rect 7646 17390 7698 17442
rect 7698 17390 7700 17442
rect 7644 17388 7700 17390
rect 7868 17388 7924 17444
rect 8428 19234 8484 19236
rect 8428 19182 8430 19234
rect 8430 19182 8482 19234
rect 8482 19182 8484 19234
rect 8428 19180 8484 19182
rect 8092 17948 8148 18004
rect 7644 15932 7700 15988
rect 7868 15708 7924 15764
rect 7868 15260 7924 15316
rect 7532 14028 7588 14084
rect 7980 15148 8036 15204
rect 7756 14530 7812 14532
rect 7756 14478 7758 14530
rect 7758 14478 7810 14530
rect 7810 14478 7812 14530
rect 7756 14476 7812 14478
rect 7980 14306 8036 14308
rect 7980 14254 7982 14306
rect 7982 14254 8034 14306
rect 8034 14254 8036 14306
rect 7980 14252 8036 14254
rect 7868 14140 7924 14196
rect 7532 12796 7588 12852
rect 7644 13468 7700 13524
rect 7980 13916 8036 13972
rect 7420 12348 7476 12404
rect 7644 12572 7700 12628
rect 7308 12236 7364 12292
rect 7980 13468 8036 13524
rect 7868 12124 7924 12180
rect 7980 12684 8036 12740
rect 7196 11900 7252 11956
rect 7532 11900 7588 11956
rect 7196 11676 7252 11732
rect 6972 11116 7028 11172
rect 7196 10834 7252 10836
rect 7196 10782 7198 10834
rect 7198 10782 7250 10834
rect 7250 10782 7252 10834
rect 7196 10780 7252 10782
rect 6972 10722 7028 10724
rect 6972 10670 6974 10722
rect 6974 10670 7026 10722
rect 7026 10670 7028 10722
rect 6972 10668 7028 10670
rect 6412 9212 6468 9268
rect 6636 10220 6692 10276
rect 6524 8988 6580 9044
rect 6300 8204 6356 8260
rect 6972 10108 7028 10164
rect 7868 11676 7924 11732
rect 7308 10108 7364 10164
rect 6972 9212 7028 9268
rect 7644 9884 7700 9940
rect 7868 9660 7924 9716
rect 7196 8988 7252 9044
rect 7532 9436 7588 9492
rect 6860 8428 6916 8484
rect 9100 19122 9156 19124
rect 9100 19070 9102 19122
rect 9102 19070 9154 19122
rect 9154 19070 9156 19122
rect 9100 19068 9156 19070
rect 8428 18226 8484 18228
rect 8428 18174 8430 18226
rect 8430 18174 8482 18226
rect 8482 18174 8484 18226
rect 8428 18172 8484 18174
rect 8204 17666 8260 17668
rect 8204 17614 8206 17666
rect 8206 17614 8258 17666
rect 8258 17614 8260 17666
rect 8204 17612 8260 17614
rect 8428 16828 8484 16884
rect 8988 17554 9044 17556
rect 8988 17502 8990 17554
rect 8990 17502 9042 17554
rect 9042 17502 9044 17554
rect 8988 17500 9044 17502
rect 10108 28140 10164 28196
rect 10556 33292 10612 33348
rect 10892 35868 10948 35924
rect 11004 35084 11060 35140
rect 12460 40460 12516 40516
rect 14028 40572 14084 40628
rect 13468 40514 13524 40516
rect 13468 40462 13470 40514
rect 13470 40462 13522 40514
rect 13522 40462 13524 40514
rect 13468 40460 13524 40462
rect 13132 40402 13188 40404
rect 13132 40350 13134 40402
rect 13134 40350 13186 40402
rect 13186 40350 13188 40402
rect 13132 40348 13188 40350
rect 13580 40290 13636 40292
rect 13580 40238 13582 40290
rect 13582 40238 13634 40290
rect 13634 40238 13636 40290
rect 13580 40236 13636 40238
rect 11564 37826 11620 37828
rect 11564 37774 11566 37826
rect 11566 37774 11618 37826
rect 11618 37774 11620 37826
rect 11564 37772 11620 37774
rect 11340 37212 11396 37268
rect 11900 37324 11956 37380
rect 12124 37826 12180 37828
rect 12124 37774 12126 37826
rect 12126 37774 12178 37826
rect 12178 37774 12180 37826
rect 12124 37772 12180 37774
rect 13020 39618 13076 39620
rect 13020 39566 13022 39618
rect 13022 39566 13074 39618
rect 13074 39566 13076 39618
rect 13020 39564 13076 39566
rect 13804 39618 13860 39620
rect 13804 39566 13806 39618
rect 13806 39566 13858 39618
rect 13858 39566 13860 39618
rect 13804 39564 13860 39566
rect 12124 37212 12180 37268
rect 12012 36428 12068 36484
rect 12460 37212 12516 37268
rect 11788 35532 11844 35588
rect 11900 35644 11956 35700
rect 11116 34972 11172 35028
rect 11116 34636 11172 34692
rect 11004 34018 11060 34020
rect 11004 33966 11006 34018
rect 11006 33966 11058 34018
rect 11058 33966 11060 34018
rect 11004 33964 11060 33966
rect 10892 33740 10948 33796
rect 10892 32396 10948 32452
rect 11004 32620 11060 32676
rect 10892 32060 10948 32116
rect 10556 30156 10612 30212
rect 10556 29596 10612 29652
rect 10332 29036 10388 29092
rect 10444 29484 10500 29540
rect 9660 27804 9716 27860
rect 10108 27916 10164 27972
rect 9660 27468 9716 27524
rect 10332 27020 10388 27076
rect 9548 25340 9604 25396
rect 10220 25340 10276 25396
rect 9548 24892 9604 24948
rect 9660 23938 9716 23940
rect 9660 23886 9662 23938
rect 9662 23886 9714 23938
rect 9714 23886 9716 23938
rect 9660 23884 9716 23886
rect 9660 23212 9716 23268
rect 10108 23212 10164 23268
rect 10220 23324 10276 23380
rect 9772 20860 9828 20916
rect 9884 20412 9940 20468
rect 9996 20188 10052 20244
rect 9884 20018 9940 20020
rect 9884 19966 9886 20018
rect 9886 19966 9938 20018
rect 9938 19966 9940 20018
rect 9884 19964 9940 19966
rect 9660 18172 9716 18228
rect 8652 16604 8708 16660
rect 8316 15426 8372 15428
rect 8316 15374 8318 15426
rect 8318 15374 8370 15426
rect 8370 15374 8372 15426
rect 8316 15372 8372 15374
rect 8204 14364 8260 14420
rect 8316 14700 8372 14756
rect 8092 12348 8148 12404
rect 8204 13020 8260 13076
rect 8092 11394 8148 11396
rect 8092 11342 8094 11394
rect 8094 11342 8146 11394
rect 8146 11342 8148 11394
rect 8092 11340 8148 11342
rect 8764 15314 8820 15316
rect 8764 15262 8766 15314
rect 8766 15262 8818 15314
rect 8818 15262 8820 15314
rect 8764 15260 8820 15262
rect 8988 15148 9044 15204
rect 8652 13916 8708 13972
rect 8428 13746 8484 13748
rect 8428 13694 8430 13746
rect 8430 13694 8482 13746
rect 8482 13694 8484 13746
rect 8428 13692 8484 13694
rect 8540 13468 8596 13524
rect 8652 13132 8708 13188
rect 8316 12684 8372 12740
rect 9436 14642 9492 14644
rect 9436 14590 9438 14642
rect 9438 14590 9490 14642
rect 9490 14590 9492 14642
rect 9436 14588 9492 14590
rect 9212 14530 9268 14532
rect 9212 14478 9214 14530
rect 9214 14478 9266 14530
rect 9266 14478 9268 14530
rect 9212 14476 9268 14478
rect 10220 21868 10276 21924
rect 10556 28700 10612 28756
rect 10668 29148 10724 29204
rect 10668 28364 10724 28420
rect 10780 27916 10836 27972
rect 11900 35084 11956 35140
rect 12460 36482 12516 36484
rect 12460 36430 12462 36482
rect 12462 36430 12514 36482
rect 12514 36430 12516 36482
rect 12460 36428 12516 36430
rect 13020 38834 13076 38836
rect 13020 38782 13022 38834
rect 13022 38782 13074 38834
rect 13074 38782 13076 38834
rect 13020 38780 13076 38782
rect 12908 37996 12964 38052
rect 12908 37548 12964 37604
rect 13020 37324 13076 37380
rect 12684 35922 12740 35924
rect 12684 35870 12686 35922
rect 12686 35870 12738 35922
rect 12738 35870 12740 35922
rect 12684 35868 12740 35870
rect 12572 35698 12628 35700
rect 12572 35646 12574 35698
rect 12574 35646 12626 35698
rect 12626 35646 12628 35698
rect 12572 35644 12628 35646
rect 12012 34748 12068 34804
rect 12572 34860 12628 34916
rect 11676 34636 11732 34692
rect 11676 34242 11732 34244
rect 11676 34190 11678 34242
rect 11678 34190 11730 34242
rect 11730 34190 11732 34242
rect 11676 34188 11732 34190
rect 11676 33346 11732 33348
rect 11676 33294 11678 33346
rect 11678 33294 11730 33346
rect 11730 33294 11732 33346
rect 11676 33292 11732 33294
rect 12012 33346 12068 33348
rect 12012 33294 12014 33346
rect 12014 33294 12066 33346
rect 12066 33294 12068 33346
rect 12012 33292 12068 33294
rect 11452 33122 11508 33124
rect 11452 33070 11454 33122
rect 11454 33070 11506 33122
rect 11506 33070 11508 33122
rect 11452 33068 11508 33070
rect 11228 32732 11284 32788
rect 11340 31836 11396 31892
rect 11340 31276 11396 31332
rect 11900 32786 11956 32788
rect 11900 32734 11902 32786
rect 11902 32734 11954 32786
rect 11954 32734 11956 32786
rect 11900 32732 11956 32734
rect 11788 32002 11844 32004
rect 11788 31950 11790 32002
rect 11790 31950 11842 32002
rect 11842 31950 11844 32002
rect 11788 31948 11844 31950
rect 11564 31500 11620 31556
rect 11564 30716 11620 30772
rect 11004 30044 11060 30100
rect 11004 29036 11060 29092
rect 11900 29820 11956 29876
rect 11228 28812 11284 28868
rect 11340 29708 11396 29764
rect 11116 28476 11172 28532
rect 11788 29650 11844 29652
rect 11788 29598 11790 29650
rect 11790 29598 11842 29650
rect 11842 29598 11844 29650
rect 11788 29596 11844 29598
rect 12348 34354 12404 34356
rect 12348 34302 12350 34354
rect 12350 34302 12402 34354
rect 12402 34302 12404 34354
rect 12348 34300 12404 34302
rect 12796 35420 12852 35476
rect 12236 33628 12292 33684
rect 12684 32508 12740 32564
rect 12572 32450 12628 32452
rect 12572 32398 12574 32450
rect 12574 32398 12626 32450
rect 12626 32398 12628 32450
rect 12572 32396 12628 32398
rect 12460 31778 12516 31780
rect 12460 31726 12462 31778
rect 12462 31726 12514 31778
rect 12514 31726 12516 31778
rect 12460 31724 12516 31726
rect 12124 31052 12180 31108
rect 12236 30604 12292 30660
rect 11676 28812 11732 28868
rect 11340 28140 11396 28196
rect 11228 28082 11284 28084
rect 11228 28030 11230 28082
rect 11230 28030 11282 28082
rect 11282 28030 11284 28082
rect 11228 28028 11284 28030
rect 11788 27916 11844 27972
rect 10556 25900 10612 25956
rect 10668 26012 10724 26068
rect 10556 24220 10612 24276
rect 10780 25676 10836 25732
rect 11340 27468 11396 27524
rect 11564 26290 11620 26292
rect 11564 26238 11566 26290
rect 11566 26238 11618 26290
rect 11618 26238 11620 26290
rect 11564 26236 11620 26238
rect 10892 24108 10948 24164
rect 10780 23436 10836 23492
rect 10444 21868 10500 21924
rect 10220 20524 10276 20580
rect 10780 21810 10836 21812
rect 10780 21758 10782 21810
rect 10782 21758 10834 21810
rect 10834 21758 10836 21810
rect 10780 21756 10836 21758
rect 10892 22652 10948 22708
rect 10668 21532 10724 21588
rect 10556 20524 10612 20580
rect 10220 18396 10276 18452
rect 10668 19180 10724 19236
rect 10780 21196 10836 21252
rect 10108 17500 10164 17556
rect 10108 17276 10164 17332
rect 9884 15596 9940 15652
rect 9100 14364 9156 14420
rect 9100 13916 9156 13972
rect 8092 9884 8148 9940
rect 8316 9436 8372 9492
rect 7980 9042 8036 9044
rect 7980 8990 7982 9042
rect 7982 8990 8034 9042
rect 8034 8990 8036 9042
rect 7980 8988 8036 8990
rect 7420 8764 7476 8820
rect 6524 7756 6580 7812
rect 6860 7644 6916 7700
rect 6972 8034 7028 8036
rect 6972 7982 6974 8034
rect 6974 7982 7026 8034
rect 7026 7982 7028 8034
rect 6972 7980 7028 7982
rect 7532 7980 7588 8036
rect 7868 8930 7924 8932
rect 7868 8878 7870 8930
rect 7870 8878 7922 8930
rect 7922 8878 7924 8930
rect 7868 8876 7924 8878
rect 7980 8652 8036 8708
rect 7868 7980 7924 8036
rect 7644 7868 7700 7924
rect 6972 7474 7028 7476
rect 6972 7422 6974 7474
rect 6974 7422 7026 7474
rect 7026 7422 7028 7474
rect 6972 7420 7028 7422
rect 6748 6748 6804 6804
rect 6076 6412 6132 6468
rect 6188 6076 6244 6132
rect 6412 6466 6468 6468
rect 6412 6414 6414 6466
rect 6414 6414 6466 6466
rect 6466 6414 6468 6466
rect 6412 6412 6468 6414
rect 6300 5740 6356 5796
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 6188 5180 6244 5236
rect 7532 7474 7588 7476
rect 7532 7422 7534 7474
rect 7534 7422 7586 7474
rect 7586 7422 7588 7474
rect 7532 7420 7588 7422
rect 7420 6690 7476 6692
rect 7420 6638 7422 6690
rect 7422 6638 7474 6690
rect 7474 6638 7476 6690
rect 7420 6636 7476 6638
rect 7084 6466 7140 6468
rect 7084 6414 7086 6466
rect 7086 6414 7138 6466
rect 7138 6414 7140 6466
rect 7084 6412 7140 6414
rect 7420 6412 7476 6468
rect 7084 6130 7140 6132
rect 7084 6078 7086 6130
rect 7086 6078 7138 6130
rect 7138 6078 7140 6130
rect 7084 6076 7140 6078
rect 7308 5740 7364 5796
rect 8204 8258 8260 8260
rect 8204 8206 8206 8258
rect 8206 8206 8258 8258
rect 8258 8206 8260 8258
rect 8204 8204 8260 8206
rect 8092 8146 8148 8148
rect 8092 8094 8094 8146
rect 8094 8094 8146 8146
rect 8146 8094 8148 8146
rect 8092 8092 8148 8094
rect 8652 12290 8708 12292
rect 8652 12238 8654 12290
rect 8654 12238 8706 12290
rect 8706 12238 8708 12290
rect 8652 12236 8708 12238
rect 10780 18508 10836 18564
rect 10332 16604 10388 16660
rect 10332 16044 10388 16100
rect 10444 15986 10500 15988
rect 10444 15934 10446 15986
rect 10446 15934 10498 15986
rect 10498 15934 10500 15986
rect 10444 15932 10500 15934
rect 9884 15036 9940 15092
rect 9996 14700 10052 14756
rect 10220 14924 10276 14980
rect 9772 14364 9828 14420
rect 9100 13468 9156 13524
rect 9100 12908 9156 12964
rect 9660 12908 9716 12964
rect 9548 12460 9604 12516
rect 9100 12124 9156 12180
rect 8988 12012 9044 12068
rect 9660 11788 9716 11844
rect 9884 13132 9940 13188
rect 9996 12908 10052 12964
rect 10220 13804 10276 13860
rect 10444 14700 10500 14756
rect 11340 26124 11396 26180
rect 11116 22316 11172 22372
rect 11116 21698 11172 21700
rect 11116 21646 11118 21698
rect 11118 21646 11170 21698
rect 11170 21646 11172 21698
rect 11116 21644 11172 21646
rect 11116 21420 11172 21476
rect 11788 24892 11844 24948
rect 12460 30156 12516 30212
rect 12348 29708 12404 29764
rect 12908 30380 12964 30436
rect 13132 36764 13188 36820
rect 13580 38892 13636 38948
rect 16940 42530 16996 42532
rect 16940 42478 16942 42530
rect 16942 42478 16994 42530
rect 16994 42478 16996 42530
rect 16940 42476 16996 42478
rect 16828 41970 16884 41972
rect 16828 41918 16830 41970
rect 16830 41918 16882 41970
rect 16882 41918 16884 41970
rect 16828 41916 16884 41918
rect 14476 40290 14532 40292
rect 14476 40238 14478 40290
rect 14478 40238 14530 40290
rect 14530 40238 14532 40290
rect 14476 40236 14532 40238
rect 14924 39228 14980 39284
rect 13916 39116 13972 39172
rect 14028 38780 14084 38836
rect 13580 38050 13636 38052
rect 13580 37998 13582 38050
rect 13582 37998 13634 38050
rect 13634 37998 13636 38050
rect 13580 37996 13636 37998
rect 14140 37212 14196 37268
rect 14588 37996 14644 38052
rect 14364 36652 14420 36708
rect 14700 36706 14756 36708
rect 14700 36654 14702 36706
rect 14702 36654 14754 36706
rect 14754 36654 14756 36706
rect 14700 36652 14756 36654
rect 13132 35868 13188 35924
rect 13244 36092 13300 36148
rect 13468 35532 13524 35588
rect 13244 35084 13300 35140
rect 13244 31836 13300 31892
rect 13132 31612 13188 31668
rect 12684 29596 12740 29652
rect 12348 29426 12404 29428
rect 12348 29374 12350 29426
rect 12350 29374 12402 29426
rect 12402 29374 12404 29426
rect 12348 29372 12404 29374
rect 12908 29596 12964 29652
rect 12908 28140 12964 28196
rect 12684 27132 12740 27188
rect 12236 27020 12292 27076
rect 12796 26962 12852 26964
rect 12796 26910 12798 26962
rect 12798 26910 12850 26962
rect 12850 26910 12852 26962
rect 12796 26908 12852 26910
rect 13692 35922 13748 35924
rect 13692 35870 13694 35922
rect 13694 35870 13746 35922
rect 13746 35870 13748 35922
rect 13692 35868 13748 35870
rect 13580 35308 13636 35364
rect 14028 35810 14084 35812
rect 14028 35758 14030 35810
rect 14030 35758 14082 35810
rect 14082 35758 14084 35810
rect 14028 35756 14084 35758
rect 13804 35196 13860 35252
rect 14028 35420 14084 35476
rect 13804 34748 13860 34804
rect 13916 34860 13972 34916
rect 14476 35980 14532 36036
rect 14140 35084 14196 35140
rect 14252 35644 14308 35700
rect 14364 35532 14420 35588
rect 14364 35196 14420 35252
rect 13580 33852 13636 33908
rect 14364 34300 14420 34356
rect 14364 34130 14420 34132
rect 14364 34078 14366 34130
rect 14366 34078 14418 34130
rect 14418 34078 14420 34130
rect 14364 34076 14420 34078
rect 14028 33852 14084 33908
rect 14252 33628 14308 33684
rect 14028 33516 14084 33572
rect 13468 31612 13524 31668
rect 13580 33404 13636 33460
rect 13580 33180 13636 33236
rect 13244 31052 13300 31108
rect 13468 30380 13524 30436
rect 13244 29820 13300 29876
rect 13020 27356 13076 27412
rect 13020 27074 13076 27076
rect 13020 27022 13022 27074
rect 13022 27022 13074 27074
rect 13074 27022 13076 27074
rect 13020 27020 13076 27022
rect 12012 26124 12068 26180
rect 12348 26236 12404 26292
rect 12236 24668 12292 24724
rect 12012 24050 12068 24052
rect 12012 23998 12014 24050
rect 12014 23998 12066 24050
rect 12066 23998 12068 24050
rect 12012 23996 12068 23998
rect 11676 23436 11732 23492
rect 11564 23212 11620 23268
rect 11676 22988 11732 23044
rect 11900 23884 11956 23940
rect 11676 21756 11732 21812
rect 11676 20636 11732 20692
rect 11564 20130 11620 20132
rect 11564 20078 11566 20130
rect 11566 20078 11618 20130
rect 11618 20078 11620 20130
rect 11564 20076 11620 20078
rect 12124 23772 12180 23828
rect 12124 23436 12180 23492
rect 12460 26178 12516 26180
rect 12460 26126 12462 26178
rect 12462 26126 12514 26178
rect 12514 26126 12516 26178
rect 12460 26124 12516 26126
rect 12796 25730 12852 25732
rect 12796 25678 12798 25730
rect 12798 25678 12850 25730
rect 12850 25678 12852 25730
rect 12796 25676 12852 25678
rect 12572 25564 12628 25620
rect 13020 24946 13076 24948
rect 13020 24894 13022 24946
rect 13022 24894 13074 24946
rect 13074 24894 13076 24946
rect 13020 24892 13076 24894
rect 12236 23212 12292 23268
rect 12012 22876 12068 22932
rect 11900 20412 11956 20468
rect 12012 21586 12068 21588
rect 12012 21534 12014 21586
rect 12014 21534 12066 21586
rect 12066 21534 12068 21586
rect 12012 21532 12068 21534
rect 11228 19964 11284 20020
rect 12348 22146 12404 22148
rect 12348 22094 12350 22146
rect 12350 22094 12402 22146
rect 12402 22094 12404 22146
rect 12348 22092 12404 22094
rect 12236 21532 12292 21588
rect 13020 23660 13076 23716
rect 12796 22652 12852 22708
rect 12908 22540 12964 22596
rect 12908 21980 12964 22036
rect 12572 20748 12628 20804
rect 11004 18284 11060 18340
rect 11228 19068 11284 19124
rect 11452 19068 11508 19124
rect 11452 18508 11508 18564
rect 11228 16828 11284 16884
rect 10668 14924 10724 14980
rect 11340 18284 11396 18340
rect 10892 14700 10948 14756
rect 9884 12012 9940 12068
rect 10108 12348 10164 12404
rect 10332 12962 10388 12964
rect 10332 12910 10334 12962
rect 10334 12910 10386 12962
rect 10386 12910 10388 12962
rect 10332 12908 10388 12910
rect 10668 13746 10724 13748
rect 10668 13694 10670 13746
rect 10670 13694 10722 13746
rect 10722 13694 10724 13746
rect 10668 13692 10724 13694
rect 10556 13132 10612 13188
rect 10668 13020 10724 13076
rect 10892 13580 10948 13636
rect 10668 12796 10724 12852
rect 10556 12738 10612 12740
rect 10556 12686 10558 12738
rect 10558 12686 10610 12738
rect 10610 12686 10612 12738
rect 10556 12684 10612 12686
rect 10556 12236 10612 12292
rect 10220 12124 10276 12180
rect 8988 11394 9044 11396
rect 8988 11342 8990 11394
rect 8990 11342 9042 11394
rect 9042 11342 9044 11394
rect 8988 11340 9044 11342
rect 8652 11228 8708 11284
rect 8876 11170 8932 11172
rect 8876 11118 8878 11170
rect 8878 11118 8930 11170
rect 8930 11118 8932 11170
rect 8876 11116 8932 11118
rect 9100 10498 9156 10500
rect 9100 10446 9102 10498
rect 9102 10446 9154 10498
rect 9154 10446 9156 10498
rect 9100 10444 9156 10446
rect 8764 9996 8820 10052
rect 8428 9548 8484 9604
rect 8428 7980 8484 8036
rect 9772 9996 9828 10052
rect 9660 9660 9716 9716
rect 11228 14588 11284 14644
rect 11116 14530 11172 14532
rect 11116 14478 11118 14530
rect 11118 14478 11170 14530
rect 11170 14478 11172 14530
rect 11116 14476 11172 14478
rect 11788 18396 11844 18452
rect 11676 17724 11732 17780
rect 11788 17612 11844 17668
rect 11452 17052 11508 17108
rect 11900 16098 11956 16100
rect 11900 16046 11902 16098
rect 11902 16046 11954 16098
rect 11954 16046 11956 16098
rect 11900 16044 11956 16046
rect 11788 15202 11844 15204
rect 11788 15150 11790 15202
rect 11790 15150 11842 15202
rect 11842 15150 11844 15202
rect 11788 15148 11844 15150
rect 12460 19122 12516 19124
rect 12460 19070 12462 19122
rect 12462 19070 12514 19122
rect 12514 19070 12516 19122
rect 12460 19068 12516 19070
rect 12348 18844 12404 18900
rect 12236 17836 12292 17892
rect 12572 18172 12628 18228
rect 12124 17442 12180 17444
rect 12124 17390 12126 17442
rect 12126 17390 12178 17442
rect 12178 17390 12180 17442
rect 12124 17388 12180 17390
rect 12572 17554 12628 17556
rect 12572 17502 12574 17554
rect 12574 17502 12626 17554
rect 12626 17502 12628 17554
rect 12572 17500 12628 17502
rect 12460 16268 12516 16324
rect 13020 21196 13076 21252
rect 12908 20802 12964 20804
rect 12908 20750 12910 20802
rect 12910 20750 12962 20802
rect 12962 20750 12964 20802
rect 12908 20748 12964 20750
rect 13356 27356 13412 27412
rect 13692 33122 13748 33124
rect 13692 33070 13694 33122
rect 13694 33070 13746 33122
rect 13746 33070 13748 33122
rect 13692 33068 13748 33070
rect 14812 36428 14868 36484
rect 14812 35138 14868 35140
rect 14812 35086 14814 35138
rect 14814 35086 14866 35138
rect 14866 35086 14868 35138
rect 14812 35084 14868 35086
rect 14700 34860 14756 34916
rect 15036 38892 15092 38948
rect 15260 39452 15316 39508
rect 15596 39340 15652 39396
rect 15260 38892 15316 38948
rect 15484 38892 15540 38948
rect 15372 38050 15428 38052
rect 15372 37998 15374 38050
rect 15374 37998 15426 38050
rect 15426 37998 15428 38050
rect 15372 37996 15428 37998
rect 15036 36988 15092 37044
rect 15036 36482 15092 36484
rect 15036 36430 15038 36482
rect 15038 36430 15090 36482
rect 15090 36430 15092 36482
rect 15036 36428 15092 36430
rect 15148 36092 15204 36148
rect 15596 37884 15652 37940
rect 16828 40684 16884 40740
rect 17612 44044 17668 44100
rect 17500 42530 17556 42532
rect 17500 42478 17502 42530
rect 17502 42478 17554 42530
rect 17554 42478 17556 42530
rect 17500 42476 17556 42478
rect 17388 41804 17444 41860
rect 18620 44994 18676 44996
rect 18620 44942 18622 44994
rect 18622 44942 18674 44994
rect 18674 44942 18676 44994
rect 18620 44940 18676 44942
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 17948 44044 18004 44100
rect 20076 44098 20132 44100
rect 20076 44046 20078 44098
rect 20078 44046 20130 44098
rect 20130 44046 20132 44098
rect 20076 44044 20132 44046
rect 20524 44098 20580 44100
rect 20524 44046 20526 44098
rect 20526 44046 20578 44098
rect 20578 44046 20580 44098
rect 20524 44044 20580 44046
rect 21308 44940 21364 44996
rect 21868 44994 21924 44996
rect 21868 44942 21870 44994
rect 21870 44942 21922 44994
rect 21922 44942 21924 44994
rect 21868 44940 21924 44942
rect 21084 44044 21140 44100
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 18172 43426 18228 43428
rect 18172 43374 18174 43426
rect 18174 43374 18226 43426
rect 18226 43374 18228 43426
rect 18172 43372 18228 43374
rect 17948 42924 18004 42980
rect 18956 42978 19012 42980
rect 18956 42926 18958 42978
rect 18958 42926 19010 42978
rect 19010 42926 19012 42978
rect 18956 42924 19012 42926
rect 20860 43426 20916 43428
rect 20860 43374 20862 43426
rect 20862 43374 20914 43426
rect 20914 43374 20916 43426
rect 20860 43372 20916 43374
rect 20300 42700 20356 42756
rect 17500 41916 17556 41972
rect 19180 42476 19236 42532
rect 18396 41970 18452 41972
rect 18396 41918 18398 41970
rect 18398 41918 18450 41970
rect 18450 41918 18452 41970
rect 18396 41916 18452 41918
rect 17500 40908 17556 40964
rect 15820 40124 15876 40180
rect 15932 39058 15988 39060
rect 15932 39006 15934 39058
rect 15934 39006 15986 39058
rect 15986 39006 15988 39058
rect 15932 39004 15988 39006
rect 16044 38834 16100 38836
rect 16044 38782 16046 38834
rect 16046 38782 16098 38834
rect 16098 38782 16100 38834
rect 16044 38780 16100 38782
rect 16604 40012 16660 40068
rect 16380 38892 16436 38948
rect 16940 38780 16996 38836
rect 17276 39676 17332 39732
rect 17388 39394 17444 39396
rect 17388 39342 17390 39394
rect 17390 39342 17442 39394
rect 17442 39342 17444 39394
rect 17388 39340 17444 39342
rect 19068 41858 19124 41860
rect 19068 41806 19070 41858
rect 19070 41806 19122 41858
rect 19122 41806 19124 41858
rect 19068 41804 19124 41806
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 25228 46114 25284 46116
rect 25228 46062 25230 46114
rect 25230 46062 25282 46114
rect 25282 46062 25284 46114
rect 25228 46060 25284 46062
rect 27132 45388 27188 45444
rect 30940 45330 30996 45332
rect 30940 45278 30942 45330
rect 30942 45278 30994 45330
rect 30994 45278 30996 45330
rect 30940 45276 30996 45278
rect 21868 44098 21924 44100
rect 21868 44046 21870 44098
rect 21870 44046 21922 44098
rect 21922 44046 21924 44098
rect 21868 44044 21924 44046
rect 22316 44098 22372 44100
rect 22316 44046 22318 44098
rect 22318 44046 22370 44098
rect 22370 44046 22372 44098
rect 22316 44044 22372 44046
rect 22988 44098 23044 44100
rect 22988 44046 22990 44098
rect 22990 44046 23042 44098
rect 23042 44046 23044 44098
rect 22988 44044 23044 44046
rect 21420 43484 21476 43540
rect 21420 42754 21476 42756
rect 21420 42702 21422 42754
rect 21422 42702 21474 42754
rect 21474 42702 21476 42754
rect 21420 42700 21476 42702
rect 21308 42530 21364 42532
rect 21308 42478 21310 42530
rect 21310 42478 21362 42530
rect 21362 42478 21364 42530
rect 21308 42476 21364 42478
rect 20524 41970 20580 41972
rect 20524 41918 20526 41970
rect 20526 41918 20578 41970
rect 20578 41918 20580 41970
rect 20524 41916 20580 41918
rect 21420 41916 21476 41972
rect 19404 41804 19460 41860
rect 21532 41804 21588 41860
rect 18284 40684 18340 40740
rect 18396 40908 18452 40964
rect 20524 40962 20580 40964
rect 20524 40910 20526 40962
rect 20526 40910 20578 40962
rect 20578 40910 20580 40962
rect 20524 40908 20580 40910
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 18172 40012 18228 40068
rect 17724 38834 17780 38836
rect 17724 38782 17726 38834
rect 17726 38782 17778 38834
rect 17778 38782 17780 38834
rect 17724 38780 17780 38782
rect 16268 38332 16324 38388
rect 15708 37772 15764 37828
rect 15484 36092 15540 36148
rect 15036 35308 15092 35364
rect 15260 34524 15316 34580
rect 15372 34972 15428 35028
rect 15036 34412 15092 34468
rect 15148 34188 15204 34244
rect 15036 33628 15092 33684
rect 14028 32844 14084 32900
rect 16268 37100 16324 37156
rect 16604 38332 16660 38388
rect 16380 36988 16436 37044
rect 15820 34188 15876 34244
rect 13692 31612 13748 31668
rect 13692 30716 13748 30772
rect 14476 32284 14532 32340
rect 14476 31836 14532 31892
rect 14140 29986 14196 29988
rect 14140 29934 14142 29986
rect 14142 29934 14194 29986
rect 14194 29934 14196 29986
rect 14140 29932 14196 29934
rect 14252 31724 14308 31780
rect 13916 29708 13972 29764
rect 13580 29538 13636 29540
rect 13580 29486 13582 29538
rect 13582 29486 13634 29538
rect 13634 29486 13636 29538
rect 13580 29484 13636 29486
rect 13580 28754 13636 28756
rect 13580 28702 13582 28754
rect 13582 28702 13634 28754
rect 13634 28702 13636 28754
rect 13580 28700 13636 28702
rect 14588 31778 14644 31780
rect 14588 31726 14590 31778
rect 14590 31726 14642 31778
rect 14642 31726 14644 31778
rect 14588 31724 14644 31726
rect 14476 31052 14532 31108
rect 16044 34412 16100 34468
rect 16156 35308 16212 35364
rect 16044 34076 16100 34132
rect 14924 33234 14980 33236
rect 14924 33182 14926 33234
rect 14926 33182 14978 33234
rect 14978 33182 14980 33234
rect 14924 33180 14980 33182
rect 15372 32786 15428 32788
rect 15372 32734 15374 32786
rect 15374 32734 15426 32786
rect 15426 32734 15428 32786
rect 15372 32732 15428 32734
rect 14924 32284 14980 32340
rect 14924 30940 14980 30996
rect 15260 32562 15316 32564
rect 15260 32510 15262 32562
rect 15262 32510 15314 32562
rect 15314 32510 15316 32562
rect 15260 32508 15316 32510
rect 15596 32284 15652 32340
rect 15596 31612 15652 31668
rect 15372 30994 15428 30996
rect 15372 30942 15374 30994
rect 15374 30942 15426 30994
rect 15426 30942 15428 30994
rect 15372 30940 15428 30942
rect 15260 30380 15316 30436
rect 15148 30268 15204 30324
rect 14812 29820 14868 29876
rect 14252 27970 14308 27972
rect 14252 27918 14254 27970
rect 14254 27918 14306 27970
rect 14306 27918 14308 27970
rect 14252 27916 14308 27918
rect 13580 27468 13636 27524
rect 13356 26348 13412 26404
rect 13692 25564 13748 25620
rect 13692 25394 13748 25396
rect 13692 25342 13694 25394
rect 13694 25342 13746 25394
rect 13746 25342 13748 25394
rect 13692 25340 13748 25342
rect 14140 27804 14196 27860
rect 13916 25788 13972 25844
rect 13804 24780 13860 24836
rect 13580 24444 13636 24500
rect 13468 23938 13524 23940
rect 13468 23886 13470 23938
rect 13470 23886 13522 23938
rect 13522 23886 13524 23938
rect 13468 23884 13524 23886
rect 14028 24722 14084 24724
rect 14028 24670 14030 24722
rect 14030 24670 14082 24722
rect 14082 24670 14084 24722
rect 14028 24668 14084 24670
rect 13804 24220 13860 24276
rect 13468 23660 13524 23716
rect 13692 22316 13748 22372
rect 13244 21644 13300 21700
rect 13244 20972 13300 21028
rect 13132 20524 13188 20580
rect 13468 19964 13524 20020
rect 12796 18284 12852 18340
rect 13356 18284 13412 18340
rect 13244 17836 13300 17892
rect 13132 16770 13188 16772
rect 13132 16718 13134 16770
rect 13134 16718 13186 16770
rect 13186 16718 13188 16770
rect 13132 16716 13188 16718
rect 12348 15820 12404 15876
rect 12348 15596 12404 15652
rect 11116 13580 11172 13636
rect 11340 13634 11396 13636
rect 11340 13582 11342 13634
rect 11342 13582 11394 13634
rect 11394 13582 11396 13634
rect 11340 13580 11396 13582
rect 11228 13244 11284 13300
rect 11564 14812 11620 14868
rect 11900 14700 11956 14756
rect 11452 13074 11508 13076
rect 11452 13022 11454 13074
rect 11454 13022 11506 13074
rect 11506 13022 11508 13074
rect 11452 13020 11508 13022
rect 10892 12124 10948 12180
rect 10220 11788 10276 11844
rect 10108 9938 10164 9940
rect 10108 9886 10110 9938
rect 10110 9886 10162 9938
rect 10162 9886 10164 9938
rect 10108 9884 10164 9886
rect 10332 9772 10388 9828
rect 10556 11676 10612 11732
rect 11228 11900 11284 11956
rect 11788 12684 11844 12740
rect 11676 12402 11732 12404
rect 11676 12350 11678 12402
rect 11678 12350 11730 12402
rect 11730 12350 11732 12402
rect 11676 12348 11732 12350
rect 11452 11788 11508 11844
rect 10668 11394 10724 11396
rect 10668 11342 10670 11394
rect 10670 11342 10722 11394
rect 10722 11342 10724 11394
rect 10668 11340 10724 11342
rect 10556 11228 10612 11284
rect 11116 11394 11172 11396
rect 11116 11342 11118 11394
rect 11118 11342 11170 11394
rect 11170 11342 11172 11394
rect 11116 11340 11172 11342
rect 11340 11340 11396 11396
rect 11228 11282 11284 11284
rect 11228 11230 11230 11282
rect 11230 11230 11282 11282
rect 11282 11230 11284 11282
rect 11228 11228 11284 11230
rect 12124 14252 12180 14308
rect 12236 14700 12292 14756
rect 12236 14028 12292 14084
rect 12124 13580 12180 13636
rect 12236 13020 12292 13076
rect 12684 15596 12740 15652
rect 12572 14924 12628 14980
rect 12572 14476 12628 14532
rect 12684 14812 12740 14868
rect 13244 15484 13300 15540
rect 12796 14418 12852 14420
rect 12796 14366 12798 14418
rect 12798 14366 12850 14418
rect 12850 14366 12852 14418
rect 12796 14364 12852 14366
rect 12908 14306 12964 14308
rect 12908 14254 12910 14306
rect 12910 14254 12962 14306
rect 12962 14254 12964 14306
rect 12908 14252 12964 14254
rect 11900 12572 11956 12628
rect 12236 12684 12292 12740
rect 11788 11900 11844 11956
rect 12348 12178 12404 12180
rect 12348 12126 12350 12178
rect 12350 12126 12402 12178
rect 12402 12126 12404 12178
rect 12348 12124 12404 12126
rect 12572 12850 12628 12852
rect 12572 12798 12574 12850
rect 12574 12798 12626 12850
rect 12626 12798 12628 12850
rect 12572 12796 12628 12798
rect 12236 11676 12292 11732
rect 11900 11340 11956 11396
rect 12124 11564 12180 11620
rect 12460 11506 12516 11508
rect 12460 11454 12462 11506
rect 12462 11454 12514 11506
rect 12514 11454 12516 11506
rect 12460 11452 12516 11454
rect 12012 11282 12068 11284
rect 12012 11230 12014 11282
rect 12014 11230 12066 11282
rect 12066 11230 12068 11282
rect 12012 11228 12068 11230
rect 11788 11116 11844 11172
rect 11452 10892 11508 10948
rect 11340 10556 11396 10612
rect 8764 8818 8820 8820
rect 8764 8766 8766 8818
rect 8766 8766 8818 8818
rect 8818 8766 8820 8818
rect 8764 8764 8820 8766
rect 8876 8652 8932 8708
rect 9324 9436 9380 9492
rect 7980 6972 8036 7028
rect 7756 5964 7812 6020
rect 7644 5906 7700 5908
rect 7644 5854 7646 5906
rect 7646 5854 7698 5906
rect 7698 5854 7700 5906
rect 7644 5852 7700 5854
rect 7644 5404 7700 5460
rect 7868 6748 7924 6804
rect 8092 6076 8148 6132
rect 8316 6466 8372 6468
rect 8316 6414 8318 6466
rect 8318 6414 8370 6466
rect 8370 6414 8372 6466
rect 8316 6412 8372 6414
rect 8540 6300 8596 6356
rect 8428 6018 8484 6020
rect 8428 5966 8430 6018
rect 8430 5966 8482 6018
rect 8482 5966 8484 6018
rect 8428 5964 8484 5966
rect 8540 5852 8596 5908
rect 8092 5292 8148 5348
rect 7980 5122 8036 5124
rect 7980 5070 7982 5122
rect 7982 5070 8034 5122
rect 8034 5070 8036 5122
rect 7980 5068 8036 5070
rect 8652 5740 8708 5796
rect 8764 5404 8820 5460
rect 8652 5068 8708 5124
rect 8764 4956 8820 5012
rect 8316 4844 8372 4900
rect 8428 4732 8484 4788
rect 9100 8258 9156 8260
rect 9100 8206 9102 8258
rect 9102 8206 9154 8258
rect 9154 8206 9156 8258
rect 9100 8204 9156 8206
rect 8988 7308 9044 7364
rect 9212 7420 9268 7476
rect 9100 6860 9156 6916
rect 9324 6748 9380 6804
rect 9436 7868 9492 7924
rect 9212 6690 9268 6692
rect 9212 6638 9214 6690
rect 9214 6638 9266 6690
rect 9266 6638 9268 6690
rect 9212 6636 9268 6638
rect 8988 6524 9044 6580
rect 9324 6466 9380 6468
rect 9324 6414 9326 6466
rect 9326 6414 9378 6466
rect 9378 6414 9380 6466
rect 9324 6412 9380 6414
rect 8988 6076 9044 6132
rect 8988 5906 9044 5908
rect 8988 5854 8990 5906
rect 8990 5854 9042 5906
rect 9042 5854 9044 5906
rect 8988 5852 9044 5854
rect 8876 3666 8932 3668
rect 8876 3614 8878 3666
rect 8878 3614 8930 3666
rect 8930 3614 8932 3666
rect 8876 3612 8932 3614
rect 4060 3276 4116 3332
rect 3388 2828 3444 2884
rect 9324 2940 9380 2996
rect 9772 7532 9828 7588
rect 10332 9548 10388 9604
rect 12012 9938 12068 9940
rect 12012 9886 12014 9938
rect 12014 9886 12066 9938
rect 12066 9886 12068 9938
rect 12012 9884 12068 9886
rect 11004 9436 11060 9492
rect 11228 8988 11284 9044
rect 10220 8540 10276 8596
rect 10780 8316 10836 8372
rect 10108 8204 10164 8260
rect 10444 8146 10500 8148
rect 10444 8094 10446 8146
rect 10446 8094 10498 8146
rect 10498 8094 10500 8146
rect 10444 8092 10500 8094
rect 10220 8034 10276 8036
rect 10220 7982 10222 8034
rect 10222 7982 10274 8034
rect 10274 7982 10276 8034
rect 10220 7980 10276 7982
rect 10332 7698 10388 7700
rect 10332 7646 10334 7698
rect 10334 7646 10386 7698
rect 10386 7646 10388 7698
rect 10332 7644 10388 7646
rect 9996 7420 10052 7476
rect 10892 7698 10948 7700
rect 10892 7646 10894 7698
rect 10894 7646 10946 7698
rect 10946 7646 10948 7698
rect 10892 7644 10948 7646
rect 10780 7586 10836 7588
rect 10780 7534 10782 7586
rect 10782 7534 10834 7586
rect 10834 7534 10836 7586
rect 10780 7532 10836 7534
rect 9772 6748 9828 6804
rect 10668 7308 10724 7364
rect 9548 6690 9604 6692
rect 9548 6638 9550 6690
rect 9550 6638 9602 6690
rect 9602 6638 9604 6690
rect 9548 6636 9604 6638
rect 9660 6524 9716 6580
rect 10108 6300 10164 6356
rect 12460 10892 12516 10948
rect 11676 8316 11732 8372
rect 11228 7084 11284 7140
rect 9772 6130 9828 6132
rect 9772 6078 9774 6130
rect 9774 6078 9826 6130
rect 9826 6078 9828 6130
rect 9772 6076 9828 6078
rect 9660 5852 9716 5908
rect 9548 5122 9604 5124
rect 9548 5070 9550 5122
rect 9550 5070 9602 5122
rect 9602 5070 9604 5122
rect 9548 5068 9604 5070
rect 10220 5906 10276 5908
rect 10220 5854 10222 5906
rect 10222 5854 10274 5906
rect 10274 5854 10276 5906
rect 10220 5852 10276 5854
rect 10668 6300 10724 6356
rect 9996 5628 10052 5684
rect 11004 6578 11060 6580
rect 11004 6526 11006 6578
rect 11006 6526 11058 6578
rect 11058 6526 11060 6578
rect 11004 6524 11060 6526
rect 10892 6076 10948 6132
rect 10668 5628 10724 5684
rect 10892 5852 10948 5908
rect 10892 5516 10948 5572
rect 11004 5180 11060 5236
rect 11228 6412 11284 6468
rect 11452 6018 11508 6020
rect 11452 5966 11454 6018
rect 11454 5966 11506 6018
rect 11506 5966 11508 6018
rect 11452 5964 11508 5966
rect 11228 5740 11284 5796
rect 11116 5292 11172 5348
rect 10220 5068 10276 5124
rect 9772 4732 9828 4788
rect 9884 4956 9940 5012
rect 9884 4562 9940 4564
rect 9884 4510 9886 4562
rect 9886 4510 9938 4562
rect 9938 4510 9940 4562
rect 9884 4508 9940 4510
rect 10444 4732 10500 4788
rect 9996 3724 10052 3780
rect 10780 4620 10836 4676
rect 11452 5740 11508 5796
rect 10780 3612 10836 3668
rect 9548 3442 9604 3444
rect 9548 3390 9550 3442
rect 9550 3390 9602 3442
rect 9602 3390 9604 3442
rect 9548 3388 9604 3390
rect 9548 2716 9604 2772
rect 6748 2268 6804 2324
rect 12012 8316 12068 8372
rect 12348 7644 12404 7700
rect 11676 5964 11732 6020
rect 12684 10668 12740 10724
rect 13020 11954 13076 11956
rect 13020 11902 13022 11954
rect 13022 11902 13074 11954
rect 13074 11902 13076 11954
rect 13020 11900 13076 11902
rect 13132 11788 13188 11844
rect 12908 10444 12964 10500
rect 13020 11676 13076 11732
rect 12908 9996 12964 10052
rect 12908 8930 12964 8932
rect 12908 8878 12910 8930
rect 12910 8878 12962 8930
rect 12962 8878 12964 8930
rect 12908 8876 12964 8878
rect 12684 8652 12740 8708
rect 12796 8540 12852 8596
rect 12796 8146 12852 8148
rect 12796 8094 12798 8146
rect 12798 8094 12850 8146
rect 12850 8094 12852 8146
rect 12796 8092 12852 8094
rect 12572 6578 12628 6580
rect 12572 6526 12574 6578
rect 12574 6526 12626 6578
rect 12626 6526 12628 6578
rect 12572 6524 12628 6526
rect 12572 5682 12628 5684
rect 12572 5630 12574 5682
rect 12574 5630 12626 5682
rect 12626 5630 12628 5682
rect 12572 5628 12628 5630
rect 12236 5404 12292 5460
rect 12460 5516 12516 5572
rect 12348 5180 12404 5236
rect 12572 5404 12628 5460
rect 12684 5068 12740 5124
rect 12908 7756 12964 7812
rect 13468 17164 13524 17220
rect 14252 26402 14308 26404
rect 14252 26350 14254 26402
rect 14254 26350 14306 26402
rect 14306 26350 14308 26402
rect 14252 26348 14308 26350
rect 14252 25618 14308 25620
rect 14252 25566 14254 25618
rect 14254 25566 14306 25618
rect 14306 25566 14308 25618
rect 14252 25564 14308 25566
rect 16268 35084 16324 35140
rect 15932 32844 15988 32900
rect 15820 30994 15876 30996
rect 15820 30942 15822 30994
rect 15822 30942 15874 30994
rect 15874 30942 15876 30994
rect 15820 30940 15876 30942
rect 16156 32732 16212 32788
rect 16268 33852 16324 33908
rect 16156 31724 16212 31780
rect 16380 32562 16436 32564
rect 16380 32510 16382 32562
rect 16382 32510 16434 32562
rect 16434 32510 16436 32562
rect 16380 32508 16436 32510
rect 16604 35196 16660 35252
rect 16716 35420 16772 35476
rect 16604 34914 16660 34916
rect 16604 34862 16606 34914
rect 16606 34862 16658 34914
rect 16658 34862 16660 34914
rect 16604 34860 16660 34862
rect 16156 31106 16212 31108
rect 16156 31054 16158 31106
rect 16158 31054 16210 31106
rect 16210 31054 16212 31106
rect 16156 31052 16212 31054
rect 15932 30210 15988 30212
rect 15932 30158 15934 30210
rect 15934 30158 15986 30210
rect 15986 30158 15988 30210
rect 15932 30156 15988 30158
rect 16268 30716 16324 30772
rect 15820 29820 15876 29876
rect 15148 27858 15204 27860
rect 15148 27806 15150 27858
rect 15150 27806 15202 27858
rect 15202 27806 15204 27858
rect 15148 27804 15204 27806
rect 15260 28476 15316 28532
rect 14364 25228 14420 25284
rect 14588 26684 14644 26740
rect 14140 24610 14196 24612
rect 14140 24558 14142 24610
rect 14142 24558 14194 24610
rect 14194 24558 14196 24610
rect 14140 24556 14196 24558
rect 15148 26348 15204 26404
rect 14700 25676 14756 25732
rect 15036 25228 15092 25284
rect 14812 24780 14868 24836
rect 14588 24332 14644 24388
rect 14140 24050 14196 24052
rect 14140 23998 14142 24050
rect 14142 23998 14194 24050
rect 14194 23998 14196 24050
rect 14140 23996 14196 23998
rect 14252 23436 14308 23492
rect 14140 21980 14196 22036
rect 14476 23042 14532 23044
rect 14476 22990 14478 23042
rect 14478 22990 14530 23042
rect 14530 22990 14532 23042
rect 14476 22988 14532 22990
rect 14028 20578 14084 20580
rect 14028 20526 14030 20578
rect 14030 20526 14082 20578
rect 14082 20526 14084 20578
rect 14028 20524 14084 20526
rect 14252 20076 14308 20132
rect 14700 24668 14756 24724
rect 14924 24556 14980 24612
rect 15148 22594 15204 22596
rect 15148 22542 15150 22594
rect 15150 22542 15202 22594
rect 15202 22542 15204 22594
rect 15148 22540 15204 22542
rect 15484 28924 15540 28980
rect 15484 27746 15540 27748
rect 15484 27694 15486 27746
rect 15486 27694 15538 27746
rect 15538 27694 15540 27746
rect 15484 27692 15540 27694
rect 15932 28812 15988 28868
rect 15596 26684 15652 26740
rect 15708 26908 15764 26964
rect 16268 30156 16324 30212
rect 19068 40290 19124 40292
rect 19068 40238 19070 40290
rect 19070 40238 19122 40290
rect 19122 40238 19124 40290
rect 19068 40236 19124 40238
rect 20188 40124 20244 40180
rect 19404 40012 19460 40068
rect 19964 39730 20020 39732
rect 19964 39678 19966 39730
rect 19966 39678 20018 39730
rect 20018 39678 20020 39730
rect 19964 39676 20020 39678
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 18844 38780 18900 38836
rect 18172 37938 18228 37940
rect 18172 37886 18174 37938
rect 18174 37886 18226 37938
rect 18226 37886 18228 37938
rect 18172 37884 18228 37886
rect 17948 37660 18004 37716
rect 17500 37266 17556 37268
rect 17500 37214 17502 37266
rect 17502 37214 17554 37266
rect 17554 37214 17556 37266
rect 17500 37212 17556 37214
rect 17500 36988 17556 37044
rect 17388 35698 17444 35700
rect 17388 35646 17390 35698
rect 17390 35646 17442 35698
rect 17442 35646 17444 35698
rect 17388 35644 17444 35646
rect 17276 34860 17332 34916
rect 17164 33292 17220 33348
rect 16716 32844 16772 32900
rect 16716 32620 16772 32676
rect 16604 31778 16660 31780
rect 16604 31726 16606 31778
rect 16606 31726 16658 31778
rect 16658 31726 16660 31778
rect 16604 31724 16660 31726
rect 16492 30210 16548 30212
rect 16492 30158 16494 30210
rect 16494 30158 16546 30210
rect 16546 30158 16548 30210
rect 16492 30156 16548 30158
rect 17612 34524 17668 34580
rect 17724 34242 17780 34244
rect 17724 34190 17726 34242
rect 17726 34190 17778 34242
rect 17778 34190 17780 34242
rect 17724 34188 17780 34190
rect 17836 34130 17892 34132
rect 17836 34078 17838 34130
rect 17838 34078 17890 34130
rect 17890 34078 17892 34130
rect 17836 34076 17892 34078
rect 17500 32508 17556 32564
rect 17388 31724 17444 31780
rect 16492 28252 16548 28308
rect 15820 26460 15876 26516
rect 15932 26684 15988 26740
rect 16156 26572 16212 26628
rect 16156 26236 16212 26292
rect 15484 25116 15540 25172
rect 15596 23772 15652 23828
rect 15932 23772 15988 23828
rect 15708 23548 15764 23604
rect 15372 22764 15428 22820
rect 15484 22988 15540 23044
rect 15372 22146 15428 22148
rect 15372 22094 15374 22146
rect 15374 22094 15426 22146
rect 15426 22094 15428 22146
rect 15372 22092 15428 22094
rect 14924 21756 14980 21812
rect 14924 21084 14980 21140
rect 14812 20412 14868 20468
rect 15372 21420 15428 21476
rect 14588 18620 14644 18676
rect 13804 17164 13860 17220
rect 14588 18450 14644 18452
rect 14588 18398 14590 18450
rect 14590 18398 14642 18450
rect 14642 18398 14644 18450
rect 14588 18396 14644 18398
rect 14588 18060 14644 18116
rect 14140 17778 14196 17780
rect 14140 17726 14142 17778
rect 14142 17726 14194 17778
rect 14194 17726 14196 17778
rect 14140 17724 14196 17726
rect 14364 17724 14420 17780
rect 14924 17666 14980 17668
rect 14924 17614 14926 17666
rect 14926 17614 14978 17666
rect 14978 17614 14980 17666
rect 14924 17612 14980 17614
rect 14700 17554 14756 17556
rect 14700 17502 14702 17554
rect 14702 17502 14754 17554
rect 14754 17502 14756 17554
rect 14700 17500 14756 17502
rect 14364 16940 14420 16996
rect 14700 17164 14756 17220
rect 13804 16882 13860 16884
rect 13804 16830 13806 16882
rect 13806 16830 13858 16882
rect 13858 16830 13860 16882
rect 13804 16828 13860 16830
rect 14588 16716 14644 16772
rect 14140 16268 14196 16324
rect 13580 15932 13636 15988
rect 13468 15148 13524 15204
rect 13916 15260 13972 15316
rect 13804 14028 13860 14084
rect 13916 13692 13972 13748
rect 13356 12348 13412 12404
rect 13804 13244 13860 13300
rect 13468 12124 13524 12180
rect 14028 13356 14084 13412
rect 13916 12572 13972 12628
rect 13804 12460 13860 12516
rect 13804 11676 13860 11732
rect 13356 10892 13412 10948
rect 14028 12124 14084 12180
rect 14252 14418 14308 14420
rect 14252 14366 14254 14418
rect 14254 14366 14306 14418
rect 14306 14366 14308 14418
rect 14252 14364 14308 14366
rect 14812 16940 14868 16996
rect 14700 16380 14756 16436
rect 14476 14140 14532 14196
rect 15260 20972 15316 21028
rect 16044 22876 16100 22932
rect 15484 20188 15540 20244
rect 15596 22092 15652 22148
rect 15820 20860 15876 20916
rect 15932 20972 15988 21028
rect 15708 20636 15764 20692
rect 15708 20242 15764 20244
rect 15708 20190 15710 20242
rect 15710 20190 15762 20242
rect 15762 20190 15764 20242
rect 15708 20188 15764 20190
rect 15932 20412 15988 20468
rect 15596 19628 15652 19684
rect 15036 15708 15092 15764
rect 15148 18508 15204 18564
rect 15372 16828 15428 16884
rect 14812 14252 14868 14308
rect 14364 13580 14420 13636
rect 14252 13244 14308 13300
rect 14364 13132 14420 13188
rect 14588 12850 14644 12852
rect 14588 12798 14590 12850
rect 14590 12798 14642 12850
rect 14642 12798 14644 12850
rect 14588 12796 14644 12798
rect 14588 12402 14644 12404
rect 14588 12350 14590 12402
rect 14590 12350 14642 12402
rect 14642 12350 14644 12402
rect 14588 12348 14644 12350
rect 14476 12290 14532 12292
rect 14476 12238 14478 12290
rect 14478 12238 14530 12290
rect 14530 12238 14532 12290
rect 14476 12236 14532 12238
rect 14364 12124 14420 12180
rect 14364 11676 14420 11732
rect 14588 11564 14644 11620
rect 14028 10834 14084 10836
rect 14028 10782 14030 10834
rect 14030 10782 14082 10834
rect 14082 10782 14084 10834
rect 14028 10780 14084 10782
rect 13468 10444 13524 10500
rect 13580 10668 13636 10724
rect 13804 10444 13860 10500
rect 13804 8652 13860 8708
rect 13244 8540 13300 8596
rect 12908 6076 12964 6132
rect 11564 4620 11620 4676
rect 12236 4620 12292 4676
rect 12796 4844 12852 4900
rect 14028 8764 14084 8820
rect 13916 8428 13972 8484
rect 13468 8092 13524 8148
rect 13468 7532 13524 7588
rect 13804 8204 13860 8260
rect 14476 11004 14532 11060
rect 14588 10780 14644 10836
rect 14476 10610 14532 10612
rect 14476 10558 14478 10610
rect 14478 10558 14530 10610
rect 14530 10558 14532 10610
rect 14476 10556 14532 10558
rect 14812 11228 14868 11284
rect 15260 13970 15316 13972
rect 15260 13918 15262 13970
rect 15262 13918 15314 13970
rect 15314 13918 15316 13970
rect 15260 13916 15316 13918
rect 15036 12348 15092 12404
rect 15148 12796 15204 12852
rect 15484 13468 15540 13524
rect 15036 11900 15092 11956
rect 14812 11004 14868 11060
rect 14476 8930 14532 8932
rect 14476 8878 14478 8930
rect 14478 8878 14530 8930
rect 14530 8878 14532 8930
rect 14476 8876 14532 8878
rect 14252 7308 14308 7364
rect 15036 11676 15092 11732
rect 15708 16716 15764 16772
rect 16604 26684 16660 26740
rect 16940 30380 16996 30436
rect 16492 26572 16548 26628
rect 16380 26460 16436 26516
rect 16940 28924 16996 28980
rect 17164 31164 17220 31220
rect 17500 30828 17556 30884
rect 17276 30770 17332 30772
rect 17276 30718 17278 30770
rect 17278 30718 17330 30770
rect 17330 30718 17332 30770
rect 17276 30716 17332 30718
rect 20076 38780 20132 38836
rect 18396 37660 18452 37716
rect 18396 36988 18452 37044
rect 18172 36204 18228 36260
rect 18284 35644 18340 35700
rect 18060 34076 18116 34132
rect 18284 34130 18340 34132
rect 18284 34078 18286 34130
rect 18286 34078 18338 34130
rect 18338 34078 18340 34130
rect 18284 34076 18340 34078
rect 18172 33292 18228 33348
rect 18172 31948 18228 32004
rect 18844 37100 18900 37156
rect 18844 36482 18900 36484
rect 18844 36430 18846 36482
rect 18846 36430 18898 36482
rect 18898 36430 18900 36482
rect 18844 36428 18900 36430
rect 19068 36764 19124 36820
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19404 36652 19460 36708
rect 19852 36988 19908 37044
rect 20524 39788 20580 39844
rect 20972 40348 21028 40404
rect 20748 39618 20804 39620
rect 20748 39566 20750 39618
rect 20750 39566 20802 39618
rect 20802 39566 20804 39618
rect 20748 39564 20804 39566
rect 21532 40348 21588 40404
rect 21196 39788 21252 39844
rect 21420 40236 21476 40292
rect 21756 42476 21812 42532
rect 22428 43426 22484 43428
rect 22428 43374 22430 43426
rect 22430 43374 22482 43426
rect 22482 43374 22484 43426
rect 22428 43372 22484 43374
rect 22316 42476 22372 42532
rect 24220 43650 24276 43652
rect 24220 43598 24222 43650
rect 24222 43598 24274 43650
rect 24274 43598 24276 43650
rect 24220 43596 24276 43598
rect 22876 42140 22932 42196
rect 24332 43484 24388 43540
rect 23996 43372 24052 43428
rect 23436 43260 23492 43316
rect 23660 42866 23716 42868
rect 23660 42814 23662 42866
rect 23662 42814 23714 42866
rect 23714 42814 23716 42866
rect 23660 42812 23716 42814
rect 23324 42194 23380 42196
rect 23324 42142 23326 42194
rect 23326 42142 23378 42194
rect 23378 42142 23380 42194
rect 23324 42140 23380 42142
rect 22204 41804 22260 41860
rect 23212 41858 23268 41860
rect 23212 41806 23214 41858
rect 23214 41806 23266 41858
rect 23266 41806 23268 41858
rect 23212 41804 23268 41806
rect 23772 41692 23828 41748
rect 21980 40402 22036 40404
rect 21980 40350 21982 40402
rect 21982 40350 22034 40402
rect 22034 40350 22036 40402
rect 21980 40348 22036 40350
rect 20748 38834 20804 38836
rect 20748 38782 20750 38834
rect 20750 38782 20802 38834
rect 20802 38782 20804 38834
rect 20748 38780 20804 38782
rect 20412 38722 20468 38724
rect 20412 38670 20414 38722
rect 20414 38670 20466 38722
rect 20466 38670 20468 38722
rect 20412 38668 20468 38670
rect 20300 38556 20356 38612
rect 20972 38556 21028 38612
rect 21420 38668 21476 38724
rect 20748 37826 20804 37828
rect 20748 37774 20750 37826
rect 20750 37774 20802 37826
rect 20802 37774 20804 37826
rect 20748 37772 20804 37774
rect 19180 36540 19236 36596
rect 19068 36258 19124 36260
rect 19068 36206 19070 36258
rect 19070 36206 19122 36258
rect 19122 36206 19124 36258
rect 19068 36204 19124 36206
rect 18956 35644 19012 35700
rect 19180 35532 19236 35588
rect 19516 36204 19572 36260
rect 19740 36370 19796 36372
rect 19740 36318 19742 36370
rect 19742 36318 19794 36370
rect 19794 36318 19796 36370
rect 19740 36316 19796 36318
rect 20188 36764 20244 36820
rect 19964 36482 20020 36484
rect 19964 36430 19966 36482
rect 19966 36430 20018 36482
rect 20018 36430 20020 36482
rect 19964 36428 20020 36430
rect 19852 36204 19908 36260
rect 20748 36988 20804 37044
rect 20412 36540 20468 36596
rect 20188 36204 20244 36260
rect 19836 36090 19892 36092
rect 19628 35980 19684 36036
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19516 35138 19572 35140
rect 19516 35086 19518 35138
rect 19518 35086 19570 35138
rect 19570 35086 19572 35138
rect 19516 35084 19572 35086
rect 19180 34354 19236 34356
rect 19180 34302 19182 34354
rect 19182 34302 19234 34354
rect 19234 34302 19236 34354
rect 19180 34300 19236 34302
rect 18508 34076 18564 34132
rect 18732 34076 18788 34132
rect 18060 31836 18116 31892
rect 18172 31666 18228 31668
rect 18172 31614 18174 31666
rect 18174 31614 18226 31666
rect 18226 31614 18228 31666
rect 18172 31612 18228 31614
rect 18060 31500 18116 31556
rect 17948 30716 18004 30772
rect 18172 31388 18228 31444
rect 17836 30268 17892 30324
rect 17500 30044 17556 30100
rect 17388 29820 17444 29876
rect 18396 30828 18452 30884
rect 18732 32060 18788 32116
rect 18396 30604 18452 30660
rect 17948 29538 18004 29540
rect 17948 29486 17950 29538
rect 17950 29486 18002 29538
rect 18002 29486 18004 29538
rect 17948 29484 18004 29486
rect 17612 29372 17668 29428
rect 17164 27916 17220 27972
rect 17276 27692 17332 27748
rect 16828 26908 16884 26964
rect 16940 27580 16996 27636
rect 16268 25116 16324 25172
rect 17052 26850 17108 26852
rect 17052 26798 17054 26850
rect 17054 26798 17106 26850
rect 17106 26798 17108 26850
rect 17052 26796 17108 26798
rect 17052 25788 17108 25844
rect 17052 25452 17108 25508
rect 16828 25116 16884 25172
rect 16828 24946 16884 24948
rect 16828 24894 16830 24946
rect 16830 24894 16882 24946
rect 16882 24894 16884 24946
rect 16828 24892 16884 24894
rect 16380 23772 16436 23828
rect 16604 23436 16660 23492
rect 16604 22540 16660 22596
rect 16716 21756 16772 21812
rect 16604 21644 16660 21700
rect 16492 21532 16548 21588
rect 16492 21362 16548 21364
rect 16492 21310 16494 21362
rect 16494 21310 16546 21362
rect 16546 21310 16548 21362
rect 16492 21308 16548 21310
rect 16716 21532 16772 21588
rect 16380 19234 16436 19236
rect 16380 19182 16382 19234
rect 16382 19182 16434 19234
rect 16434 19182 16436 19234
rect 16380 19180 16436 19182
rect 17836 29426 17892 29428
rect 17836 29374 17838 29426
rect 17838 29374 17890 29426
rect 17890 29374 17892 29426
rect 17836 29372 17892 29374
rect 18396 29372 18452 29428
rect 18508 30380 18564 30436
rect 18172 28812 18228 28868
rect 18060 28754 18116 28756
rect 18060 28702 18062 28754
rect 18062 28702 18114 28754
rect 18114 28702 18116 28754
rect 18060 28700 18116 28702
rect 18060 28364 18116 28420
rect 17948 28252 18004 28308
rect 17388 27020 17444 27076
rect 17276 26012 17332 26068
rect 17724 27970 17780 27972
rect 17724 27918 17726 27970
rect 17726 27918 17778 27970
rect 17778 27918 17780 27970
rect 17724 27916 17780 27918
rect 17500 26348 17556 26404
rect 17724 27132 17780 27188
rect 18396 28812 18452 28868
rect 18732 30994 18788 30996
rect 18732 30942 18734 30994
rect 18734 30942 18786 30994
rect 18786 30942 18788 30994
rect 18732 30940 18788 30942
rect 19180 33852 19236 33908
rect 18620 28700 18676 28756
rect 18396 28642 18452 28644
rect 18396 28590 18398 28642
rect 18398 28590 18450 28642
rect 18450 28590 18452 28642
rect 18396 28588 18452 28590
rect 19068 33292 19124 33348
rect 18844 30098 18900 30100
rect 18844 30046 18846 30098
rect 18846 30046 18898 30098
rect 18898 30046 18900 30098
rect 18844 30044 18900 30046
rect 20748 36428 20804 36484
rect 20636 36258 20692 36260
rect 20636 36206 20638 36258
rect 20638 36206 20690 36258
rect 20690 36206 20692 36258
rect 20636 36204 20692 36206
rect 20300 35644 20356 35700
rect 20636 35586 20692 35588
rect 20636 35534 20638 35586
rect 20638 35534 20690 35586
rect 20690 35534 20692 35586
rect 20636 35532 20692 35534
rect 21532 37938 21588 37940
rect 21532 37886 21534 37938
rect 21534 37886 21586 37938
rect 21586 37886 21588 37938
rect 21532 37884 21588 37886
rect 21308 36652 21364 36708
rect 21756 36652 21812 36708
rect 21532 36482 21588 36484
rect 21532 36430 21534 36482
rect 21534 36430 21586 36482
rect 21586 36430 21588 36482
rect 21532 36428 21588 36430
rect 21084 35698 21140 35700
rect 21084 35646 21086 35698
rect 21086 35646 21138 35698
rect 21138 35646 21140 35698
rect 21084 35644 21140 35646
rect 20076 34860 20132 34916
rect 19964 34802 20020 34804
rect 19964 34750 19966 34802
rect 19966 34750 20018 34802
rect 20018 34750 20020 34802
rect 19964 34748 20020 34750
rect 20188 34748 20244 34804
rect 19852 34636 19908 34692
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19740 34130 19796 34132
rect 19740 34078 19742 34130
rect 19742 34078 19794 34130
rect 19794 34078 19796 34130
rect 19740 34076 19796 34078
rect 19404 32396 19460 32452
rect 19292 31500 19348 31556
rect 20188 33852 20244 33908
rect 20636 34690 20692 34692
rect 20636 34638 20638 34690
rect 20638 34638 20690 34690
rect 20690 34638 20692 34690
rect 20636 34636 20692 34638
rect 20748 33516 20804 33572
rect 21420 34860 21476 34916
rect 21532 33628 21588 33684
rect 20524 33404 20580 33460
rect 20300 33292 20356 33348
rect 19516 31724 19572 31780
rect 19516 31388 19572 31444
rect 20412 33122 20468 33124
rect 20412 33070 20414 33122
rect 20414 33070 20466 33122
rect 20466 33070 20468 33122
rect 20412 33068 20468 33070
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 20524 32844 20580 32900
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20300 31388 20356 31444
rect 20044 31332 20100 31334
rect 20636 32060 20692 32116
rect 20636 31554 20692 31556
rect 20636 31502 20638 31554
rect 20638 31502 20690 31554
rect 20690 31502 20692 31554
rect 20636 31500 20692 31502
rect 20748 31388 20804 31444
rect 19740 30940 19796 30996
rect 20076 30882 20132 30884
rect 20076 30830 20078 30882
rect 20078 30830 20130 30882
rect 20130 30830 20132 30882
rect 20076 30828 20132 30830
rect 19852 30322 19908 30324
rect 19852 30270 19854 30322
rect 19854 30270 19906 30322
rect 19906 30270 19908 30322
rect 19852 30268 19908 30270
rect 21196 31778 21252 31780
rect 21196 31726 21198 31778
rect 21198 31726 21250 31778
rect 21250 31726 21252 31778
rect 21196 31724 21252 31726
rect 21420 31666 21476 31668
rect 21420 31614 21422 31666
rect 21422 31614 21474 31666
rect 21474 31614 21476 31666
rect 21420 31612 21476 31614
rect 20300 30322 20356 30324
rect 20300 30270 20302 30322
rect 20302 30270 20354 30322
rect 20354 30270 20356 30322
rect 20300 30268 20356 30270
rect 18732 29820 18788 29876
rect 18956 29426 19012 29428
rect 18956 29374 18958 29426
rect 18958 29374 19010 29426
rect 19010 29374 19012 29426
rect 18956 29372 19012 29374
rect 19068 28812 19124 28868
rect 18732 28364 18788 28420
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19852 29260 19908 29316
rect 19180 28252 19236 28308
rect 19292 29148 19348 29204
rect 19068 28140 19124 28196
rect 19068 27916 19124 27972
rect 18620 27858 18676 27860
rect 18620 27806 18622 27858
rect 18622 27806 18674 27858
rect 18674 27806 18676 27858
rect 18620 27804 18676 27806
rect 18844 27804 18900 27860
rect 18508 27692 18564 27748
rect 18172 27132 18228 27188
rect 18508 27020 18564 27076
rect 18844 27020 18900 27076
rect 17836 26012 17892 26068
rect 18396 26460 18452 26516
rect 17836 25116 17892 25172
rect 17500 24722 17556 24724
rect 17500 24670 17502 24722
rect 17502 24670 17554 24722
rect 17554 24670 17556 24722
rect 17500 24668 17556 24670
rect 17164 23996 17220 24052
rect 17612 23772 17668 23828
rect 17388 21868 17444 21924
rect 18284 25282 18340 25284
rect 18284 25230 18286 25282
rect 18286 25230 18338 25282
rect 18338 25230 18340 25282
rect 18284 25228 18340 25230
rect 18284 25004 18340 25060
rect 17948 24780 18004 24836
rect 18284 24834 18340 24836
rect 18284 24782 18286 24834
rect 18286 24782 18338 24834
rect 18338 24782 18340 24834
rect 18284 24780 18340 24782
rect 18172 24556 18228 24612
rect 17500 21810 17556 21812
rect 17500 21758 17502 21810
rect 17502 21758 17554 21810
rect 17554 21758 17556 21810
rect 17500 21756 17556 21758
rect 16940 21196 16996 21252
rect 16940 20636 16996 20692
rect 16828 19740 16884 19796
rect 17500 20412 17556 20468
rect 17388 19516 17444 19572
rect 17500 19404 17556 19460
rect 17164 19346 17220 19348
rect 17164 19294 17166 19346
rect 17166 19294 17218 19346
rect 17218 19294 17220 19346
rect 17164 19292 17220 19294
rect 16492 19010 16548 19012
rect 16492 18958 16494 19010
rect 16494 18958 16546 19010
rect 16546 18958 16548 19010
rect 16492 18956 16548 18958
rect 16156 17724 16212 17780
rect 17052 19180 17108 19236
rect 16716 17500 16772 17556
rect 16044 16940 16100 16996
rect 16156 16828 16212 16884
rect 15820 15314 15876 15316
rect 15820 15262 15822 15314
rect 15822 15262 15874 15314
rect 15874 15262 15876 15314
rect 15820 15260 15876 15262
rect 15932 15148 15988 15204
rect 15708 13916 15764 13972
rect 15260 11452 15316 11508
rect 15372 12236 15428 12292
rect 15708 12236 15764 12292
rect 14812 9714 14868 9716
rect 14812 9662 14814 9714
rect 14814 9662 14866 9714
rect 14866 9662 14868 9714
rect 14812 9660 14868 9662
rect 15148 9660 15204 9716
rect 15260 10610 15316 10612
rect 15260 10558 15262 10610
rect 15262 10558 15314 10610
rect 15314 10558 15316 10610
rect 15260 10556 15316 10558
rect 14700 9212 14756 9268
rect 15596 10556 15652 10612
rect 15932 12348 15988 12404
rect 15932 9996 15988 10052
rect 14700 9042 14756 9044
rect 14700 8990 14702 9042
rect 14702 8990 14754 9042
rect 14754 8990 14756 9042
rect 14700 8988 14756 8990
rect 14924 8540 14980 8596
rect 14812 8428 14868 8484
rect 15260 9042 15316 9044
rect 15260 8990 15262 9042
rect 15262 8990 15314 9042
rect 15314 8990 15316 9042
rect 15260 8988 15316 8990
rect 15036 8204 15092 8260
rect 13468 6466 13524 6468
rect 13468 6414 13470 6466
rect 13470 6414 13522 6466
rect 13522 6414 13524 6466
rect 13468 6412 13524 6414
rect 14140 6636 14196 6692
rect 13692 6188 13748 6244
rect 13916 6412 13972 6468
rect 13468 6130 13524 6132
rect 13468 6078 13470 6130
rect 13470 6078 13522 6130
rect 13522 6078 13524 6130
rect 13468 6076 13524 6078
rect 13132 5964 13188 6020
rect 13692 6018 13748 6020
rect 13692 5966 13694 6018
rect 13694 5966 13746 6018
rect 13746 5966 13748 6018
rect 13692 5964 13748 5966
rect 14588 6300 14644 6356
rect 14364 6188 14420 6244
rect 14140 5906 14196 5908
rect 14140 5854 14142 5906
rect 14142 5854 14194 5906
rect 14194 5854 14196 5906
rect 14140 5852 14196 5854
rect 14476 6130 14532 6132
rect 14476 6078 14478 6130
rect 14478 6078 14530 6130
rect 14530 6078 14532 6130
rect 14476 6076 14532 6078
rect 14364 5516 14420 5572
rect 14028 5180 14084 5236
rect 13580 5122 13636 5124
rect 13580 5070 13582 5122
rect 13582 5070 13634 5122
rect 13634 5070 13636 5122
rect 13580 5068 13636 5070
rect 13804 5010 13860 5012
rect 13804 4958 13806 5010
rect 13806 4958 13858 5010
rect 13858 4958 13860 5010
rect 13804 4956 13860 4958
rect 13020 4396 13076 4452
rect 13244 4844 13300 4900
rect 10892 3442 10948 3444
rect 10892 3390 10894 3442
rect 10894 3390 10946 3442
rect 10946 3390 10948 3442
rect 10892 3388 10948 3390
rect 11788 3442 11844 3444
rect 11788 3390 11790 3442
rect 11790 3390 11842 3442
rect 11842 3390 11844 3442
rect 11788 3388 11844 3390
rect 12684 3442 12740 3444
rect 12684 3390 12686 3442
rect 12686 3390 12738 3442
rect 12738 3390 12740 3442
rect 12684 3388 12740 3390
rect 13580 4508 13636 4564
rect 14252 5404 14308 5460
rect 14364 5292 14420 5348
rect 14252 4898 14308 4900
rect 14252 4846 14254 4898
rect 14254 4846 14306 4898
rect 14306 4846 14308 4898
rect 14252 4844 14308 4846
rect 14140 4172 14196 4228
rect 13580 3612 13636 3668
rect 14700 5906 14756 5908
rect 14700 5854 14702 5906
rect 14702 5854 14754 5906
rect 14754 5854 14756 5906
rect 14700 5852 14756 5854
rect 14924 6188 14980 6244
rect 14924 5292 14980 5348
rect 15148 8428 15204 8484
rect 14924 4620 14980 4676
rect 15036 4508 15092 4564
rect 15148 3836 15204 3892
rect 12796 1596 12852 1652
rect 15260 5068 15316 5124
rect 15708 9826 15764 9828
rect 15708 9774 15710 9826
rect 15710 9774 15762 9826
rect 15762 9774 15764 9826
rect 15708 9772 15764 9774
rect 16044 9884 16100 9940
rect 15596 8146 15652 8148
rect 15596 8094 15598 8146
rect 15598 8094 15650 8146
rect 15650 8094 15652 8146
rect 15596 8092 15652 8094
rect 15484 5906 15540 5908
rect 15484 5854 15486 5906
rect 15486 5854 15538 5906
rect 15538 5854 15540 5906
rect 15484 5852 15540 5854
rect 15932 7980 15988 8036
rect 16492 16322 16548 16324
rect 16492 16270 16494 16322
rect 16494 16270 16546 16322
rect 16546 16270 16548 16322
rect 16492 16268 16548 16270
rect 16604 16156 16660 16212
rect 16716 15932 16772 15988
rect 16268 15538 16324 15540
rect 16268 15486 16270 15538
rect 16270 15486 16322 15538
rect 16322 15486 16324 15538
rect 16268 15484 16324 15486
rect 16492 15148 16548 15204
rect 16492 14754 16548 14756
rect 16492 14702 16494 14754
rect 16494 14702 16546 14754
rect 16546 14702 16548 14754
rect 16492 14700 16548 14702
rect 16604 14530 16660 14532
rect 16604 14478 16606 14530
rect 16606 14478 16658 14530
rect 16658 14478 16660 14530
rect 16604 14476 16660 14478
rect 16492 14306 16548 14308
rect 16492 14254 16494 14306
rect 16494 14254 16546 14306
rect 16546 14254 16548 14306
rect 16492 14252 16548 14254
rect 16268 13858 16324 13860
rect 16268 13806 16270 13858
rect 16270 13806 16322 13858
rect 16322 13806 16324 13858
rect 16268 13804 16324 13806
rect 16604 14140 16660 14196
rect 16492 13692 16548 13748
rect 17052 15596 17108 15652
rect 17052 15260 17108 15316
rect 17388 18620 17444 18676
rect 17388 18396 17444 18452
rect 17388 18172 17444 18228
rect 17388 17948 17444 18004
rect 17276 17052 17332 17108
rect 17836 21308 17892 21364
rect 17948 21756 18004 21812
rect 17948 21196 18004 21252
rect 19180 27132 19236 27188
rect 19068 26572 19124 26628
rect 19180 26012 19236 26068
rect 18620 25004 18676 25060
rect 18620 23772 18676 23828
rect 18844 24780 18900 24836
rect 18956 24498 19012 24500
rect 18956 24446 18958 24498
rect 18958 24446 19010 24498
rect 19010 24446 19012 24498
rect 18956 24444 19012 24446
rect 19068 23996 19124 24052
rect 18844 22876 18900 22932
rect 18732 22482 18788 22484
rect 18732 22430 18734 22482
rect 18734 22430 18786 22482
rect 18786 22430 18788 22482
rect 18732 22428 18788 22430
rect 19180 23436 19236 23492
rect 19068 22988 19124 23044
rect 19516 29036 19572 29092
rect 19404 28530 19460 28532
rect 19404 28478 19406 28530
rect 19406 28478 19458 28530
rect 19458 28478 19460 28530
rect 19404 28476 19460 28478
rect 20300 29148 20356 29204
rect 20412 29484 20468 29540
rect 20188 29036 20244 29092
rect 19964 28754 20020 28756
rect 19964 28702 19966 28754
rect 19966 28702 20018 28754
rect 20018 28702 20020 28754
rect 19964 28700 20020 28702
rect 20076 28476 20132 28532
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19404 26460 19460 26516
rect 20076 27074 20132 27076
rect 20076 27022 20078 27074
rect 20078 27022 20130 27074
rect 20130 27022 20132 27074
rect 20076 27020 20132 27022
rect 21532 30716 21588 30772
rect 21644 32450 21700 32452
rect 21644 32398 21646 32450
rect 21646 32398 21698 32450
rect 21698 32398 21700 32450
rect 21644 32396 21700 32398
rect 21644 30604 21700 30660
rect 21980 34860 22036 34916
rect 22316 40962 22372 40964
rect 22316 40910 22318 40962
rect 22318 40910 22370 40962
rect 22370 40910 22372 40962
rect 22316 40908 22372 40910
rect 22204 39788 22260 39844
rect 22316 39618 22372 39620
rect 22316 39566 22318 39618
rect 22318 39566 22370 39618
rect 22370 39566 22372 39618
rect 22316 39564 22372 39566
rect 22428 39452 22484 39508
rect 22204 38780 22260 38836
rect 22428 38946 22484 38948
rect 22428 38894 22430 38946
rect 22430 38894 22482 38946
rect 22482 38894 22484 38946
rect 22428 38892 22484 38894
rect 22316 38668 22372 38724
rect 25228 44044 25284 44100
rect 25116 43650 25172 43652
rect 25116 43598 25118 43650
rect 25118 43598 25170 43650
rect 25170 43598 25172 43650
rect 25116 43596 25172 43598
rect 26348 45106 26404 45108
rect 26348 45054 26350 45106
rect 26350 45054 26402 45106
rect 26402 45054 26404 45106
rect 26348 45052 26404 45054
rect 27468 45052 27524 45108
rect 26124 44994 26180 44996
rect 26124 44942 26126 44994
rect 26126 44942 26178 44994
rect 26178 44942 26180 44994
rect 26124 44940 26180 44942
rect 26908 44322 26964 44324
rect 26908 44270 26910 44322
rect 26910 44270 26962 44322
rect 26962 44270 26964 44322
rect 26908 44268 26964 44270
rect 27132 44156 27188 44212
rect 25676 43650 25732 43652
rect 25676 43598 25678 43650
rect 25678 43598 25730 43650
rect 25730 43598 25732 43650
rect 25676 43596 25732 43598
rect 24668 43484 24724 43540
rect 25452 43538 25508 43540
rect 25452 43486 25454 43538
rect 25454 43486 25506 43538
rect 25506 43486 25508 43538
rect 25452 43484 25508 43486
rect 28364 44322 28420 44324
rect 28364 44270 28366 44322
rect 28366 44270 28418 44322
rect 28418 44270 28420 44322
rect 28364 44268 28420 44270
rect 27468 43820 27524 43876
rect 26572 43650 26628 43652
rect 26572 43598 26574 43650
rect 26574 43598 26626 43650
rect 26626 43598 26628 43650
rect 26572 43596 26628 43598
rect 28252 44210 28308 44212
rect 28252 44158 28254 44210
rect 28254 44158 28306 44210
rect 28306 44158 28308 44210
rect 28252 44156 28308 44158
rect 28028 44098 28084 44100
rect 28028 44046 28030 44098
rect 28030 44046 28082 44098
rect 28082 44046 28084 44098
rect 28028 44044 28084 44046
rect 28364 43820 28420 43876
rect 23996 41244 24052 41300
rect 23884 41074 23940 41076
rect 23884 41022 23886 41074
rect 23886 41022 23938 41074
rect 23938 41022 23940 41074
rect 23884 41020 23940 41022
rect 25340 42642 25396 42644
rect 25340 42590 25342 42642
rect 25342 42590 25394 42642
rect 25394 42590 25396 42642
rect 25340 42588 25396 42590
rect 26684 42700 26740 42756
rect 27916 42754 27972 42756
rect 27916 42702 27918 42754
rect 27918 42702 27970 42754
rect 27970 42702 27972 42754
rect 27916 42700 27972 42702
rect 28252 43708 28308 43764
rect 25788 42642 25844 42644
rect 25788 42590 25790 42642
rect 25790 42590 25842 42642
rect 25842 42590 25844 42642
rect 25788 42588 25844 42590
rect 26124 42642 26180 42644
rect 26124 42590 26126 42642
rect 26126 42590 26178 42642
rect 26178 42590 26180 42642
rect 26124 42588 26180 42590
rect 26796 42642 26852 42644
rect 26796 42590 26798 42642
rect 26798 42590 26850 42642
rect 26850 42590 26852 42642
rect 26796 42588 26852 42590
rect 24332 41692 24388 41748
rect 25228 42530 25284 42532
rect 25228 42478 25230 42530
rect 25230 42478 25282 42530
rect 25282 42478 25284 42530
rect 25228 42476 25284 42478
rect 26236 42252 26292 42308
rect 24668 41970 24724 41972
rect 24668 41918 24670 41970
rect 24670 41918 24722 41970
rect 24722 41918 24724 41970
rect 24668 41916 24724 41918
rect 26684 42252 26740 42308
rect 24108 40908 24164 40964
rect 23324 40572 23380 40628
rect 22988 40460 23044 40516
rect 22876 39676 22932 39732
rect 22652 39452 22708 39508
rect 22652 37826 22708 37828
rect 22652 37774 22654 37826
rect 22654 37774 22706 37826
rect 22706 37774 22708 37826
rect 22652 37772 22708 37774
rect 22204 36204 22260 36260
rect 24108 40236 24164 40292
rect 23100 39788 23156 39844
rect 22988 39564 23044 39620
rect 23212 39058 23268 39060
rect 23212 39006 23214 39058
rect 23214 39006 23266 39058
rect 23266 39006 23268 39058
rect 23212 39004 23268 39006
rect 22876 38834 22932 38836
rect 22876 38782 22878 38834
rect 22878 38782 22930 38834
rect 22930 38782 22932 38834
rect 22876 38780 22932 38782
rect 23660 38892 23716 38948
rect 24108 38722 24164 38724
rect 24108 38670 24110 38722
rect 24110 38670 24162 38722
rect 24162 38670 24164 38722
rect 24108 38668 24164 38670
rect 22988 38556 23044 38612
rect 24220 38108 24276 38164
rect 25564 41580 25620 41636
rect 24892 40962 24948 40964
rect 24892 40910 24894 40962
rect 24894 40910 24946 40962
rect 24946 40910 24948 40962
rect 24892 40908 24948 40910
rect 25788 40962 25844 40964
rect 25788 40910 25790 40962
rect 25790 40910 25842 40962
rect 25842 40910 25844 40962
rect 25788 40908 25844 40910
rect 25340 40626 25396 40628
rect 25340 40574 25342 40626
rect 25342 40574 25394 40626
rect 25394 40574 25396 40626
rect 25340 40572 25396 40574
rect 24780 40236 24836 40292
rect 25116 40236 25172 40292
rect 23548 38050 23604 38052
rect 23548 37998 23550 38050
rect 23550 37998 23602 38050
rect 23602 37998 23604 38050
rect 23548 37996 23604 37998
rect 22764 36652 22820 36708
rect 22764 36482 22820 36484
rect 22764 36430 22766 36482
rect 22766 36430 22818 36482
rect 22818 36430 22820 36482
rect 22764 36428 22820 36430
rect 22428 35868 22484 35924
rect 22652 36204 22708 36260
rect 22316 34972 22372 35028
rect 22204 34748 22260 34804
rect 24332 38050 24388 38052
rect 24332 37998 24334 38050
rect 24334 37998 24386 38050
rect 24386 37998 24388 38050
rect 24332 37996 24388 37998
rect 23884 37772 23940 37828
rect 23772 37548 23828 37604
rect 23772 36594 23828 36596
rect 23772 36542 23774 36594
rect 23774 36542 23826 36594
rect 23826 36542 23828 36594
rect 23772 36540 23828 36542
rect 23100 35980 23156 36036
rect 23660 35922 23716 35924
rect 23660 35870 23662 35922
rect 23662 35870 23714 35922
rect 23714 35870 23716 35922
rect 23660 35868 23716 35870
rect 23212 35698 23268 35700
rect 23212 35646 23214 35698
rect 23214 35646 23266 35698
rect 23266 35646 23268 35698
rect 23212 35644 23268 35646
rect 21980 33740 22036 33796
rect 21868 30492 21924 30548
rect 21308 30210 21364 30212
rect 21308 30158 21310 30210
rect 21310 30158 21362 30210
rect 21362 30158 21364 30210
rect 21308 30156 21364 30158
rect 20636 29820 20692 29876
rect 20860 29932 20916 29988
rect 22092 32508 22148 32564
rect 23548 34748 23604 34804
rect 23100 34636 23156 34692
rect 22876 33404 22932 33460
rect 23324 34076 23380 34132
rect 22428 32562 22484 32564
rect 22428 32510 22430 32562
rect 22430 32510 22482 32562
rect 22482 32510 22484 32562
rect 22428 32508 22484 32510
rect 21532 29932 21588 29988
rect 21308 29820 21364 29876
rect 20748 29372 20804 29428
rect 20636 29260 20692 29316
rect 21196 29036 21252 29092
rect 20524 28418 20580 28420
rect 20524 28366 20526 28418
rect 20526 28366 20578 28418
rect 20578 28366 20580 28418
rect 20524 28364 20580 28366
rect 20524 28140 20580 28196
rect 20636 27746 20692 27748
rect 20636 27694 20638 27746
rect 20638 27694 20690 27746
rect 20690 27694 20692 27746
rect 20636 27692 20692 27694
rect 20636 27468 20692 27524
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19516 26402 19572 26404
rect 19516 26350 19518 26402
rect 19518 26350 19570 26402
rect 19570 26350 19572 26402
rect 19516 26348 19572 26350
rect 19404 25900 19460 25956
rect 19628 25788 19684 25844
rect 19516 25676 19572 25732
rect 19516 25452 19572 25508
rect 19292 22876 19348 22932
rect 19404 25228 19460 25284
rect 18956 22316 19012 22372
rect 19068 22764 19124 22820
rect 20076 26066 20132 26068
rect 20076 26014 20078 26066
rect 20078 26014 20130 26066
rect 20130 26014 20132 26066
rect 20076 26012 20132 26014
rect 19740 25452 19796 25508
rect 19964 25228 20020 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20300 25116 20356 25172
rect 20076 24668 20132 24724
rect 19740 23938 19796 23940
rect 19740 23886 19742 23938
rect 19742 23886 19794 23938
rect 19794 23886 19796 23938
rect 19740 23884 19796 23886
rect 20188 23660 20244 23716
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 20076 23324 20132 23380
rect 19404 22764 19460 22820
rect 19516 22540 19572 22596
rect 19628 22428 19684 22484
rect 20524 26290 20580 26292
rect 20524 26238 20526 26290
rect 20526 26238 20578 26290
rect 20578 26238 20580 26290
rect 20524 26236 20580 26238
rect 20860 27692 20916 27748
rect 21084 28364 21140 28420
rect 21084 27468 21140 27524
rect 21196 27692 21252 27748
rect 21196 27020 21252 27076
rect 20748 25564 20804 25620
rect 20860 26796 20916 26852
rect 21084 26124 21140 26180
rect 20860 25340 20916 25396
rect 20636 25228 20692 25284
rect 20748 25116 20804 25172
rect 20412 23324 20468 23380
rect 20524 23884 20580 23940
rect 20076 22764 20132 22820
rect 20076 22370 20132 22372
rect 20076 22318 20078 22370
rect 20078 22318 20130 22370
rect 20130 22318 20132 22370
rect 20076 22316 20132 22318
rect 18732 21810 18788 21812
rect 18732 21758 18734 21810
rect 18734 21758 18786 21810
rect 18786 21758 18788 21810
rect 18732 21756 18788 21758
rect 17724 20300 17780 20356
rect 17724 19404 17780 19460
rect 17612 18732 17668 18788
rect 18284 20748 18340 20804
rect 18172 19852 18228 19908
rect 18172 19516 18228 19572
rect 18396 20300 18452 20356
rect 18508 20860 18564 20916
rect 18620 20524 18676 20580
rect 18956 21196 19012 21252
rect 19068 20860 19124 20916
rect 19292 21868 19348 21924
rect 19404 21698 19460 21700
rect 19404 21646 19406 21698
rect 19406 21646 19458 21698
rect 19458 21646 19460 21698
rect 19404 21644 19460 21646
rect 19292 20860 19348 20916
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20412 22652 20468 22708
rect 20188 21644 20244 21700
rect 20636 23772 20692 23828
rect 19740 21586 19796 21588
rect 19740 21534 19742 21586
rect 19742 21534 19794 21586
rect 19794 21534 19796 21586
rect 19740 21532 19796 21534
rect 20076 21586 20132 21588
rect 20076 21534 20078 21586
rect 20078 21534 20130 21586
rect 20130 21534 20132 21586
rect 20076 21532 20132 21534
rect 19628 21084 19684 21140
rect 18956 20802 19012 20804
rect 18956 20750 18958 20802
rect 18958 20750 19010 20802
rect 19010 20750 19012 20802
rect 18956 20748 19012 20750
rect 19068 20690 19124 20692
rect 19068 20638 19070 20690
rect 19070 20638 19122 20690
rect 19122 20638 19124 20690
rect 19068 20636 19124 20638
rect 19292 20636 19348 20692
rect 18396 19404 18452 19460
rect 17948 18508 18004 18564
rect 18620 19628 18676 19684
rect 19404 20412 19460 20468
rect 19180 20130 19236 20132
rect 19180 20078 19182 20130
rect 19182 20078 19234 20130
rect 19234 20078 19236 20130
rect 19180 20076 19236 20078
rect 19292 19964 19348 20020
rect 19068 19852 19124 19908
rect 19292 19628 19348 19684
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20188 20188 20244 20244
rect 20524 21698 20580 21700
rect 20524 21646 20526 21698
rect 20526 21646 20578 21698
rect 20578 21646 20580 21698
rect 20524 21644 20580 21646
rect 20412 20972 20468 21028
rect 18508 19180 18564 19236
rect 18060 18620 18116 18676
rect 17612 18284 17668 18340
rect 18060 18226 18116 18228
rect 18060 18174 18062 18226
rect 18062 18174 18114 18226
rect 18114 18174 18116 18226
rect 18060 18172 18116 18174
rect 18284 18844 18340 18900
rect 18508 18956 18564 19012
rect 18172 17612 18228 17668
rect 17500 17052 17556 17108
rect 17948 17052 18004 17108
rect 17500 16770 17556 16772
rect 17500 16718 17502 16770
rect 17502 16718 17554 16770
rect 17554 16718 17556 16770
rect 17500 16716 17556 16718
rect 16940 13916 16996 13972
rect 17500 16380 17556 16436
rect 16716 13356 16772 13412
rect 16380 13020 16436 13076
rect 16268 12402 16324 12404
rect 16268 12350 16270 12402
rect 16270 12350 16322 12402
rect 16322 12350 16324 12402
rect 16268 12348 16324 12350
rect 16828 12572 16884 12628
rect 16940 13132 16996 13188
rect 16380 12290 16436 12292
rect 16380 12238 16382 12290
rect 16382 12238 16434 12290
rect 16434 12238 16436 12290
rect 16380 12236 16436 12238
rect 16716 12460 16772 12516
rect 17276 13804 17332 13860
rect 17612 15986 17668 15988
rect 17612 15934 17614 15986
rect 17614 15934 17666 15986
rect 17666 15934 17668 15986
rect 17612 15932 17668 15934
rect 17500 15538 17556 15540
rect 17500 15486 17502 15538
rect 17502 15486 17554 15538
rect 17554 15486 17556 15538
rect 17500 15484 17556 15486
rect 18060 16882 18116 16884
rect 18060 16830 18062 16882
rect 18062 16830 18114 16882
rect 18114 16830 18116 16882
rect 18060 16828 18116 16830
rect 18284 17052 18340 17108
rect 18396 18284 18452 18340
rect 19852 19516 19908 19572
rect 20188 20018 20244 20020
rect 20188 19966 20190 20018
rect 20190 19966 20242 20018
rect 20242 19966 20244 20018
rect 20188 19964 20244 19966
rect 19740 19404 19796 19460
rect 19740 19234 19796 19236
rect 19740 19182 19742 19234
rect 19742 19182 19794 19234
rect 19794 19182 19796 19234
rect 19740 19180 19796 19182
rect 20860 23884 20916 23940
rect 21084 25228 21140 25284
rect 20636 19964 20692 20020
rect 20748 20524 20804 20580
rect 20748 20076 20804 20132
rect 20524 19346 20580 19348
rect 20524 19294 20526 19346
rect 20526 19294 20578 19346
rect 20578 19294 20580 19346
rect 20524 19292 20580 19294
rect 20076 18956 20132 19012
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 20524 18844 20580 18900
rect 19404 18338 19460 18340
rect 19404 18286 19406 18338
rect 19406 18286 19458 18338
rect 19458 18286 19460 18338
rect 19404 18284 19460 18286
rect 18620 17106 18676 17108
rect 18620 17054 18622 17106
rect 18622 17054 18674 17106
rect 18674 17054 18676 17106
rect 18620 17052 18676 17054
rect 18284 15596 18340 15652
rect 17948 15036 18004 15092
rect 17724 14364 17780 14420
rect 17500 13804 17556 13860
rect 17164 12850 17220 12852
rect 17164 12798 17166 12850
rect 17166 12798 17218 12850
rect 17218 12798 17220 12850
rect 17164 12796 17220 12798
rect 17724 13692 17780 13748
rect 17164 12012 17220 12068
rect 16492 11676 16548 11732
rect 16940 11788 16996 11844
rect 16268 10834 16324 10836
rect 16268 10782 16270 10834
rect 16270 10782 16322 10834
rect 16322 10782 16324 10834
rect 16268 10780 16324 10782
rect 16380 10610 16436 10612
rect 16380 10558 16382 10610
rect 16382 10558 16434 10610
rect 16434 10558 16436 10610
rect 16380 10556 16436 10558
rect 16828 11282 16884 11284
rect 16828 11230 16830 11282
rect 16830 11230 16882 11282
rect 16882 11230 16884 11282
rect 16828 11228 16884 11230
rect 16380 9938 16436 9940
rect 16380 9886 16382 9938
rect 16382 9886 16434 9938
rect 16434 9886 16436 9938
rect 16380 9884 16436 9886
rect 16268 9772 16324 9828
rect 15820 7586 15876 7588
rect 15820 7534 15822 7586
rect 15822 7534 15874 7586
rect 15874 7534 15876 7586
rect 15820 7532 15876 7534
rect 16268 7308 16324 7364
rect 17164 11282 17220 11284
rect 17164 11230 17166 11282
rect 17166 11230 17218 11282
rect 17218 11230 17220 11282
rect 17164 11228 17220 11230
rect 17948 13468 18004 13524
rect 18844 17164 18900 17220
rect 19740 18338 19796 18340
rect 19740 18286 19742 18338
rect 19742 18286 19794 18338
rect 19794 18286 19796 18338
rect 19740 18284 19796 18286
rect 19068 17052 19124 17108
rect 18732 16268 18788 16324
rect 20300 18450 20356 18452
rect 20300 18398 20302 18450
rect 20302 18398 20354 18450
rect 20354 18398 20356 18450
rect 20300 18396 20356 18398
rect 19852 17836 19908 17892
rect 19628 17666 19684 17668
rect 19628 17614 19630 17666
rect 19630 17614 19682 17666
rect 19682 17614 19684 17666
rect 19628 17612 19684 17614
rect 19516 17388 19572 17444
rect 20076 17442 20132 17444
rect 20076 17390 20078 17442
rect 20078 17390 20130 17442
rect 20130 17390 20132 17442
rect 20076 17388 20132 17390
rect 19628 17164 19684 17220
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20076 16940 20132 16996
rect 19740 15874 19796 15876
rect 19740 15822 19742 15874
rect 19742 15822 19794 15874
rect 19794 15822 19796 15874
rect 19740 15820 19796 15822
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19068 15484 19124 15540
rect 19404 15314 19460 15316
rect 19404 15262 19406 15314
rect 19406 15262 19458 15314
rect 19458 15262 19460 15314
rect 19404 15260 19460 15262
rect 18508 14476 18564 14532
rect 19628 14812 19684 14868
rect 18620 14418 18676 14420
rect 18620 14366 18622 14418
rect 18622 14366 18674 14418
rect 18674 14366 18676 14418
rect 18620 14364 18676 14366
rect 20300 14252 20356 14308
rect 19628 14140 19684 14196
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20636 17890 20692 17892
rect 20636 17838 20638 17890
rect 20638 17838 20690 17890
rect 20690 17838 20692 17890
rect 20636 17836 20692 17838
rect 20636 17442 20692 17444
rect 20636 17390 20638 17442
rect 20638 17390 20690 17442
rect 20690 17390 20692 17442
rect 20636 17388 20692 17390
rect 20636 16940 20692 16996
rect 20524 15932 20580 15988
rect 20412 14028 20468 14084
rect 19740 13916 19796 13972
rect 18060 13244 18116 13300
rect 18060 12908 18116 12964
rect 19180 13132 19236 13188
rect 18508 13020 18564 13076
rect 18732 13020 18788 13076
rect 18172 12572 18228 12628
rect 18620 12684 18676 12740
rect 17612 11900 17668 11956
rect 17276 10780 17332 10836
rect 18508 12402 18564 12404
rect 18508 12350 18510 12402
rect 18510 12350 18562 12402
rect 18562 12350 18564 12402
rect 18508 12348 18564 12350
rect 18620 12124 18676 12180
rect 18508 11900 18564 11956
rect 17948 11452 18004 11508
rect 18060 11788 18116 11844
rect 17724 10834 17780 10836
rect 17724 10782 17726 10834
rect 17726 10782 17778 10834
rect 17778 10782 17780 10834
rect 17724 10780 17780 10782
rect 18396 11788 18452 11844
rect 18396 11564 18452 11620
rect 18284 11452 18340 11508
rect 17836 10610 17892 10612
rect 17836 10558 17838 10610
rect 17838 10558 17890 10610
rect 17890 10558 17892 10610
rect 17836 10556 17892 10558
rect 19068 12124 19124 12180
rect 18956 11900 19012 11956
rect 18620 10892 18676 10948
rect 17724 9772 17780 9828
rect 16828 9212 16884 9268
rect 16828 8146 16884 8148
rect 16828 8094 16830 8146
rect 16830 8094 16882 8146
rect 16882 8094 16884 8146
rect 16828 8092 16884 8094
rect 17052 8146 17108 8148
rect 17052 8094 17054 8146
rect 17054 8094 17106 8146
rect 17106 8094 17108 8146
rect 17052 8092 17108 8094
rect 16940 8034 16996 8036
rect 16940 7982 16942 8034
rect 16942 7982 16994 8034
rect 16994 7982 16996 8034
rect 16940 7980 16996 7982
rect 16940 7698 16996 7700
rect 16940 7646 16942 7698
rect 16942 7646 16994 7698
rect 16994 7646 16996 7698
rect 16940 7644 16996 7646
rect 16716 7420 16772 7476
rect 17276 7474 17332 7476
rect 17276 7422 17278 7474
rect 17278 7422 17330 7474
rect 17330 7422 17332 7474
rect 17276 7420 17332 7422
rect 17500 7532 17556 7588
rect 16716 6860 16772 6916
rect 16380 6636 16436 6692
rect 16716 6524 16772 6580
rect 16828 6130 16884 6132
rect 16828 6078 16830 6130
rect 16830 6078 16882 6130
rect 16882 6078 16884 6130
rect 16828 6076 16884 6078
rect 15484 5122 15540 5124
rect 15484 5070 15486 5122
rect 15486 5070 15538 5122
rect 15538 5070 15540 5122
rect 15484 5068 15540 5070
rect 16604 5180 16660 5236
rect 17500 7362 17556 7364
rect 17500 7310 17502 7362
rect 17502 7310 17554 7362
rect 17554 7310 17556 7362
rect 17500 7308 17556 7310
rect 17500 6636 17556 6692
rect 17052 5068 17108 5124
rect 15596 4732 15652 4788
rect 16044 4956 16100 5012
rect 16492 4732 16548 4788
rect 17724 9548 17780 9604
rect 18172 9548 18228 9604
rect 18284 9266 18340 9268
rect 18284 9214 18286 9266
rect 18286 9214 18338 9266
rect 18338 9214 18340 9266
rect 18284 9212 18340 9214
rect 18956 10722 19012 10724
rect 18956 10670 18958 10722
rect 18958 10670 19010 10722
rect 19010 10670 19012 10722
rect 18956 10668 19012 10670
rect 18732 9884 18788 9940
rect 18620 9772 18676 9828
rect 18620 8428 18676 8484
rect 17836 8034 17892 8036
rect 17836 7982 17838 8034
rect 17838 7982 17890 8034
rect 17890 7982 17892 8034
rect 17836 7980 17892 7982
rect 17724 6972 17780 7028
rect 18508 7980 18564 8036
rect 18620 7756 18676 7812
rect 18620 7532 18676 7588
rect 18172 7420 18228 7476
rect 17724 6466 17780 6468
rect 17724 6414 17726 6466
rect 17726 6414 17778 6466
rect 17778 6414 17780 6466
rect 17724 6412 17780 6414
rect 17500 6130 17556 6132
rect 17500 6078 17502 6130
rect 17502 6078 17554 6130
rect 17554 6078 17556 6130
rect 17500 6076 17556 6078
rect 17612 5906 17668 5908
rect 17612 5854 17614 5906
rect 17614 5854 17666 5906
rect 17666 5854 17668 5906
rect 17612 5852 17668 5854
rect 17724 5740 17780 5796
rect 17276 4732 17332 4788
rect 17724 3666 17780 3668
rect 17724 3614 17726 3666
rect 17726 3614 17778 3666
rect 17778 3614 17780 3666
rect 17724 3612 17780 3614
rect 15260 3388 15316 3444
rect 10780 1372 10836 1428
rect 17948 6076 18004 6132
rect 18060 6636 18116 6692
rect 18508 7362 18564 7364
rect 18508 7310 18510 7362
rect 18510 7310 18562 7362
rect 18562 7310 18564 7362
rect 18508 7308 18564 7310
rect 18284 6972 18340 7028
rect 18844 8146 18900 8148
rect 18844 8094 18846 8146
rect 18846 8094 18898 8146
rect 18898 8094 18900 8146
rect 18844 8092 18900 8094
rect 18844 7698 18900 7700
rect 18844 7646 18846 7698
rect 18846 7646 18898 7698
rect 18898 7646 18900 7698
rect 18844 7644 18900 7646
rect 18844 7084 18900 7140
rect 18284 5740 18340 5796
rect 18060 4172 18116 4228
rect 18172 5180 18228 5236
rect 18620 6412 18676 6468
rect 18620 5964 18676 6020
rect 18396 4956 18452 5012
rect 18508 5516 18564 5572
rect 18284 4226 18340 4228
rect 18284 4174 18286 4226
rect 18286 4174 18338 4226
rect 18338 4174 18340 4226
rect 18284 4172 18340 4174
rect 18844 6578 18900 6580
rect 18844 6526 18846 6578
rect 18846 6526 18898 6578
rect 18898 6526 18900 6578
rect 18844 6524 18900 6526
rect 19180 10610 19236 10612
rect 19180 10558 19182 10610
rect 19182 10558 19234 10610
rect 19234 10558 19236 10610
rect 19180 10556 19236 10558
rect 21756 29314 21812 29316
rect 21756 29262 21758 29314
rect 21758 29262 21810 29314
rect 21810 29262 21812 29314
rect 21756 29260 21812 29262
rect 21420 29148 21476 29204
rect 21644 28812 21700 28868
rect 21420 27970 21476 27972
rect 21420 27918 21422 27970
rect 21422 27918 21474 27970
rect 21474 27918 21476 27970
rect 21420 27916 21476 27918
rect 22316 31276 22372 31332
rect 23660 34242 23716 34244
rect 23660 34190 23662 34242
rect 23662 34190 23714 34242
rect 23714 34190 23716 34242
rect 23660 34188 23716 34190
rect 23436 33628 23492 33684
rect 23436 33404 23492 33460
rect 23436 32732 23492 32788
rect 22988 31948 23044 32004
rect 22540 31500 22596 31556
rect 22652 31836 22708 31892
rect 22428 31106 22484 31108
rect 22428 31054 22430 31106
rect 22430 31054 22482 31106
rect 22482 31054 22484 31106
rect 22428 31052 22484 31054
rect 22876 31276 22932 31332
rect 23100 31890 23156 31892
rect 23100 31838 23102 31890
rect 23102 31838 23154 31890
rect 23154 31838 23156 31890
rect 23100 31836 23156 31838
rect 23324 32284 23380 32340
rect 22988 31052 23044 31108
rect 22652 30268 22708 30324
rect 22316 30156 22372 30212
rect 22764 28700 22820 28756
rect 22204 28364 22260 28420
rect 22428 28364 22484 28420
rect 22428 27692 22484 27748
rect 22540 28140 22596 28196
rect 22204 27356 22260 27412
rect 22092 27074 22148 27076
rect 22092 27022 22094 27074
rect 22094 27022 22146 27074
rect 22146 27022 22148 27074
rect 22092 27020 22148 27022
rect 21532 26850 21588 26852
rect 21532 26798 21534 26850
rect 21534 26798 21586 26850
rect 21586 26798 21588 26850
rect 21532 26796 21588 26798
rect 21420 26178 21476 26180
rect 21420 26126 21422 26178
rect 21422 26126 21474 26178
rect 21474 26126 21476 26178
rect 21420 26124 21476 26126
rect 21532 25676 21588 25732
rect 22092 26124 22148 26180
rect 21868 25618 21924 25620
rect 21868 25566 21870 25618
rect 21870 25566 21922 25618
rect 21922 25566 21924 25618
rect 21868 25564 21924 25566
rect 21756 25228 21812 25284
rect 21420 23938 21476 23940
rect 21420 23886 21422 23938
rect 21422 23886 21474 23938
rect 21474 23886 21476 23938
rect 21420 23884 21476 23886
rect 21196 21698 21252 21700
rect 21196 21646 21198 21698
rect 21198 21646 21250 21698
rect 21250 21646 21252 21698
rect 21196 21644 21252 21646
rect 20860 19628 20916 19684
rect 20860 18732 20916 18788
rect 21420 21756 21476 21812
rect 21420 21196 21476 21252
rect 23996 36482 24052 36484
rect 23996 36430 23998 36482
rect 23998 36430 24050 36482
rect 24050 36430 24052 36482
rect 23996 36428 24052 36430
rect 24892 39506 24948 39508
rect 24892 39454 24894 39506
rect 24894 39454 24946 39506
rect 24946 39454 24948 39506
rect 24892 39452 24948 39454
rect 25004 39004 25060 39060
rect 24668 38780 24724 38836
rect 24668 38556 24724 38612
rect 25228 38610 25284 38612
rect 25228 38558 25230 38610
rect 25230 38558 25282 38610
rect 25282 38558 25284 38610
rect 25228 38556 25284 38558
rect 25564 40626 25620 40628
rect 25564 40574 25566 40626
rect 25566 40574 25618 40626
rect 25618 40574 25620 40626
rect 25564 40572 25620 40574
rect 27916 41804 27972 41860
rect 25788 40514 25844 40516
rect 25788 40462 25790 40514
rect 25790 40462 25842 40514
rect 25842 40462 25844 40514
rect 25788 40460 25844 40462
rect 26124 39676 26180 39732
rect 27468 40626 27524 40628
rect 27468 40574 27470 40626
rect 27470 40574 27522 40626
rect 27522 40574 27524 40626
rect 27468 40572 27524 40574
rect 27804 40572 27860 40628
rect 26796 39506 26852 39508
rect 26796 39454 26798 39506
rect 26798 39454 26850 39506
rect 26850 39454 26852 39506
rect 26796 39452 26852 39454
rect 25452 38556 25508 38612
rect 26012 38556 26068 38612
rect 25676 38444 25732 38500
rect 27356 39730 27412 39732
rect 27356 39678 27358 39730
rect 27358 39678 27410 39730
rect 27410 39678 27412 39730
rect 27356 39676 27412 39678
rect 27916 40402 27972 40404
rect 27916 40350 27918 40402
rect 27918 40350 27970 40402
rect 27970 40350 27972 40402
rect 27916 40348 27972 40350
rect 28252 39842 28308 39844
rect 28252 39790 28254 39842
rect 28254 39790 28306 39842
rect 28306 39790 28308 39842
rect 28252 39788 28308 39790
rect 27804 38834 27860 38836
rect 27804 38782 27806 38834
rect 27806 38782 27858 38834
rect 27858 38782 27860 38834
rect 27804 38780 27860 38782
rect 27132 38556 27188 38612
rect 26348 37884 26404 37940
rect 27020 38108 27076 38164
rect 25228 36876 25284 36932
rect 25900 36652 25956 36708
rect 23996 35698 24052 35700
rect 23996 35646 23998 35698
rect 23998 35646 24050 35698
rect 24050 35646 24052 35698
rect 23996 35644 24052 35646
rect 23884 34524 23940 34580
rect 23996 34412 24052 34468
rect 24108 34860 24164 34916
rect 24108 34300 24164 34356
rect 23212 29932 23268 29988
rect 23548 30210 23604 30212
rect 23548 30158 23550 30210
rect 23550 30158 23602 30210
rect 23602 30158 23604 30210
rect 23548 30156 23604 30158
rect 23436 29708 23492 29764
rect 24108 32786 24164 32788
rect 24108 32734 24110 32786
rect 24110 32734 24162 32786
rect 24162 32734 24164 32786
rect 24108 32732 24164 32734
rect 24108 31778 24164 31780
rect 24108 31726 24110 31778
rect 24110 31726 24162 31778
rect 24162 31726 24164 31778
rect 24108 31724 24164 31726
rect 23996 31612 24052 31668
rect 23996 31164 24052 31220
rect 23772 30492 23828 30548
rect 23996 30716 24052 30772
rect 23772 30268 23828 30324
rect 24108 30604 24164 30660
rect 24332 35026 24388 35028
rect 24332 34974 24334 35026
rect 24334 34974 24386 35026
rect 24386 34974 24388 35026
rect 24332 34972 24388 34974
rect 24332 34188 24388 34244
rect 24668 35084 24724 35140
rect 24556 34130 24612 34132
rect 24556 34078 24558 34130
rect 24558 34078 24610 34130
rect 24610 34078 24612 34130
rect 24556 34076 24612 34078
rect 24668 33628 24724 33684
rect 25004 35644 25060 35700
rect 24444 33234 24500 33236
rect 24444 33182 24446 33234
rect 24446 33182 24498 33234
rect 24498 33182 24500 33234
rect 24444 33180 24500 33182
rect 24444 32844 24500 32900
rect 24444 30716 24500 30772
rect 24892 32172 24948 32228
rect 24780 31836 24836 31892
rect 24220 29932 24276 29988
rect 23100 29036 23156 29092
rect 23436 29148 23492 29204
rect 23100 27020 23156 27076
rect 23212 27804 23268 27860
rect 22316 26290 22372 26292
rect 22316 26238 22318 26290
rect 22318 26238 22370 26290
rect 22370 26238 22372 26290
rect 22316 26236 22372 26238
rect 22204 24892 22260 24948
rect 22876 26796 22932 26852
rect 22764 25788 22820 25844
rect 23324 26348 23380 26404
rect 22540 24220 22596 24276
rect 22764 25228 22820 25284
rect 22092 22204 22148 22260
rect 22764 24668 22820 24724
rect 21868 21756 21924 21812
rect 21532 20802 21588 20804
rect 21532 20750 21534 20802
rect 21534 20750 21586 20802
rect 21586 20750 21588 20802
rect 21532 20748 21588 20750
rect 21756 20914 21812 20916
rect 21756 20862 21758 20914
rect 21758 20862 21810 20914
rect 21810 20862 21812 20914
rect 21756 20860 21812 20862
rect 21644 20076 21700 20132
rect 21532 19740 21588 19796
rect 21420 19628 21476 19684
rect 21868 19180 21924 19236
rect 21756 19122 21812 19124
rect 21756 19070 21758 19122
rect 21758 19070 21810 19122
rect 21810 19070 21812 19122
rect 21756 19068 21812 19070
rect 21644 18956 21700 19012
rect 21532 18284 21588 18340
rect 20748 15932 20804 15988
rect 20748 15484 20804 15540
rect 20860 15260 20916 15316
rect 20748 14642 20804 14644
rect 20748 14590 20750 14642
rect 20750 14590 20802 14642
rect 20802 14590 20804 14642
rect 20748 14588 20804 14590
rect 20748 13916 20804 13972
rect 20412 12908 20468 12964
rect 19836 12570 19892 12572
rect 19628 12460 19684 12516
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19964 12402 20020 12404
rect 19964 12350 19966 12402
rect 19966 12350 20018 12402
rect 20018 12350 20020 12402
rect 19964 12348 20020 12350
rect 19628 11900 19684 11956
rect 19404 9772 19460 9828
rect 19516 10892 19572 10948
rect 20300 11564 20356 11620
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 21420 16380 21476 16436
rect 20972 15036 21028 15092
rect 20860 13468 20916 13524
rect 20748 13074 20804 13076
rect 20748 13022 20750 13074
rect 20750 13022 20802 13074
rect 20802 13022 20804 13074
rect 20748 13020 20804 13022
rect 20636 11452 20692 11508
rect 20748 12572 20804 12628
rect 20972 12178 21028 12180
rect 20972 12126 20974 12178
rect 20974 12126 21026 12178
rect 21026 12126 21028 12178
rect 20972 12124 21028 12126
rect 20412 10834 20468 10836
rect 20412 10782 20414 10834
rect 20414 10782 20466 10834
rect 20466 10782 20468 10834
rect 20412 10780 20468 10782
rect 19852 9996 19908 10052
rect 19404 9324 19460 9380
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19292 8930 19348 8932
rect 19292 8878 19294 8930
rect 19294 8878 19346 8930
rect 19346 8878 19348 8930
rect 19292 8876 19348 8878
rect 19180 8370 19236 8372
rect 19180 8318 19182 8370
rect 19182 8318 19234 8370
rect 19234 8318 19236 8370
rect 19180 8316 19236 8318
rect 19292 7698 19348 7700
rect 19292 7646 19294 7698
rect 19294 7646 19346 7698
rect 19346 7646 19348 7698
rect 19292 7644 19348 7646
rect 19068 7532 19124 7588
rect 20300 9212 20356 9268
rect 19516 8876 19572 8932
rect 19852 8316 19908 8372
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19964 7250 20020 7252
rect 19964 7198 19966 7250
rect 19966 7198 20018 7250
rect 20018 7198 20020 7250
rect 19964 7196 20020 7198
rect 19852 7084 19908 7140
rect 19516 6690 19572 6692
rect 19516 6638 19518 6690
rect 19518 6638 19570 6690
rect 19570 6638 19572 6690
rect 19516 6636 19572 6638
rect 19292 6130 19348 6132
rect 19292 6078 19294 6130
rect 19294 6078 19346 6130
rect 19346 6078 19348 6130
rect 19292 6076 19348 6078
rect 18956 5740 19012 5796
rect 19180 5292 19236 5348
rect 19292 4732 19348 4788
rect 18844 3666 18900 3668
rect 18844 3614 18846 3666
rect 18846 3614 18898 3666
rect 18898 3614 18900 3666
rect 18844 3612 18900 3614
rect 20748 10892 20804 10948
rect 20860 11788 20916 11844
rect 20748 10722 20804 10724
rect 20748 10670 20750 10722
rect 20750 10670 20802 10722
rect 20802 10670 20804 10722
rect 20748 10668 20804 10670
rect 20748 9714 20804 9716
rect 20748 9662 20750 9714
rect 20750 9662 20802 9714
rect 20802 9662 20804 9714
rect 20748 9660 20804 9662
rect 20636 9100 20692 9156
rect 21420 15708 21476 15764
rect 21196 14476 21252 14532
rect 21868 18508 21924 18564
rect 22204 21196 22260 21252
rect 22316 21084 22372 21140
rect 22092 20636 22148 20692
rect 22204 19852 22260 19908
rect 21980 17836 22036 17892
rect 22092 19234 22148 19236
rect 22092 19182 22094 19234
rect 22094 19182 22146 19234
rect 22146 19182 22148 19234
rect 22092 19180 22148 19182
rect 22092 18508 22148 18564
rect 22876 23266 22932 23268
rect 22876 23214 22878 23266
rect 22878 23214 22930 23266
rect 22930 23214 22932 23266
rect 22876 23212 22932 23214
rect 22764 21868 22820 21924
rect 23772 27132 23828 27188
rect 23772 26178 23828 26180
rect 23772 26126 23774 26178
rect 23774 26126 23826 26178
rect 23826 26126 23828 26178
rect 23772 26124 23828 26126
rect 23548 25788 23604 25844
rect 23436 25228 23492 25284
rect 23772 25228 23828 25284
rect 23548 24722 23604 24724
rect 23548 24670 23550 24722
rect 23550 24670 23602 24722
rect 23602 24670 23604 24722
rect 23548 24668 23604 24670
rect 23100 23938 23156 23940
rect 23100 23886 23102 23938
rect 23102 23886 23154 23938
rect 23154 23886 23156 23938
rect 23100 23884 23156 23886
rect 23436 23826 23492 23828
rect 23436 23774 23438 23826
rect 23438 23774 23490 23826
rect 23490 23774 23492 23826
rect 23436 23772 23492 23774
rect 23212 23378 23268 23380
rect 23212 23326 23214 23378
rect 23214 23326 23266 23378
rect 23266 23326 23268 23378
rect 23212 23324 23268 23326
rect 22988 22540 23044 22596
rect 22540 21586 22596 21588
rect 22540 21534 22542 21586
rect 22542 21534 22594 21586
rect 22594 21534 22596 21586
rect 22540 21532 22596 21534
rect 22764 21420 22820 21476
rect 22540 19628 22596 19684
rect 22428 19010 22484 19012
rect 22428 18958 22430 19010
rect 22430 18958 22482 19010
rect 22482 18958 22484 19010
rect 22428 18956 22484 18958
rect 22540 18060 22596 18116
rect 22428 17106 22484 17108
rect 22428 17054 22430 17106
rect 22430 17054 22482 17106
rect 22482 17054 22484 17106
rect 22428 17052 22484 17054
rect 22764 19180 22820 19236
rect 22764 18844 22820 18900
rect 22764 18172 22820 18228
rect 22764 17612 22820 17668
rect 22764 17052 22820 17108
rect 22540 16882 22596 16884
rect 22540 16830 22542 16882
rect 22542 16830 22594 16882
rect 22594 16830 22596 16882
rect 22540 16828 22596 16830
rect 23324 21308 23380 21364
rect 23212 20748 23268 20804
rect 23100 19628 23156 19684
rect 23660 23324 23716 23380
rect 24108 29708 24164 29764
rect 24220 28812 24276 28868
rect 23996 28700 24052 28756
rect 24108 28642 24164 28644
rect 24108 28590 24110 28642
rect 24110 28590 24162 28642
rect 24162 28590 24164 28642
rect 24108 28588 24164 28590
rect 24108 27970 24164 27972
rect 24108 27918 24110 27970
rect 24110 27918 24162 27970
rect 24162 27918 24164 27970
rect 24108 27916 24164 27918
rect 24668 29036 24724 29092
rect 24444 27858 24500 27860
rect 24444 27806 24446 27858
rect 24446 27806 24498 27858
rect 24498 27806 24500 27858
rect 24444 27804 24500 27806
rect 24220 27692 24276 27748
rect 23996 27244 24052 27300
rect 24332 26514 24388 26516
rect 24332 26462 24334 26514
rect 24334 26462 24386 26514
rect 24386 26462 24388 26514
rect 24332 26460 24388 26462
rect 25900 35868 25956 35924
rect 25116 34748 25172 34804
rect 25340 34130 25396 34132
rect 25340 34078 25342 34130
rect 25342 34078 25394 34130
rect 25394 34078 25396 34130
rect 25340 34076 25396 34078
rect 25452 33180 25508 33236
rect 25452 32956 25508 33012
rect 25228 31500 25284 31556
rect 25452 32732 25508 32788
rect 25676 32172 25732 32228
rect 25564 31836 25620 31892
rect 25564 31388 25620 31444
rect 25340 30882 25396 30884
rect 25340 30830 25342 30882
rect 25342 30830 25394 30882
rect 25394 30830 25396 30882
rect 25340 30828 25396 30830
rect 25340 30604 25396 30660
rect 25116 27186 25172 27188
rect 25116 27134 25118 27186
rect 25118 27134 25170 27186
rect 25170 27134 25172 27186
rect 25116 27132 25172 27134
rect 25004 25900 25060 25956
rect 23772 23212 23828 23268
rect 23772 23042 23828 23044
rect 23772 22990 23774 23042
rect 23774 22990 23826 23042
rect 23826 22990 23828 23042
rect 23772 22988 23828 22990
rect 23772 22092 23828 22148
rect 23660 21698 23716 21700
rect 23660 21646 23662 21698
rect 23662 21646 23714 21698
rect 23714 21646 23716 21698
rect 23660 21644 23716 21646
rect 23548 21532 23604 21588
rect 24108 23324 24164 23380
rect 24556 23324 24612 23380
rect 24332 23212 24388 23268
rect 25340 28700 25396 28756
rect 25340 28252 25396 28308
rect 25340 27804 25396 27860
rect 25340 27074 25396 27076
rect 25340 27022 25342 27074
rect 25342 27022 25394 27074
rect 25394 27022 25396 27074
rect 25340 27020 25396 27022
rect 26124 37212 26180 37268
rect 26348 36876 26404 36932
rect 26572 36482 26628 36484
rect 26572 36430 26574 36482
rect 26574 36430 26626 36482
rect 26626 36430 26628 36482
rect 26572 36428 26628 36430
rect 26796 36652 26852 36708
rect 28140 39506 28196 39508
rect 28140 39454 28142 39506
rect 28142 39454 28194 39506
rect 28194 39454 28196 39506
rect 28140 39452 28196 39454
rect 29932 44940 29988 44996
rect 29260 43708 29316 43764
rect 30492 44268 30548 44324
rect 28700 43148 28756 43204
rect 28476 40572 28532 40628
rect 28588 39340 28644 39396
rect 28364 38668 28420 38724
rect 27916 38108 27972 38164
rect 27580 37938 27636 37940
rect 27580 37886 27582 37938
rect 27582 37886 27634 37938
rect 27634 37886 27636 37938
rect 27580 37884 27636 37886
rect 28252 37324 28308 37380
rect 28476 37660 28532 37716
rect 27580 36706 27636 36708
rect 27580 36654 27582 36706
rect 27582 36654 27634 36706
rect 27634 36654 27636 36706
rect 27580 36652 27636 36654
rect 27020 36370 27076 36372
rect 27020 36318 27022 36370
rect 27022 36318 27074 36370
rect 27074 36318 27076 36370
rect 27020 36316 27076 36318
rect 26796 36204 26852 36260
rect 26460 35868 26516 35924
rect 26796 35586 26852 35588
rect 26796 35534 26798 35586
rect 26798 35534 26850 35586
rect 26850 35534 26852 35586
rect 26796 35532 26852 35534
rect 26572 33964 26628 34020
rect 26236 33628 26292 33684
rect 26348 33068 26404 33124
rect 26012 32956 26068 33012
rect 26684 32732 26740 32788
rect 27356 36482 27412 36484
rect 27356 36430 27358 36482
rect 27358 36430 27410 36482
rect 27410 36430 27412 36482
rect 27356 36428 27412 36430
rect 27692 35810 27748 35812
rect 27692 35758 27694 35810
rect 27694 35758 27746 35810
rect 27746 35758 27748 35810
rect 27692 35756 27748 35758
rect 27468 35532 27524 35588
rect 28588 36258 28644 36260
rect 28588 36206 28590 36258
rect 28590 36206 28642 36258
rect 28642 36206 28644 36258
rect 28588 36204 28644 36206
rect 28588 35698 28644 35700
rect 28588 35646 28590 35698
rect 28590 35646 28642 35698
rect 28642 35646 28644 35698
rect 28588 35644 28644 35646
rect 27244 34972 27300 35028
rect 27580 34914 27636 34916
rect 27580 34862 27582 34914
rect 27582 34862 27634 34914
rect 27634 34862 27636 34914
rect 27580 34860 27636 34862
rect 27356 34748 27412 34804
rect 27468 33516 27524 33572
rect 26684 32284 26740 32340
rect 26460 31778 26516 31780
rect 26460 31726 26462 31778
rect 26462 31726 26514 31778
rect 26514 31726 26516 31778
rect 26460 31724 26516 31726
rect 27020 32284 27076 32340
rect 26796 31724 26852 31780
rect 27132 31778 27188 31780
rect 27132 31726 27134 31778
rect 27134 31726 27186 31778
rect 27186 31726 27188 31778
rect 27132 31724 27188 31726
rect 26012 30716 26068 30772
rect 25900 30380 25956 30436
rect 25676 29260 25732 29316
rect 27132 29372 27188 29428
rect 26572 29314 26628 29316
rect 26572 29262 26574 29314
rect 26574 29262 26626 29314
rect 26626 29262 26628 29314
rect 26572 29260 26628 29262
rect 28812 41858 28868 41860
rect 28812 41806 28814 41858
rect 28814 41806 28866 41858
rect 28866 41806 28868 41858
rect 28812 41804 28868 41806
rect 29260 42866 29316 42868
rect 29260 42814 29262 42866
rect 29262 42814 29314 42866
rect 29314 42814 29316 42866
rect 29260 42812 29316 42814
rect 29036 41692 29092 41748
rect 29148 42476 29204 42532
rect 29484 42700 29540 42756
rect 29484 42530 29540 42532
rect 29484 42478 29486 42530
rect 29486 42478 29538 42530
rect 29538 42478 29540 42530
rect 29484 42476 29540 42478
rect 30268 44210 30324 44212
rect 30268 44158 30270 44210
rect 30270 44158 30322 44210
rect 30322 44158 30324 44210
rect 30268 44156 30324 44158
rect 31388 44994 31444 44996
rect 31388 44942 31390 44994
rect 31390 44942 31442 44994
rect 31442 44942 31444 44994
rect 31388 44940 31444 44942
rect 33404 46060 33460 46116
rect 31836 44492 31892 44548
rect 30828 43932 30884 43988
rect 29708 43538 29764 43540
rect 29708 43486 29710 43538
rect 29710 43486 29762 43538
rect 29762 43486 29764 43538
rect 29708 43484 29764 43486
rect 30044 42866 30100 42868
rect 30044 42814 30046 42866
rect 30046 42814 30098 42866
rect 30098 42814 30100 42866
rect 30044 42812 30100 42814
rect 30044 42252 30100 42308
rect 29260 41916 29316 41972
rect 29260 41356 29316 41412
rect 29148 41020 29204 41076
rect 29036 39788 29092 39844
rect 29932 41692 29988 41748
rect 31052 43708 31108 43764
rect 30940 43650 30996 43652
rect 30940 43598 30942 43650
rect 30942 43598 30994 43650
rect 30994 43598 30996 43650
rect 30940 43596 30996 43598
rect 31164 43538 31220 43540
rect 31164 43486 31166 43538
rect 31166 43486 31218 43538
rect 31218 43486 31220 43538
rect 31164 43484 31220 43486
rect 30828 43036 30884 43092
rect 30268 42476 30324 42532
rect 30716 42028 30772 42084
rect 30156 41410 30212 41412
rect 30156 41358 30158 41410
rect 30158 41358 30210 41410
rect 30210 41358 30212 41410
rect 30156 41356 30212 41358
rect 30604 41692 30660 41748
rect 29596 40684 29652 40740
rect 30268 40236 30324 40292
rect 30156 39900 30212 39956
rect 29372 39676 29428 39732
rect 29036 39452 29092 39508
rect 30156 39618 30212 39620
rect 30156 39566 30158 39618
rect 30158 39566 30210 39618
rect 30210 39566 30212 39618
rect 30156 39564 30212 39566
rect 29484 39340 29540 39396
rect 29148 38946 29204 38948
rect 29148 38894 29150 38946
rect 29150 38894 29202 38946
rect 29202 38894 29204 38946
rect 29148 38892 29204 38894
rect 30044 38892 30100 38948
rect 29260 37660 29316 37716
rect 29596 37772 29652 37828
rect 29708 38108 29764 38164
rect 29484 37548 29540 37604
rect 29260 37378 29316 37380
rect 29260 37326 29262 37378
rect 29262 37326 29314 37378
rect 29314 37326 29316 37378
rect 29260 37324 29316 37326
rect 28924 36540 28980 36596
rect 29148 36370 29204 36372
rect 29148 36318 29150 36370
rect 29150 36318 29202 36370
rect 29202 36318 29204 36370
rect 29148 36316 29204 36318
rect 29260 35756 29316 35812
rect 29148 35644 29204 35700
rect 29372 35644 29428 35700
rect 30940 42924 30996 42980
rect 30828 37996 30884 38052
rect 30268 37660 30324 37716
rect 30828 37772 30884 37828
rect 30044 37548 30100 37604
rect 30044 37266 30100 37268
rect 30044 37214 30046 37266
rect 30046 37214 30098 37266
rect 30098 37214 30100 37266
rect 30044 37212 30100 37214
rect 31276 42754 31332 42756
rect 31276 42702 31278 42754
rect 31278 42702 31330 42754
rect 31330 42702 31332 42754
rect 31276 42700 31332 42702
rect 31500 42028 31556 42084
rect 31164 41858 31220 41860
rect 31164 41806 31166 41858
rect 31166 41806 31218 41858
rect 31218 41806 31220 41858
rect 31164 41804 31220 41806
rect 31836 42252 31892 42308
rect 32172 44940 32228 44996
rect 32284 44156 32340 44212
rect 32060 43596 32116 43652
rect 32060 43036 32116 43092
rect 32172 42700 32228 42756
rect 31948 41074 32004 41076
rect 31948 41022 31950 41074
rect 31950 41022 32002 41074
rect 32002 41022 32004 41074
rect 31948 41020 32004 41022
rect 31948 40796 32004 40852
rect 31388 40236 31444 40292
rect 31836 40236 31892 40292
rect 31164 39618 31220 39620
rect 31164 39566 31166 39618
rect 31166 39566 31218 39618
rect 31218 39566 31220 39618
rect 31164 39564 31220 39566
rect 31948 39564 32004 39620
rect 31276 38946 31332 38948
rect 31276 38894 31278 38946
rect 31278 38894 31330 38946
rect 31330 38894 31332 38946
rect 31276 38892 31332 38894
rect 31836 38668 31892 38724
rect 31388 37660 31444 37716
rect 31500 37548 31556 37604
rect 31052 37436 31108 37492
rect 29148 34412 29204 34468
rect 30044 35868 30100 35924
rect 30156 34972 30212 35028
rect 30492 35644 30548 35700
rect 32060 39676 32116 39732
rect 32172 39506 32228 39508
rect 32172 39454 32174 39506
rect 32174 39454 32226 39506
rect 32226 39454 32228 39506
rect 32172 39452 32228 39454
rect 32844 43708 32900 43764
rect 32508 43426 32564 43428
rect 32508 43374 32510 43426
rect 32510 43374 32562 43426
rect 32562 43374 32564 43426
rect 32508 43372 32564 43374
rect 32508 41970 32564 41972
rect 32508 41918 32510 41970
rect 32510 41918 32562 41970
rect 32562 41918 32564 41970
rect 32508 41916 32564 41918
rect 32396 41132 32452 41188
rect 32508 40684 32564 40740
rect 32508 40514 32564 40516
rect 32508 40462 32510 40514
rect 32510 40462 32562 40514
rect 32562 40462 32564 40514
rect 32508 40460 32564 40462
rect 33180 44940 33236 44996
rect 33740 44546 33796 44548
rect 33740 44494 33742 44546
rect 33742 44494 33794 44546
rect 33794 44494 33796 44546
rect 33740 44492 33796 44494
rect 33964 44044 34020 44100
rect 34860 44156 34916 44212
rect 33180 42812 33236 42868
rect 33068 41692 33124 41748
rect 33068 41132 33124 41188
rect 34076 43260 34132 43316
rect 34748 43650 34804 43652
rect 34748 43598 34750 43650
rect 34750 43598 34802 43650
rect 34802 43598 34804 43650
rect 34748 43596 34804 43598
rect 33964 42812 34020 42868
rect 34076 43036 34132 43092
rect 34188 42754 34244 42756
rect 34188 42702 34190 42754
rect 34190 42702 34242 42754
rect 34242 42702 34244 42754
rect 34188 42700 34244 42702
rect 33628 42364 33684 42420
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35084 45836 35140 45892
rect 35980 45890 36036 45892
rect 35980 45838 35982 45890
rect 35982 45838 36034 45890
rect 36034 45838 36036 45890
rect 35980 45836 36036 45838
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 36428 44940 36484 44996
rect 36988 46114 37044 46116
rect 36988 46062 36990 46114
rect 36990 46062 37042 46114
rect 37042 46062 37044 46114
rect 36988 46060 37044 46062
rect 38108 46060 38164 46116
rect 36540 44492 36596 44548
rect 37212 44546 37268 44548
rect 37212 44494 37214 44546
rect 37214 44494 37266 44546
rect 37266 44494 37268 44546
rect 37212 44492 37268 44494
rect 35868 43596 35924 43652
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35308 42924 35364 42980
rect 35868 42924 35924 42980
rect 34748 42588 34804 42644
rect 33628 41916 33684 41972
rect 34412 41858 34468 41860
rect 34412 41806 34414 41858
rect 34414 41806 34466 41858
rect 34466 41806 34468 41858
rect 34412 41804 34468 41806
rect 36316 44156 36372 44212
rect 37548 43538 37604 43540
rect 37548 43486 37550 43538
rect 37550 43486 37602 43538
rect 37602 43486 37604 43538
rect 37548 43484 37604 43486
rect 37548 43036 37604 43092
rect 37100 42978 37156 42980
rect 37100 42926 37102 42978
rect 37102 42926 37154 42978
rect 37154 42926 37156 42978
rect 37100 42924 37156 42926
rect 37100 42642 37156 42644
rect 37100 42590 37102 42642
rect 37102 42590 37154 42642
rect 37154 42590 37156 42642
rect 37100 42588 37156 42590
rect 37212 42140 37268 42196
rect 36428 42082 36484 42084
rect 36428 42030 36430 42082
rect 36430 42030 36482 42082
rect 36482 42030 36484 42082
rect 36428 42028 36484 42030
rect 35532 41804 35588 41860
rect 33404 41580 33460 41636
rect 33740 41580 33796 41636
rect 33292 40684 33348 40740
rect 32956 40124 33012 40180
rect 33404 39900 33460 39956
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35196 41132 35252 41188
rect 34300 41074 34356 41076
rect 34300 41022 34302 41074
rect 34302 41022 34354 41074
rect 34354 41022 34356 41074
rect 34300 41020 34356 41022
rect 35196 40460 35252 40516
rect 35084 40402 35140 40404
rect 35084 40350 35086 40402
rect 35086 40350 35138 40402
rect 35138 40350 35140 40402
rect 35084 40348 35140 40350
rect 35980 41020 36036 41076
rect 36428 41020 36484 41076
rect 36316 40908 36372 40964
rect 36204 40684 36260 40740
rect 36316 40348 36372 40404
rect 33516 39676 33572 39732
rect 33964 40124 34020 40180
rect 32284 39004 32340 39060
rect 32508 38892 32564 38948
rect 32732 38668 32788 38724
rect 33740 39452 33796 39508
rect 33404 38892 33460 38948
rect 33180 38722 33236 38724
rect 33180 38670 33182 38722
rect 33182 38670 33234 38722
rect 33234 38670 33236 38722
rect 33180 38668 33236 38670
rect 31948 38444 32004 38500
rect 33852 38556 33908 38612
rect 32396 38444 32452 38500
rect 32284 37996 32340 38052
rect 31948 37212 32004 37268
rect 30940 35644 30996 35700
rect 31052 36370 31108 36372
rect 31052 36318 31054 36370
rect 31054 36318 31106 36370
rect 31106 36318 31108 36370
rect 31052 36316 31108 36318
rect 29596 34300 29652 34356
rect 30940 34748 30996 34804
rect 29708 34076 29764 34132
rect 27916 32620 27972 32676
rect 28700 32562 28756 32564
rect 28700 32510 28702 32562
rect 28702 32510 28754 32562
rect 28754 32510 28756 32562
rect 28700 32508 28756 32510
rect 27468 32172 27524 32228
rect 27580 30828 27636 30884
rect 27468 29372 27524 29428
rect 26236 28924 26292 28980
rect 26684 28642 26740 28644
rect 26684 28590 26686 28642
rect 26686 28590 26738 28642
rect 26738 28590 26740 28642
rect 26684 28588 26740 28590
rect 26908 28530 26964 28532
rect 26908 28478 26910 28530
rect 26910 28478 26962 28530
rect 26962 28478 26964 28530
rect 26908 28476 26964 28478
rect 26796 27858 26852 27860
rect 26796 27806 26798 27858
rect 26798 27806 26850 27858
rect 26850 27806 26852 27858
rect 26796 27804 26852 27806
rect 26460 27580 26516 27636
rect 25228 25116 25284 25172
rect 27132 28588 27188 28644
rect 27244 27970 27300 27972
rect 27244 27918 27246 27970
rect 27246 27918 27298 27970
rect 27298 27918 27300 27970
rect 27244 27916 27300 27918
rect 27020 27580 27076 27636
rect 27356 27132 27412 27188
rect 27692 29148 27748 29204
rect 27804 32172 27860 32228
rect 28588 31666 28644 31668
rect 28588 31614 28590 31666
rect 28590 31614 28642 31666
rect 28642 31614 28644 31666
rect 28588 31612 28644 31614
rect 31612 35586 31668 35588
rect 31612 35534 31614 35586
rect 31614 35534 31666 35586
rect 31666 35534 31668 35586
rect 31612 35532 31668 35534
rect 31276 34972 31332 35028
rect 29148 32508 29204 32564
rect 29260 33068 29316 33124
rect 29596 32674 29652 32676
rect 29596 32622 29598 32674
rect 29598 32622 29650 32674
rect 29650 32622 29652 32674
rect 29596 32620 29652 32622
rect 30716 32620 30772 32676
rect 29148 31666 29204 31668
rect 29148 31614 29150 31666
rect 29150 31614 29202 31666
rect 29202 31614 29204 31666
rect 29148 31612 29204 31614
rect 29260 31554 29316 31556
rect 29260 31502 29262 31554
rect 29262 31502 29314 31554
rect 29314 31502 29316 31554
rect 29260 31500 29316 31502
rect 28924 31276 28980 31332
rect 28252 30828 28308 30884
rect 28700 30940 28756 30996
rect 30380 31500 30436 31556
rect 30156 31164 30212 31220
rect 28700 30156 28756 30212
rect 30492 31612 30548 31668
rect 30492 31052 30548 31108
rect 31388 34914 31444 34916
rect 31388 34862 31390 34914
rect 31390 34862 31442 34914
rect 31442 34862 31444 34914
rect 31388 34860 31444 34862
rect 31276 34748 31332 34804
rect 32732 37938 32788 37940
rect 32732 37886 32734 37938
rect 32734 37886 32786 37938
rect 32786 37886 32788 37938
rect 32732 37884 32788 37886
rect 33740 37436 33796 37492
rect 32508 37266 32564 37268
rect 32508 37214 32510 37266
rect 32510 37214 32562 37266
rect 32562 37214 32564 37266
rect 32508 37212 32564 37214
rect 33516 37266 33572 37268
rect 33516 37214 33518 37266
rect 33518 37214 33570 37266
rect 33570 37214 33572 37266
rect 33516 37212 33572 37214
rect 32396 36370 32452 36372
rect 32396 36318 32398 36370
rect 32398 36318 32450 36370
rect 32450 36318 32452 36370
rect 32396 36316 32452 36318
rect 32172 35868 32228 35924
rect 32284 35810 32340 35812
rect 32284 35758 32286 35810
rect 32286 35758 32338 35810
rect 32338 35758 32340 35810
rect 32284 35756 32340 35758
rect 31948 35698 32004 35700
rect 31948 35646 31950 35698
rect 31950 35646 32002 35698
rect 32002 35646 32004 35698
rect 31948 35644 32004 35646
rect 31948 34860 32004 34916
rect 31724 34748 31780 34804
rect 32396 34748 32452 34804
rect 32956 36482 33012 36484
rect 32956 36430 32958 36482
rect 32958 36430 33010 36482
rect 33010 36430 33012 36482
rect 32956 36428 33012 36430
rect 33628 36482 33684 36484
rect 33628 36430 33630 36482
rect 33630 36430 33682 36482
rect 33682 36430 33684 36482
rect 33628 36428 33684 36430
rect 33180 36316 33236 36372
rect 33516 35868 33572 35924
rect 32732 34972 32788 35028
rect 33292 34972 33348 35028
rect 32844 34690 32900 34692
rect 32844 34638 32846 34690
rect 32846 34638 32898 34690
rect 32898 34638 32900 34690
rect 32844 34636 32900 34638
rect 33404 34802 33460 34804
rect 33404 34750 33406 34802
rect 33406 34750 33458 34802
rect 33458 34750 33460 34802
rect 33404 34748 33460 34750
rect 33516 34636 33572 34692
rect 32060 33346 32116 33348
rect 32060 33294 32062 33346
rect 32062 33294 32114 33346
rect 32114 33294 32116 33346
rect 32060 33292 32116 33294
rect 31500 33180 31556 33236
rect 31612 31164 31668 31220
rect 30828 30994 30884 30996
rect 30828 30942 30830 30994
rect 30830 30942 30882 30994
rect 30882 30942 30884 30994
rect 30828 30940 30884 30942
rect 30380 30716 30436 30772
rect 31388 30716 31444 30772
rect 31836 31164 31892 31220
rect 31836 30882 31892 30884
rect 31836 30830 31838 30882
rect 31838 30830 31890 30882
rect 31890 30830 31892 30882
rect 31836 30828 31892 30830
rect 28588 29596 28644 29652
rect 27916 29484 27972 29540
rect 28588 29372 28644 29428
rect 28140 29314 28196 29316
rect 28140 29262 28142 29314
rect 28142 29262 28194 29314
rect 28194 29262 28196 29314
rect 28140 29260 28196 29262
rect 27580 28812 27636 28868
rect 27580 27858 27636 27860
rect 27580 27806 27582 27858
rect 27582 27806 27634 27858
rect 27634 27806 27636 27858
rect 27580 27804 27636 27806
rect 26572 26684 26628 26740
rect 26908 26572 26964 26628
rect 26684 26514 26740 26516
rect 26684 26462 26686 26514
rect 26686 26462 26738 26514
rect 26738 26462 26740 26514
rect 26684 26460 26740 26462
rect 26236 26402 26292 26404
rect 26236 26350 26238 26402
rect 26238 26350 26290 26402
rect 26290 26350 26292 26402
rect 26236 26348 26292 26350
rect 25788 26178 25844 26180
rect 25788 26126 25790 26178
rect 25790 26126 25842 26178
rect 25842 26126 25844 26178
rect 25788 26124 25844 26126
rect 26572 26124 26628 26180
rect 26012 25506 26068 25508
rect 26012 25454 26014 25506
rect 26014 25454 26066 25506
rect 26066 25454 26068 25506
rect 26012 25452 26068 25454
rect 26236 25452 26292 25508
rect 25228 24722 25284 24724
rect 25228 24670 25230 24722
rect 25230 24670 25282 24722
rect 25282 24670 25284 24722
rect 25228 24668 25284 24670
rect 25900 24892 25956 24948
rect 24556 22930 24612 22932
rect 24556 22878 24558 22930
rect 24558 22878 24610 22930
rect 24610 22878 24612 22930
rect 24556 22876 24612 22878
rect 24444 22092 24500 22148
rect 24332 21868 24388 21924
rect 23884 21420 23940 21476
rect 24556 21308 24612 21364
rect 23772 20802 23828 20804
rect 23772 20750 23774 20802
rect 23774 20750 23826 20802
rect 23826 20750 23828 20802
rect 23772 20748 23828 20750
rect 24892 21868 24948 21924
rect 24220 20690 24276 20692
rect 24220 20638 24222 20690
rect 24222 20638 24274 20690
rect 24274 20638 24276 20690
rect 24220 20636 24276 20638
rect 23548 19740 23604 19796
rect 23212 19404 23268 19460
rect 23436 18732 23492 18788
rect 23660 19180 23716 19236
rect 23324 18450 23380 18452
rect 23324 18398 23326 18450
rect 23326 18398 23378 18450
rect 23378 18398 23380 18450
rect 23324 18396 23380 18398
rect 23548 18172 23604 18228
rect 23100 18060 23156 18116
rect 22988 16828 23044 16884
rect 21756 15986 21812 15988
rect 21756 15934 21758 15986
rect 21758 15934 21810 15986
rect 21810 15934 21812 15986
rect 21756 15932 21812 15934
rect 21644 14924 21700 14980
rect 22092 14588 22148 14644
rect 21196 14028 21252 14084
rect 21084 11004 21140 11060
rect 21532 13746 21588 13748
rect 21532 13694 21534 13746
rect 21534 13694 21586 13746
rect 21586 13694 21588 13746
rect 21532 13692 21588 13694
rect 22764 16156 22820 16212
rect 22428 15708 22484 15764
rect 22316 14924 22372 14980
rect 21756 14364 21812 14420
rect 22092 14028 22148 14084
rect 21420 13468 21476 13524
rect 21308 11676 21364 11732
rect 21644 13020 21700 13076
rect 21756 12850 21812 12852
rect 21756 12798 21758 12850
rect 21758 12798 21810 12850
rect 21810 12798 21812 12850
rect 21756 12796 21812 12798
rect 21644 12684 21700 12740
rect 21532 11788 21588 11844
rect 21980 11788 22036 11844
rect 23772 19068 23828 19124
rect 23884 18620 23940 18676
rect 23996 18508 24052 18564
rect 24108 19292 24164 19348
rect 23884 18172 23940 18228
rect 23436 17500 23492 17556
rect 23100 16380 23156 16436
rect 23548 16604 23604 16660
rect 23324 16268 23380 16324
rect 22092 13580 22148 13636
rect 21420 11564 21476 11620
rect 21644 11452 21700 11508
rect 21196 10892 21252 10948
rect 21084 10610 21140 10612
rect 21084 10558 21086 10610
rect 21086 10558 21138 10610
rect 21138 10558 21140 10610
rect 21084 10556 21140 10558
rect 21196 10332 21252 10388
rect 20972 10220 21028 10276
rect 20860 8652 20916 8708
rect 21084 9884 21140 9940
rect 21420 8988 21476 9044
rect 21084 8428 21140 8484
rect 21644 10108 21700 10164
rect 21868 10668 21924 10724
rect 22316 13634 22372 13636
rect 22316 13582 22318 13634
rect 22318 13582 22370 13634
rect 22370 13582 22372 13634
rect 22316 13580 22372 13582
rect 24332 19740 24388 19796
rect 24444 19628 24500 19684
rect 24780 19404 24836 19460
rect 24444 18562 24500 18564
rect 24444 18510 24446 18562
rect 24446 18510 24498 18562
rect 24498 18510 24500 18562
rect 24444 18508 24500 18510
rect 24668 18338 24724 18340
rect 24668 18286 24670 18338
rect 24670 18286 24722 18338
rect 24722 18286 24724 18338
rect 24668 18284 24724 18286
rect 25340 23548 25396 23604
rect 25340 22428 25396 22484
rect 25116 22316 25172 22372
rect 25452 22316 25508 22372
rect 25228 22258 25284 22260
rect 25228 22206 25230 22258
rect 25230 22206 25282 22258
rect 25282 22206 25284 22258
rect 25228 22204 25284 22206
rect 25228 21756 25284 21812
rect 25564 22092 25620 22148
rect 25452 21084 25508 21140
rect 25564 20860 25620 20916
rect 25340 20802 25396 20804
rect 25340 20750 25342 20802
rect 25342 20750 25394 20802
rect 25394 20750 25396 20802
rect 25340 20748 25396 20750
rect 25004 20524 25060 20580
rect 25564 20300 25620 20356
rect 25116 20188 25172 20244
rect 25452 20188 25508 20244
rect 25340 20130 25396 20132
rect 25340 20078 25342 20130
rect 25342 20078 25394 20130
rect 25394 20078 25396 20130
rect 25340 20076 25396 20078
rect 25340 19794 25396 19796
rect 25340 19742 25342 19794
rect 25342 19742 25394 19794
rect 25394 19742 25396 19794
rect 25340 19740 25396 19742
rect 25116 18620 25172 18676
rect 24220 17948 24276 18004
rect 24780 17948 24836 18004
rect 24108 17500 24164 17556
rect 24668 17666 24724 17668
rect 24668 17614 24670 17666
rect 24670 17614 24722 17666
rect 24722 17614 24724 17666
rect 24668 17612 24724 17614
rect 23772 16882 23828 16884
rect 23772 16830 23774 16882
rect 23774 16830 23826 16882
rect 23826 16830 23828 16882
rect 23772 16828 23828 16830
rect 24332 17106 24388 17108
rect 24332 17054 24334 17106
rect 24334 17054 24386 17106
rect 24386 17054 24388 17106
rect 24332 17052 24388 17054
rect 24108 16604 24164 16660
rect 23884 16210 23940 16212
rect 23884 16158 23886 16210
rect 23886 16158 23938 16210
rect 23938 16158 23940 16210
rect 23884 16156 23940 16158
rect 23772 15708 23828 15764
rect 23884 14700 23940 14756
rect 23436 14364 23492 14420
rect 23548 14028 23604 14084
rect 22540 13916 22596 13972
rect 22540 13522 22596 13524
rect 22540 13470 22542 13522
rect 22542 13470 22594 13522
rect 22594 13470 22596 13522
rect 22540 13468 22596 13470
rect 22428 12796 22484 12852
rect 23324 13916 23380 13972
rect 22876 13692 22932 13748
rect 22876 13244 22932 13300
rect 22316 11676 22372 11732
rect 23212 13746 23268 13748
rect 23212 13694 23214 13746
rect 23214 13694 23266 13746
rect 23266 13694 23268 13746
rect 23212 13692 23268 13694
rect 23660 13858 23716 13860
rect 23660 13806 23662 13858
rect 23662 13806 23714 13858
rect 23714 13806 23716 13858
rect 23660 13804 23716 13806
rect 23548 13692 23604 13748
rect 22316 11116 22372 11172
rect 21980 10332 22036 10388
rect 22092 10220 22148 10276
rect 21196 8204 21252 8260
rect 20412 8146 20468 8148
rect 20412 8094 20414 8146
rect 20414 8094 20466 8146
rect 20466 8094 20468 8146
rect 20412 8092 20468 8094
rect 21532 8316 21588 8372
rect 20300 7756 20356 7812
rect 21532 7868 21588 7924
rect 20860 7756 20916 7812
rect 20412 7250 20468 7252
rect 20412 7198 20414 7250
rect 20414 7198 20466 7250
rect 20466 7198 20468 7250
rect 20412 7196 20468 7198
rect 20188 6748 20244 6804
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19964 6076 20020 6132
rect 20636 6636 20692 6692
rect 19628 5346 19684 5348
rect 19628 5294 19630 5346
rect 19630 5294 19682 5346
rect 19682 5294 19684 5346
rect 19628 5292 19684 5294
rect 20076 5740 20132 5796
rect 19516 4508 19572 4564
rect 19628 5068 19684 5124
rect 19516 4172 19572 4228
rect 20748 6076 20804 6132
rect 20748 5180 20804 5236
rect 20412 5122 20468 5124
rect 20412 5070 20414 5122
rect 20414 5070 20466 5122
rect 20466 5070 20468 5122
rect 20412 5068 20468 5070
rect 20300 5010 20356 5012
rect 20300 4958 20302 5010
rect 20302 4958 20354 5010
rect 20354 4958 20356 5010
rect 20300 4956 20356 4958
rect 19964 4844 20020 4900
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 20076 4508 20132 4564
rect 20748 4338 20804 4340
rect 20748 4286 20750 4338
rect 20750 4286 20802 4338
rect 20802 4286 20804 4338
rect 20748 4284 20804 4286
rect 21420 7756 21476 7812
rect 21084 7586 21140 7588
rect 21084 7534 21086 7586
rect 21086 7534 21138 7586
rect 21138 7534 21140 7586
rect 21084 7532 21140 7534
rect 20972 7084 21028 7140
rect 21196 7196 21252 7252
rect 21868 8930 21924 8932
rect 21868 8878 21870 8930
rect 21870 8878 21922 8930
rect 21922 8878 21924 8930
rect 21868 8876 21924 8878
rect 23100 13132 23156 13188
rect 22652 11564 22708 11620
rect 23436 12962 23492 12964
rect 23436 12910 23438 12962
rect 23438 12910 23490 12962
rect 23490 12910 23492 12962
rect 23436 12908 23492 12910
rect 23884 14252 23940 14308
rect 24220 16098 24276 16100
rect 24220 16046 24222 16098
rect 24222 16046 24274 16098
rect 24274 16046 24276 16098
rect 24220 16044 24276 16046
rect 24332 15932 24388 15988
rect 24556 17388 24612 17444
rect 24668 17164 24724 17220
rect 24780 17052 24836 17108
rect 24780 16828 24836 16884
rect 25116 17388 25172 17444
rect 25228 16770 25284 16772
rect 25228 16718 25230 16770
rect 25230 16718 25282 16770
rect 25282 16718 25284 16770
rect 25228 16716 25284 16718
rect 24668 15708 24724 15764
rect 24332 15484 24388 15540
rect 24108 13692 24164 13748
rect 24444 15148 24500 15204
rect 23772 13356 23828 13412
rect 23660 11788 23716 11844
rect 23100 11618 23156 11620
rect 23100 11566 23102 11618
rect 23102 11566 23154 11618
rect 23154 11566 23156 11618
rect 23100 11564 23156 11566
rect 23436 11676 23492 11732
rect 23324 11340 23380 11396
rect 22988 10610 23044 10612
rect 22988 10558 22990 10610
rect 22990 10558 23042 10610
rect 23042 10558 23044 10610
rect 22988 10556 23044 10558
rect 23100 9660 23156 9716
rect 23212 10220 23268 10276
rect 22428 9548 22484 9604
rect 22092 9154 22148 9156
rect 22092 9102 22094 9154
rect 22094 9102 22146 9154
rect 22146 9102 22148 9154
rect 22092 9100 22148 9102
rect 21756 8092 21812 8148
rect 22204 9042 22260 9044
rect 22204 8990 22206 9042
rect 22206 8990 22258 9042
rect 22258 8990 22260 9042
rect 22204 8988 22260 8990
rect 21644 7644 21700 7700
rect 21196 5794 21252 5796
rect 21196 5742 21198 5794
rect 21198 5742 21250 5794
rect 21250 5742 21252 5794
rect 21196 5740 21252 5742
rect 21196 5068 21252 5124
rect 21084 4956 21140 5012
rect 21756 7532 21812 7588
rect 21980 8034 22036 8036
rect 21980 7982 21982 8034
rect 21982 7982 22034 8034
rect 22034 7982 22036 8034
rect 21980 7980 22036 7982
rect 23324 10108 23380 10164
rect 23548 11564 23604 11620
rect 23548 11116 23604 11172
rect 23548 10386 23604 10388
rect 23548 10334 23550 10386
rect 23550 10334 23602 10386
rect 23602 10334 23604 10386
rect 23548 10332 23604 10334
rect 23436 9660 23492 9716
rect 22764 8652 22820 8708
rect 22764 7308 22820 7364
rect 22204 7196 22260 7252
rect 21756 6748 21812 6804
rect 22092 6860 22148 6916
rect 22316 6636 22372 6692
rect 21756 5794 21812 5796
rect 21756 5742 21758 5794
rect 21758 5742 21810 5794
rect 21810 5742 21812 5794
rect 21756 5740 21812 5742
rect 22316 5740 22372 5796
rect 22204 5122 22260 5124
rect 22204 5070 22206 5122
rect 22206 5070 22258 5122
rect 22258 5070 22260 5122
rect 22204 5068 22260 5070
rect 22540 6018 22596 6020
rect 22540 5966 22542 6018
rect 22542 5966 22594 6018
rect 22594 5966 22596 6018
rect 22540 5964 22596 5966
rect 22540 5404 22596 5460
rect 23436 8876 23492 8932
rect 22988 8428 23044 8484
rect 23324 8764 23380 8820
rect 23100 8092 23156 8148
rect 23212 7868 23268 7924
rect 23100 6524 23156 6580
rect 22988 6130 23044 6132
rect 22988 6078 22990 6130
rect 22990 6078 23042 6130
rect 23042 6078 23044 6130
rect 22988 6076 23044 6078
rect 22988 5628 23044 5684
rect 22428 4844 22484 4900
rect 21420 4284 21476 4340
rect 21420 3666 21476 3668
rect 21420 3614 21422 3666
rect 21422 3614 21474 3666
rect 21474 3614 21476 3666
rect 21420 3612 21476 3614
rect 21868 3666 21924 3668
rect 21868 3614 21870 3666
rect 21870 3614 21922 3666
rect 21922 3614 21924 3666
rect 21868 3612 21924 3614
rect 22764 5010 22820 5012
rect 22764 4958 22766 5010
rect 22766 4958 22818 5010
rect 22818 4958 22820 5010
rect 22764 4956 22820 4958
rect 23100 4844 23156 4900
rect 23100 4172 23156 4228
rect 24108 12236 24164 12292
rect 24220 12012 24276 12068
rect 24332 13244 24388 13300
rect 23996 11564 24052 11620
rect 23884 10780 23940 10836
rect 23772 10668 23828 10724
rect 23996 10108 24052 10164
rect 23884 8204 23940 8260
rect 23324 7308 23380 7364
rect 25228 16044 25284 16100
rect 24892 15874 24948 15876
rect 24892 15822 24894 15874
rect 24894 15822 24946 15874
rect 24946 15822 24948 15874
rect 24892 15820 24948 15822
rect 26012 23266 26068 23268
rect 26012 23214 26014 23266
rect 26014 23214 26066 23266
rect 26066 23214 26068 23266
rect 26012 23212 26068 23214
rect 26012 21586 26068 21588
rect 26012 21534 26014 21586
rect 26014 21534 26066 21586
rect 26066 21534 26068 21586
rect 26012 21532 26068 21534
rect 26124 20412 26180 20468
rect 26684 25506 26740 25508
rect 26684 25454 26686 25506
rect 26686 25454 26738 25506
rect 26738 25454 26740 25506
rect 26684 25452 26740 25454
rect 26572 25340 26628 25396
rect 27244 26124 27300 26180
rect 26908 25228 26964 25284
rect 27244 25788 27300 25844
rect 26572 23266 26628 23268
rect 26572 23214 26574 23266
rect 26574 23214 26626 23266
rect 26626 23214 26628 23266
rect 26572 23212 26628 23214
rect 27132 22876 27188 22932
rect 27132 22652 27188 22708
rect 27468 26850 27524 26852
rect 27468 26798 27470 26850
rect 27470 26798 27522 26850
rect 27522 26798 27524 26850
rect 27468 26796 27524 26798
rect 27468 26348 27524 26404
rect 27580 26178 27636 26180
rect 27580 26126 27582 26178
rect 27582 26126 27634 26178
rect 27634 26126 27636 26178
rect 27580 26124 27636 26126
rect 28140 28812 28196 28868
rect 28476 28754 28532 28756
rect 28476 28702 28478 28754
rect 28478 28702 28530 28754
rect 28530 28702 28532 28754
rect 28476 28700 28532 28702
rect 29260 30044 29316 30100
rect 29148 29538 29204 29540
rect 29148 29486 29150 29538
rect 29150 29486 29202 29538
rect 29202 29486 29204 29538
rect 29148 29484 29204 29486
rect 28812 29426 28868 29428
rect 28812 29374 28814 29426
rect 28814 29374 28866 29426
rect 28866 29374 28868 29426
rect 28812 29372 28868 29374
rect 27804 28028 27860 28084
rect 28364 28418 28420 28420
rect 28364 28366 28366 28418
rect 28366 28366 28418 28418
rect 28418 28366 28420 28418
rect 28364 28364 28420 28366
rect 27804 27020 27860 27076
rect 28140 27858 28196 27860
rect 28140 27806 28142 27858
rect 28142 27806 28194 27858
rect 28194 27806 28196 27858
rect 28140 27804 28196 27806
rect 28364 27356 28420 27412
rect 28252 27074 28308 27076
rect 28252 27022 28254 27074
rect 28254 27022 28306 27074
rect 28306 27022 28308 27074
rect 28252 27020 28308 27022
rect 28028 26124 28084 26180
rect 27692 25676 27748 25732
rect 27580 25618 27636 25620
rect 27580 25566 27582 25618
rect 27582 25566 27634 25618
rect 27634 25566 27636 25618
rect 27580 25564 27636 25566
rect 27356 25340 27412 25396
rect 27580 25340 27636 25396
rect 27356 25116 27412 25172
rect 28252 25282 28308 25284
rect 28252 25230 28254 25282
rect 28254 25230 28306 25282
rect 28306 25230 28308 25282
rect 28252 25228 28308 25230
rect 27916 23884 27972 23940
rect 27580 22092 27636 22148
rect 26684 21308 26740 21364
rect 27020 20578 27076 20580
rect 27020 20526 27022 20578
rect 27022 20526 27074 20578
rect 27074 20526 27076 20578
rect 27020 20524 27076 20526
rect 26796 20018 26852 20020
rect 26796 19966 26798 20018
rect 26798 19966 26850 20018
rect 26850 19966 26852 20018
rect 26796 19964 26852 19966
rect 27132 19964 27188 20020
rect 26684 19404 26740 19460
rect 27020 19292 27076 19348
rect 26908 18844 26964 18900
rect 26012 18338 26068 18340
rect 26012 18286 26014 18338
rect 26014 18286 26066 18338
rect 26066 18286 26068 18338
rect 26012 18284 26068 18286
rect 25900 17666 25956 17668
rect 25900 17614 25902 17666
rect 25902 17614 25954 17666
rect 25954 17614 25956 17666
rect 25900 17612 25956 17614
rect 25564 16098 25620 16100
rect 25564 16046 25566 16098
rect 25566 16046 25618 16098
rect 25618 16046 25620 16098
rect 25564 16044 25620 16046
rect 25228 15148 25284 15204
rect 24892 14530 24948 14532
rect 24892 14478 24894 14530
rect 24894 14478 24946 14530
rect 24946 14478 24948 14530
rect 24892 14476 24948 14478
rect 25452 14530 25508 14532
rect 25452 14478 25454 14530
rect 25454 14478 25506 14530
rect 25506 14478 25508 14530
rect 25452 14476 25508 14478
rect 25116 14306 25172 14308
rect 25116 14254 25118 14306
rect 25118 14254 25170 14306
rect 25170 14254 25172 14306
rect 25116 14252 25172 14254
rect 25116 13916 25172 13972
rect 25004 13692 25060 13748
rect 24220 7756 24276 7812
rect 24668 11788 24724 11844
rect 24780 11506 24836 11508
rect 24780 11454 24782 11506
rect 24782 11454 24834 11506
rect 24834 11454 24836 11506
rect 24780 11452 24836 11454
rect 24892 10444 24948 10500
rect 24332 9772 24388 9828
rect 24892 9826 24948 9828
rect 24892 9774 24894 9826
rect 24894 9774 24946 9826
rect 24946 9774 24948 9826
rect 24892 9772 24948 9774
rect 24220 7586 24276 7588
rect 24220 7534 24222 7586
rect 24222 7534 24274 7586
rect 24274 7534 24276 7586
rect 24220 7532 24276 7534
rect 23324 5404 23380 5460
rect 23436 5740 23492 5796
rect 23436 5346 23492 5348
rect 23436 5294 23438 5346
rect 23438 5294 23490 5346
rect 23490 5294 23492 5346
rect 23436 5292 23492 5294
rect 26012 17276 26068 17332
rect 26348 17052 26404 17108
rect 25788 16882 25844 16884
rect 25788 16830 25790 16882
rect 25790 16830 25842 16882
rect 25842 16830 25844 16882
rect 25788 16828 25844 16830
rect 26572 16882 26628 16884
rect 26572 16830 26574 16882
rect 26574 16830 26626 16882
rect 26626 16830 26628 16882
rect 26572 16828 26628 16830
rect 27692 21532 27748 21588
rect 27580 20524 27636 20580
rect 27692 20300 27748 20356
rect 27468 20018 27524 20020
rect 27468 19966 27470 20018
rect 27470 19966 27522 20018
rect 27522 19966 27524 20018
rect 27468 19964 27524 19966
rect 27580 19234 27636 19236
rect 27580 19182 27582 19234
rect 27582 19182 27634 19234
rect 27634 19182 27636 19234
rect 27580 19180 27636 19182
rect 28140 23212 28196 23268
rect 27916 21644 27972 21700
rect 28028 22876 28084 22932
rect 28700 27020 28756 27076
rect 28588 26460 28644 26516
rect 28588 25900 28644 25956
rect 28588 25394 28644 25396
rect 28588 25342 28590 25394
rect 28590 25342 28642 25394
rect 28642 25342 28644 25394
rect 28588 25340 28644 25342
rect 29596 29986 29652 29988
rect 29596 29934 29598 29986
rect 29598 29934 29650 29986
rect 29650 29934 29652 29986
rect 29596 29932 29652 29934
rect 29708 29708 29764 29764
rect 29484 28812 29540 28868
rect 29372 28588 29428 28644
rect 30156 29538 30212 29540
rect 30156 29486 30158 29538
rect 30158 29486 30210 29538
rect 30210 29486 30212 29538
rect 30156 29484 30212 29486
rect 29932 28924 29988 28980
rect 29820 28588 29876 28644
rect 29260 28476 29316 28532
rect 29148 28364 29204 28420
rect 28588 24556 28644 24612
rect 28252 22652 28308 22708
rect 28140 22370 28196 22372
rect 28140 22318 28142 22370
rect 28142 22318 28194 22370
rect 28194 22318 28196 22370
rect 28140 22316 28196 22318
rect 28476 20860 28532 20916
rect 27692 18844 27748 18900
rect 27916 20524 27972 20580
rect 27916 20076 27972 20132
rect 28252 20748 28308 20804
rect 28140 19346 28196 19348
rect 28140 19294 28142 19346
rect 28142 19294 28194 19346
rect 28194 19294 28196 19346
rect 28140 19292 28196 19294
rect 28364 20636 28420 20692
rect 28700 22146 28756 22148
rect 28700 22094 28702 22146
rect 28702 22094 28754 22146
rect 28754 22094 28756 22146
rect 28700 22092 28756 22094
rect 28700 19292 28756 19348
rect 28924 28252 28980 28308
rect 29372 27804 29428 27860
rect 29148 27186 29204 27188
rect 29148 27134 29150 27186
rect 29150 27134 29202 27186
rect 29202 27134 29204 27186
rect 29148 27132 29204 27134
rect 29820 27858 29876 27860
rect 29820 27806 29822 27858
rect 29822 27806 29874 27858
rect 29874 27806 29876 27858
rect 29820 27804 29876 27806
rect 29708 27132 29764 27188
rect 29484 27020 29540 27076
rect 29148 26348 29204 26404
rect 30940 29708 30996 29764
rect 30380 29484 30436 29540
rect 31052 29484 31108 29540
rect 31500 29708 31556 29764
rect 30828 29372 30884 29428
rect 31388 28924 31444 28980
rect 31052 28812 31108 28868
rect 30380 28700 30436 28756
rect 30604 26908 30660 26964
rect 29708 26236 29764 26292
rect 29596 25676 29652 25732
rect 29484 25506 29540 25508
rect 29484 25454 29486 25506
rect 29486 25454 29538 25506
rect 29538 25454 29540 25506
rect 29484 25452 29540 25454
rect 29148 25228 29204 25284
rect 29036 21698 29092 21700
rect 29036 21646 29038 21698
rect 29038 21646 29090 21698
rect 29090 21646 29092 21698
rect 29036 21644 29092 21646
rect 29260 21644 29316 21700
rect 30940 25900 30996 25956
rect 31276 26796 31332 26852
rect 30604 25676 30660 25732
rect 30044 25564 30100 25620
rect 29932 23884 29988 23940
rect 29708 21868 29764 21924
rect 29036 20300 29092 20356
rect 29148 20860 29204 20916
rect 30492 25004 30548 25060
rect 30156 23772 30212 23828
rect 30268 24668 30324 24724
rect 31052 25282 31108 25284
rect 31052 25230 31054 25282
rect 31054 25230 31106 25282
rect 31106 25230 31108 25282
rect 31052 25228 31108 25230
rect 31612 29372 31668 29428
rect 31836 29314 31892 29316
rect 31836 29262 31838 29314
rect 31838 29262 31890 29314
rect 31890 29262 31892 29314
rect 31836 29260 31892 29262
rect 32060 29932 32116 29988
rect 31948 28812 32004 28868
rect 31612 28754 31668 28756
rect 31612 28702 31614 28754
rect 31614 28702 31666 28754
rect 31666 28702 31668 28754
rect 31612 28700 31668 28702
rect 32508 33516 32564 33572
rect 33516 33852 33572 33908
rect 32508 32786 32564 32788
rect 32508 32734 32510 32786
rect 32510 32734 32562 32786
rect 32562 32734 32564 32786
rect 32508 32732 32564 32734
rect 32620 31890 32676 31892
rect 32620 31838 32622 31890
rect 32622 31838 32674 31890
rect 32674 31838 32676 31890
rect 32620 31836 32676 31838
rect 33068 31724 33124 31780
rect 33180 31388 33236 31444
rect 33068 31106 33124 31108
rect 33068 31054 33070 31106
rect 33070 31054 33122 31106
rect 33122 31054 33124 31106
rect 33068 31052 33124 31054
rect 33180 30994 33236 30996
rect 33180 30942 33182 30994
rect 33182 30942 33234 30994
rect 33234 30942 33236 30994
rect 33180 30940 33236 30942
rect 35532 40124 35588 40180
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35084 39730 35140 39732
rect 35084 39678 35086 39730
rect 35086 39678 35138 39730
rect 35138 39678 35140 39730
rect 35084 39676 35140 39678
rect 34412 39618 34468 39620
rect 34412 39566 34414 39618
rect 34414 39566 34466 39618
rect 34466 39566 34468 39618
rect 34412 39564 34468 39566
rect 35196 39564 35252 39620
rect 34076 39340 34132 39396
rect 35980 39730 36036 39732
rect 35980 39678 35982 39730
rect 35982 39678 36034 39730
rect 36034 39678 36036 39730
rect 35980 39676 36036 39678
rect 35644 38892 35700 38948
rect 33964 35980 34020 36036
rect 34188 37996 34244 38052
rect 34748 38108 34804 38164
rect 34412 37884 34468 37940
rect 34300 37378 34356 37380
rect 34300 37326 34302 37378
rect 34302 37326 34354 37378
rect 34354 37326 34356 37378
rect 34300 37324 34356 37326
rect 34860 37884 34916 37940
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35084 38108 35140 38164
rect 35868 38162 35924 38164
rect 35868 38110 35870 38162
rect 35870 38110 35922 38162
rect 35922 38110 35924 38162
rect 35868 38108 35924 38110
rect 35308 37826 35364 37828
rect 35308 37774 35310 37826
rect 35310 37774 35362 37826
rect 35362 37774 35364 37826
rect 35308 37772 35364 37774
rect 35196 37378 35252 37380
rect 35196 37326 35198 37378
rect 35198 37326 35250 37378
rect 35250 37326 35252 37378
rect 35196 37324 35252 37326
rect 36876 41020 36932 41076
rect 36988 40684 37044 40740
rect 37212 41804 37268 41860
rect 37100 40626 37156 40628
rect 37100 40574 37102 40626
rect 37102 40574 37154 40626
rect 37154 40574 37156 40626
rect 37100 40572 37156 40574
rect 36764 40402 36820 40404
rect 36764 40350 36766 40402
rect 36766 40350 36818 40402
rect 36818 40350 36820 40402
rect 36764 40348 36820 40350
rect 37436 41580 37492 41636
rect 37436 41186 37492 41188
rect 37436 41134 37438 41186
rect 37438 41134 37490 41186
rect 37490 41134 37492 41186
rect 37436 41132 37492 41134
rect 37660 42924 37716 42980
rect 38780 44716 38836 44772
rect 38220 44268 38276 44324
rect 38108 44156 38164 44212
rect 37996 43820 38052 43876
rect 37884 43372 37940 43428
rect 38108 43708 38164 43764
rect 38332 44156 38388 44212
rect 38332 43820 38388 43876
rect 38332 43650 38388 43652
rect 38332 43598 38334 43650
rect 38334 43598 38386 43650
rect 38386 43598 38388 43650
rect 38332 43596 38388 43598
rect 39228 44828 39284 44884
rect 40348 46060 40404 46116
rect 41244 46060 41300 46116
rect 39340 44716 39396 44772
rect 38556 43372 38612 43428
rect 39340 44044 39396 44100
rect 39228 43596 39284 43652
rect 39004 43036 39060 43092
rect 38892 42812 38948 42868
rect 38332 42028 38388 42084
rect 38668 42028 38724 42084
rect 38892 42082 38948 42084
rect 38892 42030 38894 42082
rect 38894 42030 38946 42082
rect 38946 42030 38948 42082
rect 38892 42028 38948 42030
rect 37884 41468 37940 41524
rect 37548 40908 37604 40964
rect 37772 40572 37828 40628
rect 37996 40460 38052 40516
rect 37212 40124 37268 40180
rect 36876 39788 36932 39844
rect 37772 40348 37828 40404
rect 37772 39900 37828 39956
rect 37324 39340 37380 39396
rect 37436 39788 37492 39844
rect 38108 40684 38164 40740
rect 38668 41356 38724 41412
rect 38108 40348 38164 40404
rect 39228 42530 39284 42532
rect 39228 42478 39230 42530
rect 39230 42478 39282 42530
rect 39282 42478 39284 42530
rect 39228 42476 39284 42478
rect 39116 41356 39172 41412
rect 39004 41132 39060 41188
rect 38108 39900 38164 39956
rect 36092 38220 36148 38276
rect 36876 38722 36932 38724
rect 36876 38670 36878 38722
rect 36878 38670 36930 38722
rect 36930 38670 36932 38722
rect 36876 38668 36932 38670
rect 35980 37436 36036 37492
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 34748 36428 34804 36484
rect 35084 36316 35140 36372
rect 34188 35756 34244 35812
rect 34076 35252 34132 35308
rect 33852 34972 33908 35028
rect 34188 34972 34244 35028
rect 34972 34972 35028 35028
rect 34300 34914 34356 34916
rect 34300 34862 34302 34914
rect 34302 34862 34354 34914
rect 34354 34862 34356 34914
rect 34300 34860 34356 34862
rect 33852 32956 33908 33012
rect 34188 32396 34244 32452
rect 33516 31724 33572 31780
rect 33740 31388 33796 31444
rect 33292 30716 33348 30772
rect 33852 30882 33908 30884
rect 33852 30830 33854 30882
rect 33854 30830 33906 30882
rect 33906 30830 33908 30882
rect 33852 30828 33908 30830
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35308 35084 35364 35140
rect 35196 34914 35252 34916
rect 35196 34862 35198 34914
rect 35198 34862 35250 34914
rect 35250 34862 35252 34914
rect 35196 34860 35252 34862
rect 35252 34636 35308 34692
rect 35420 34524 35476 34580
rect 36092 37884 36148 37940
rect 36204 37772 36260 37828
rect 36204 37212 36260 37268
rect 35644 36764 35700 36820
rect 36316 36764 36372 36820
rect 36652 38220 36708 38276
rect 35756 36370 35812 36372
rect 35756 36318 35758 36370
rect 35758 36318 35810 36370
rect 35810 36318 35812 36370
rect 35756 36316 35812 36318
rect 35980 36092 36036 36148
rect 35644 35868 35700 35924
rect 36540 36092 36596 36148
rect 37212 38892 37268 38948
rect 37660 39394 37716 39396
rect 37660 39342 37662 39394
rect 37662 39342 37714 39394
rect 37714 39342 37716 39394
rect 37660 39340 37716 39342
rect 37884 39004 37940 39060
rect 37212 38668 37268 38724
rect 37772 37938 37828 37940
rect 37772 37886 37774 37938
rect 37774 37886 37826 37938
rect 37826 37886 37828 37938
rect 37772 37884 37828 37886
rect 36988 37378 37044 37380
rect 36988 37326 36990 37378
rect 36990 37326 37042 37378
rect 37042 37326 37044 37378
rect 36988 37324 37044 37326
rect 37212 37212 37268 37268
rect 37436 37436 37492 37492
rect 37100 36652 37156 36708
rect 36988 36370 37044 36372
rect 36988 36318 36990 36370
rect 36990 36318 37042 36370
rect 37042 36318 37044 36370
rect 36988 36316 37044 36318
rect 38220 39788 38276 39844
rect 38780 38834 38836 38836
rect 38780 38782 38782 38834
rect 38782 38782 38834 38834
rect 38834 38782 38836 38834
rect 38780 38780 38836 38782
rect 39788 44268 39844 44324
rect 39900 44210 39956 44212
rect 39900 44158 39902 44210
rect 39902 44158 39954 44210
rect 39954 44158 39956 44210
rect 39900 44156 39956 44158
rect 40012 44828 40068 44884
rect 39676 43372 39732 43428
rect 40012 43148 40068 43204
rect 40348 44716 40404 44772
rect 40236 43484 40292 43540
rect 39788 42028 39844 42084
rect 39900 41916 39956 41972
rect 39452 41580 39508 41636
rect 39676 41186 39732 41188
rect 39676 41134 39678 41186
rect 39678 41134 39730 41186
rect 39730 41134 39732 41186
rect 39676 41132 39732 41134
rect 40124 42924 40180 42980
rect 40012 40908 40068 40964
rect 39228 40796 39284 40852
rect 40012 40402 40068 40404
rect 40012 40350 40014 40402
rect 40014 40350 40066 40402
rect 40066 40350 40068 40402
rect 40012 40348 40068 40350
rect 40012 40124 40068 40180
rect 41132 43426 41188 43428
rect 41132 43374 41134 43426
rect 41134 43374 41186 43426
rect 41186 43374 41188 43426
rect 41132 43372 41188 43374
rect 41356 42812 41412 42868
rect 40460 41804 40516 41860
rect 40572 42588 40628 42644
rect 40348 41746 40404 41748
rect 40348 41694 40350 41746
rect 40350 41694 40402 41746
rect 40402 41694 40404 41746
rect 40348 41692 40404 41694
rect 40236 40626 40292 40628
rect 40236 40574 40238 40626
rect 40238 40574 40290 40626
rect 40290 40574 40292 40626
rect 40236 40572 40292 40574
rect 40348 40514 40404 40516
rect 40348 40462 40350 40514
rect 40350 40462 40402 40514
rect 40402 40462 40404 40514
rect 40348 40460 40404 40462
rect 40236 40124 40292 40180
rect 40012 39058 40068 39060
rect 40012 39006 40014 39058
rect 40014 39006 40066 39058
rect 40066 39006 40068 39058
rect 40012 39004 40068 39006
rect 39004 38668 39060 38724
rect 40348 39004 40404 39060
rect 38220 37826 38276 37828
rect 38220 37774 38222 37826
rect 38222 37774 38274 37826
rect 38274 37774 38276 37826
rect 38220 37772 38276 37774
rect 38220 37436 38276 37492
rect 39116 37826 39172 37828
rect 39116 37774 39118 37826
rect 39118 37774 39170 37826
rect 39170 37774 39172 37826
rect 39116 37772 39172 37774
rect 39900 37826 39956 37828
rect 39900 37774 39902 37826
rect 39902 37774 39954 37826
rect 39954 37774 39956 37826
rect 39900 37772 39956 37774
rect 38780 37324 38836 37380
rect 39116 37324 39172 37380
rect 37996 36706 38052 36708
rect 37996 36654 37998 36706
rect 37998 36654 38050 36706
rect 38050 36654 38052 36706
rect 37996 36652 38052 36654
rect 37884 36316 37940 36372
rect 38556 36370 38612 36372
rect 38556 36318 38558 36370
rect 38558 36318 38610 36370
rect 38610 36318 38612 36370
rect 38556 36316 38612 36318
rect 36316 35532 36372 35588
rect 38556 35756 38612 35812
rect 37436 35308 37492 35364
rect 35980 35026 36036 35028
rect 35980 34974 35982 35026
rect 35982 34974 36034 35026
rect 36034 34974 36036 35026
rect 35980 34972 36036 34974
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35420 33458 35476 33460
rect 35420 33406 35422 33458
rect 35422 33406 35474 33458
rect 35474 33406 35476 33458
rect 35420 33404 35476 33406
rect 35868 34524 35924 34580
rect 36204 34914 36260 34916
rect 36204 34862 36206 34914
rect 36206 34862 36258 34914
rect 36258 34862 36260 34914
rect 36204 34860 36260 34862
rect 36428 34748 36484 34804
rect 36316 34636 36372 34692
rect 35868 33404 35924 33460
rect 35756 33234 35812 33236
rect 35756 33182 35758 33234
rect 35758 33182 35810 33234
rect 35810 33182 35812 33234
rect 35756 33180 35812 33182
rect 36428 33292 36484 33348
rect 36092 33180 36148 33236
rect 34636 31612 34692 31668
rect 34524 31052 34580 31108
rect 35084 32620 35140 32676
rect 34860 31164 34916 31220
rect 34860 30940 34916 30996
rect 36428 32674 36484 32676
rect 36428 32622 36430 32674
rect 36430 32622 36482 32674
rect 36482 32622 36484 32674
rect 36428 32620 36484 32622
rect 35980 32450 36036 32452
rect 35980 32398 35982 32450
rect 35982 32398 36034 32450
rect 36034 32398 36036 32450
rect 35980 32396 36036 32398
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35644 31666 35700 31668
rect 35644 31614 35646 31666
rect 35646 31614 35698 31666
rect 35698 31614 35700 31666
rect 35644 31612 35700 31614
rect 35756 31052 35812 31108
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35756 30268 35812 30324
rect 32284 29708 32340 29764
rect 33180 29426 33236 29428
rect 33180 29374 33182 29426
rect 33182 29374 33234 29426
rect 33234 29374 33236 29426
rect 33180 29372 33236 29374
rect 34188 30156 34244 30212
rect 33740 29372 33796 29428
rect 32844 28924 32900 28980
rect 34524 29596 34580 29652
rect 35868 30940 35924 30996
rect 34972 29596 35028 29652
rect 36428 30380 36484 30436
rect 36092 30268 36148 30324
rect 33068 28642 33124 28644
rect 33068 28590 33070 28642
rect 33070 28590 33122 28642
rect 33122 28590 33124 28642
rect 33068 28588 33124 28590
rect 34412 28476 34468 28532
rect 31836 27020 31892 27076
rect 32172 27186 32228 27188
rect 32172 27134 32174 27186
rect 32174 27134 32226 27186
rect 32226 27134 32228 27186
rect 32172 27132 32228 27134
rect 31276 25394 31332 25396
rect 31276 25342 31278 25394
rect 31278 25342 31330 25394
rect 31330 25342 31332 25394
rect 31276 25340 31332 25342
rect 30940 24722 30996 24724
rect 30940 24670 30942 24722
rect 30942 24670 30994 24722
rect 30994 24670 30996 24722
rect 30940 24668 30996 24670
rect 30268 23548 30324 23604
rect 29932 22652 29988 22708
rect 30268 22988 30324 23044
rect 29820 20860 29876 20916
rect 29932 20972 29988 21028
rect 29372 20802 29428 20804
rect 29372 20750 29374 20802
rect 29374 20750 29426 20802
rect 29426 20750 29428 20802
rect 29372 20748 29428 20750
rect 29708 19516 29764 19572
rect 29484 19234 29540 19236
rect 29484 19182 29486 19234
rect 29486 19182 29538 19234
rect 29538 19182 29540 19234
rect 29484 19180 29540 19182
rect 31276 25004 31332 25060
rect 30940 24220 30996 24276
rect 30828 24108 30884 24164
rect 30828 23324 30884 23380
rect 30828 23042 30884 23044
rect 30828 22990 30830 23042
rect 30830 22990 30882 23042
rect 30882 22990 30884 23042
rect 30828 22988 30884 22990
rect 31388 24108 31444 24164
rect 31388 23436 31444 23492
rect 31164 22988 31220 23044
rect 31500 23324 31556 23380
rect 32060 26460 32116 26516
rect 31836 26290 31892 26292
rect 31836 26238 31838 26290
rect 31838 26238 31890 26290
rect 31890 26238 31892 26290
rect 31836 26236 31892 26238
rect 31836 25900 31892 25956
rect 31948 25340 32004 25396
rect 31724 24108 31780 24164
rect 32172 25394 32228 25396
rect 32172 25342 32174 25394
rect 32174 25342 32226 25394
rect 32226 25342 32228 25394
rect 32172 25340 32228 25342
rect 32284 24668 32340 24724
rect 32172 24220 32228 24276
rect 33404 27916 33460 27972
rect 34076 27970 34132 27972
rect 34076 27918 34078 27970
rect 34078 27918 34130 27970
rect 34130 27918 34132 27970
rect 34076 27916 34132 27918
rect 33516 27746 33572 27748
rect 33516 27694 33518 27746
rect 33518 27694 33570 27746
rect 33570 27694 33572 27746
rect 33516 27692 33572 27694
rect 33404 27132 33460 27188
rect 32844 26572 32900 26628
rect 33628 26290 33684 26292
rect 33628 26238 33630 26290
rect 33630 26238 33682 26290
rect 33682 26238 33684 26290
rect 33628 26236 33684 26238
rect 32844 26124 32900 26180
rect 31724 23266 31780 23268
rect 31724 23214 31726 23266
rect 31726 23214 31778 23266
rect 31778 23214 31780 23266
rect 31724 23212 31780 23214
rect 31724 22540 31780 22596
rect 31276 21868 31332 21924
rect 31500 22092 31556 22148
rect 30492 21698 30548 21700
rect 30492 21646 30494 21698
rect 30494 21646 30546 21698
rect 30546 21646 30548 21698
rect 30492 21644 30548 21646
rect 30604 21532 30660 21588
rect 31052 21586 31108 21588
rect 31052 21534 31054 21586
rect 31054 21534 31106 21586
rect 31106 21534 31108 21586
rect 31052 21532 31108 21534
rect 30716 20748 30772 20804
rect 30604 20412 30660 20468
rect 30156 19346 30212 19348
rect 30156 19294 30158 19346
rect 30158 19294 30210 19346
rect 30210 19294 30212 19346
rect 30156 19292 30212 19294
rect 30268 18844 30324 18900
rect 28364 17500 28420 17556
rect 27132 17164 27188 17220
rect 27692 17052 27748 17108
rect 26908 16882 26964 16884
rect 26908 16830 26910 16882
rect 26910 16830 26962 16882
rect 26962 16830 26964 16882
rect 26908 16828 26964 16830
rect 26684 16380 26740 16436
rect 26796 16268 26852 16324
rect 25900 15986 25956 15988
rect 25900 15934 25902 15986
rect 25902 15934 25954 15986
rect 25954 15934 25956 15986
rect 25900 15932 25956 15934
rect 26012 14812 26068 14868
rect 25788 14476 25844 14532
rect 26460 14812 26516 14868
rect 25676 14028 25732 14084
rect 27132 16604 27188 16660
rect 27244 15484 27300 15540
rect 27356 15372 27412 15428
rect 26684 14306 26740 14308
rect 26684 14254 26686 14306
rect 26686 14254 26738 14306
rect 26738 14254 26740 14306
rect 26684 14252 26740 14254
rect 26124 13916 26180 13972
rect 26572 14140 26628 14196
rect 27132 14924 27188 14980
rect 25564 13580 25620 13636
rect 25676 13468 25732 13524
rect 26348 13468 26404 13524
rect 25676 13244 25732 13300
rect 25228 12962 25284 12964
rect 25228 12910 25230 12962
rect 25230 12910 25282 12962
rect 25282 12910 25284 12962
rect 25228 12908 25284 12910
rect 25340 12402 25396 12404
rect 25340 12350 25342 12402
rect 25342 12350 25394 12402
rect 25394 12350 25396 12402
rect 25340 12348 25396 12350
rect 25116 12124 25172 12180
rect 26348 12402 26404 12404
rect 26348 12350 26350 12402
rect 26350 12350 26402 12402
rect 26402 12350 26404 12402
rect 26348 12348 26404 12350
rect 26572 13244 26628 13300
rect 26012 12290 26068 12292
rect 26012 12238 26014 12290
rect 26014 12238 26066 12290
rect 26066 12238 26068 12290
rect 26012 12236 26068 12238
rect 27020 13634 27076 13636
rect 27020 13582 27022 13634
rect 27022 13582 27074 13634
rect 27074 13582 27076 13634
rect 27020 13580 27076 13582
rect 26124 12124 26180 12180
rect 25340 11228 25396 11284
rect 26796 12572 26852 12628
rect 26348 12012 26404 12068
rect 26460 11900 26516 11956
rect 26348 10668 26404 10724
rect 25228 10498 25284 10500
rect 25228 10446 25230 10498
rect 25230 10446 25282 10498
rect 25282 10446 25284 10498
rect 25228 10444 25284 10446
rect 25564 9324 25620 9380
rect 24668 8428 24724 8484
rect 24556 7474 24612 7476
rect 24556 7422 24558 7474
rect 24558 7422 24610 7474
rect 24610 7422 24612 7474
rect 24556 7420 24612 7422
rect 24556 6972 24612 7028
rect 23772 5852 23828 5908
rect 23884 5516 23940 5572
rect 24108 5906 24164 5908
rect 24108 5854 24110 5906
rect 24110 5854 24162 5906
rect 24162 5854 24164 5906
rect 24108 5852 24164 5854
rect 24556 6018 24612 6020
rect 24556 5966 24558 6018
rect 24558 5966 24610 6018
rect 24610 5966 24612 6018
rect 24556 5964 24612 5966
rect 24332 5516 24388 5572
rect 24556 5628 24612 5684
rect 23660 4956 23716 5012
rect 24444 5346 24500 5348
rect 24444 5294 24446 5346
rect 24446 5294 24498 5346
rect 24498 5294 24500 5346
rect 24444 5292 24500 5294
rect 24108 4562 24164 4564
rect 24108 4510 24110 4562
rect 24110 4510 24162 4562
rect 24162 4510 24164 4562
rect 24108 4508 24164 4510
rect 23660 4226 23716 4228
rect 23660 4174 23662 4226
rect 23662 4174 23714 4226
rect 23714 4174 23716 4226
rect 23660 4172 23716 4174
rect 24108 3666 24164 3668
rect 24108 3614 24110 3666
rect 24110 3614 24162 3666
rect 24162 3614 24164 3666
rect 24108 3612 24164 3614
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 21084 2828 21140 2884
rect 25116 7532 25172 7588
rect 25004 7308 25060 7364
rect 24892 6690 24948 6692
rect 24892 6638 24894 6690
rect 24894 6638 24946 6690
rect 24946 6638 24948 6690
rect 24892 6636 24948 6638
rect 24780 5404 24836 5460
rect 23660 3164 23716 3220
rect 18508 2492 18564 2548
rect 23660 2492 23716 2548
rect 25676 9212 25732 9268
rect 26012 9266 26068 9268
rect 26012 9214 26014 9266
rect 26014 9214 26066 9266
rect 26066 9214 26068 9266
rect 26012 9212 26068 9214
rect 25900 8258 25956 8260
rect 25900 8206 25902 8258
rect 25902 8206 25954 8258
rect 25954 8206 25956 8258
rect 25900 8204 25956 8206
rect 25788 7586 25844 7588
rect 25788 7534 25790 7586
rect 25790 7534 25842 7586
rect 25842 7534 25844 7586
rect 25788 7532 25844 7534
rect 27020 12236 27076 12292
rect 27468 16716 27524 16772
rect 27916 16658 27972 16660
rect 27916 16606 27918 16658
rect 27918 16606 27970 16658
rect 27970 16606 27972 16658
rect 27916 16604 27972 16606
rect 27468 15260 27524 15316
rect 27580 16380 27636 16436
rect 28364 16604 28420 16660
rect 28476 16828 28532 16884
rect 27916 15874 27972 15876
rect 27916 15822 27918 15874
rect 27918 15822 27970 15874
rect 27970 15822 27972 15874
rect 27916 15820 27972 15822
rect 27580 14700 27636 14756
rect 28140 14812 28196 14868
rect 28028 14642 28084 14644
rect 28028 14590 28030 14642
rect 28030 14590 28082 14642
rect 28082 14590 28084 14642
rect 28028 14588 28084 14590
rect 27692 14476 27748 14532
rect 27468 13746 27524 13748
rect 27468 13694 27470 13746
rect 27470 13694 27522 13746
rect 27522 13694 27524 13746
rect 27468 13692 27524 13694
rect 27356 13356 27412 13412
rect 27356 13132 27412 13188
rect 28140 14476 28196 14532
rect 28140 13074 28196 13076
rect 28140 13022 28142 13074
rect 28142 13022 28194 13074
rect 28194 13022 28196 13074
rect 28140 13020 28196 13022
rect 27468 12236 27524 12292
rect 27580 12124 27636 12180
rect 28364 15260 28420 15316
rect 29932 18508 29988 18564
rect 29260 18172 29316 18228
rect 29148 17836 29204 17892
rect 28812 16940 28868 16996
rect 28924 17276 28980 17332
rect 28588 16716 28644 16772
rect 28700 16882 28756 16884
rect 28700 16830 28702 16882
rect 28702 16830 28754 16882
rect 28754 16830 28756 16882
rect 28700 16828 28756 16830
rect 28588 15708 28644 15764
rect 28588 14812 28644 14868
rect 28924 16828 28980 16884
rect 29596 18450 29652 18452
rect 29596 18398 29598 18450
rect 29598 18398 29650 18450
rect 29650 18398 29652 18450
rect 29596 18396 29652 18398
rect 28700 14924 28756 14980
rect 28588 14642 28644 14644
rect 28588 14590 28590 14642
rect 28590 14590 28642 14642
rect 28642 14590 28644 14642
rect 28588 14588 28644 14590
rect 28700 13916 28756 13972
rect 29148 16716 29204 16772
rect 27356 10780 27412 10836
rect 27244 10332 27300 10388
rect 26460 9266 26516 9268
rect 26460 9214 26462 9266
rect 26462 9214 26514 9266
rect 26514 9214 26516 9266
rect 26460 9212 26516 9214
rect 26796 9100 26852 9156
rect 26348 8146 26404 8148
rect 26348 8094 26350 8146
rect 26350 8094 26402 8146
rect 26402 8094 26404 8146
rect 26348 8092 26404 8094
rect 26124 7308 26180 7364
rect 26348 7532 26404 7588
rect 25564 6018 25620 6020
rect 25564 5966 25566 6018
rect 25566 5966 25618 6018
rect 25618 5966 25620 6018
rect 25564 5964 25620 5966
rect 25340 5906 25396 5908
rect 25340 5854 25342 5906
rect 25342 5854 25394 5906
rect 25394 5854 25396 5906
rect 25340 5852 25396 5854
rect 25788 5906 25844 5908
rect 25788 5854 25790 5906
rect 25790 5854 25842 5906
rect 25842 5854 25844 5906
rect 25788 5852 25844 5854
rect 25788 5122 25844 5124
rect 25788 5070 25790 5122
rect 25790 5070 25842 5122
rect 25842 5070 25844 5122
rect 25788 5068 25844 5070
rect 25004 5010 25060 5012
rect 25004 4958 25006 5010
rect 25006 4958 25058 5010
rect 25058 4958 25060 5010
rect 25004 4956 25060 4958
rect 26124 6130 26180 6132
rect 26124 6078 26126 6130
rect 26126 6078 26178 6130
rect 26178 6078 26180 6130
rect 26124 6076 26180 6078
rect 26572 7980 26628 8036
rect 26460 7420 26516 7476
rect 26348 7362 26404 7364
rect 26348 7310 26350 7362
rect 26350 7310 26402 7362
rect 26402 7310 26404 7362
rect 26348 7308 26404 7310
rect 26684 6636 26740 6692
rect 27132 9996 27188 10052
rect 27020 8652 27076 8708
rect 27132 7980 27188 8036
rect 27580 8316 27636 8372
rect 26908 6860 26964 6916
rect 26796 6076 26852 6132
rect 26460 5234 26516 5236
rect 26460 5182 26462 5234
rect 26462 5182 26514 5234
rect 26514 5182 26516 5234
rect 26460 5180 26516 5182
rect 26236 4562 26292 4564
rect 26236 4510 26238 4562
rect 26238 4510 26290 4562
rect 26290 4510 26292 4562
rect 26236 4508 26292 4510
rect 24892 1596 24948 1652
rect 24556 1372 24612 1428
rect 15036 1260 15092 1316
rect 27020 6300 27076 6356
rect 27020 5964 27076 6020
rect 27468 7308 27524 7364
rect 27132 6748 27188 6804
rect 27356 6690 27412 6692
rect 27356 6638 27358 6690
rect 27358 6638 27410 6690
rect 27410 6638 27412 6690
rect 27356 6636 27412 6638
rect 27356 6300 27412 6356
rect 27916 11788 27972 11844
rect 27804 11170 27860 11172
rect 27804 11118 27806 11170
rect 27806 11118 27858 11170
rect 27858 11118 27860 11170
rect 27804 11116 27860 11118
rect 28140 12178 28196 12180
rect 28140 12126 28142 12178
rect 28142 12126 28194 12178
rect 28194 12126 28196 12178
rect 28140 12124 28196 12126
rect 28476 12402 28532 12404
rect 28476 12350 28478 12402
rect 28478 12350 28530 12402
rect 28530 12350 28532 12402
rect 28476 12348 28532 12350
rect 28700 12460 28756 12516
rect 28140 11116 28196 11172
rect 28140 10780 28196 10836
rect 27804 10332 27860 10388
rect 27804 9996 27860 10052
rect 27804 8652 27860 8708
rect 27804 7698 27860 7700
rect 27804 7646 27806 7698
rect 27806 7646 27858 7698
rect 27858 7646 27860 7698
rect 27804 7644 27860 7646
rect 28252 9660 28308 9716
rect 28588 9772 28644 9828
rect 28140 8764 28196 8820
rect 28476 9602 28532 9604
rect 28476 9550 28478 9602
rect 28478 9550 28530 9602
rect 28530 9550 28532 9602
rect 28476 9548 28532 9550
rect 28588 8370 28644 8372
rect 28588 8318 28590 8370
rect 28590 8318 28642 8370
rect 28642 8318 28644 8370
rect 28588 8316 28644 8318
rect 28140 8034 28196 8036
rect 28140 7982 28142 8034
rect 28142 7982 28194 8034
rect 28194 7982 28196 8034
rect 28140 7980 28196 7982
rect 29372 15986 29428 15988
rect 29372 15934 29374 15986
rect 29374 15934 29426 15986
rect 29426 15934 29428 15986
rect 29372 15932 29428 15934
rect 30044 16828 30100 16884
rect 29708 14700 29764 14756
rect 29372 14140 29428 14196
rect 29372 13970 29428 13972
rect 29372 13918 29374 13970
rect 29374 13918 29426 13970
rect 29426 13918 29428 13970
rect 29372 13916 29428 13918
rect 30940 20300 30996 20356
rect 30828 19628 30884 19684
rect 30492 19234 30548 19236
rect 30492 19182 30494 19234
rect 30494 19182 30546 19234
rect 30546 19182 30548 19234
rect 30492 19180 30548 19182
rect 31164 20412 31220 20468
rect 31052 19516 31108 19572
rect 31276 19292 31332 19348
rect 32060 23324 32116 23380
rect 32284 21868 32340 21924
rect 32508 23996 32564 24052
rect 32732 24108 32788 24164
rect 32508 23154 32564 23156
rect 32508 23102 32510 23154
rect 32510 23102 32562 23154
rect 32562 23102 32564 23154
rect 32508 23100 32564 23102
rect 32508 21586 32564 21588
rect 32508 21534 32510 21586
rect 32510 21534 32562 21586
rect 32562 21534 32564 21586
rect 32508 21532 32564 21534
rect 31836 20524 31892 20580
rect 31836 20300 31892 20356
rect 33068 25340 33124 25396
rect 34300 27692 34356 27748
rect 33964 26684 34020 26740
rect 33516 25116 33572 25172
rect 33068 24780 33124 24836
rect 34076 26178 34132 26180
rect 34076 26126 34078 26178
rect 34078 26126 34130 26178
rect 34130 26126 34132 26178
rect 34076 26124 34132 26126
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 34748 28866 34804 28868
rect 34748 28814 34750 28866
rect 34750 28814 34802 28866
rect 34802 28814 34804 28866
rect 34748 28812 34804 28814
rect 35308 28476 35364 28532
rect 35532 28140 35588 28196
rect 35868 28642 35924 28644
rect 35868 28590 35870 28642
rect 35870 28590 35922 28642
rect 35922 28590 35924 28642
rect 35868 28588 35924 28590
rect 35756 28364 35812 28420
rect 34636 27468 34692 27524
rect 34524 25900 34580 25956
rect 34524 25676 34580 25732
rect 34300 25228 34356 25284
rect 33852 24610 33908 24612
rect 33852 24558 33854 24610
rect 33854 24558 33906 24610
rect 33906 24558 33908 24610
rect 33852 24556 33908 24558
rect 34524 23548 34580 23604
rect 32956 22652 33012 22708
rect 32956 21980 33012 22036
rect 32284 20802 32340 20804
rect 32284 20750 32286 20802
rect 32286 20750 32338 20802
rect 32338 20750 32340 20802
rect 32284 20748 32340 20750
rect 31724 19404 31780 19460
rect 32060 19740 32116 19796
rect 31612 19180 31668 19236
rect 31500 19068 31556 19124
rect 31948 18508 32004 18564
rect 31388 18396 31444 18452
rect 31164 17724 31220 17780
rect 30380 16770 30436 16772
rect 30380 16718 30382 16770
rect 30382 16718 30434 16770
rect 30434 16718 30436 16770
rect 30380 16716 30436 16718
rect 30268 16098 30324 16100
rect 30268 16046 30270 16098
rect 30270 16046 30322 16098
rect 30322 16046 30324 16098
rect 30268 16044 30324 16046
rect 30156 14812 30212 14868
rect 30380 14700 30436 14756
rect 30492 15036 30548 15092
rect 30044 13916 30100 13972
rect 29036 12236 29092 12292
rect 29372 12402 29428 12404
rect 29372 12350 29374 12402
rect 29374 12350 29426 12402
rect 29426 12350 29428 12402
rect 29372 12348 29428 12350
rect 29484 12178 29540 12180
rect 29484 12126 29486 12178
rect 29486 12126 29538 12178
rect 29538 12126 29540 12178
rect 29484 12124 29540 12126
rect 29260 11788 29316 11844
rect 29260 10780 29316 10836
rect 29372 10220 29428 10276
rect 29932 13074 29988 13076
rect 29932 13022 29934 13074
rect 29934 13022 29986 13074
rect 29986 13022 29988 13074
rect 29932 13020 29988 13022
rect 29820 12290 29876 12292
rect 29820 12238 29822 12290
rect 29822 12238 29874 12290
rect 29874 12238 29876 12290
rect 29820 12236 29876 12238
rect 29708 11788 29764 11844
rect 30044 11788 30100 11844
rect 30156 12124 30212 12180
rect 29708 11394 29764 11396
rect 29708 11342 29710 11394
rect 29710 11342 29762 11394
rect 29762 11342 29764 11394
rect 29708 11340 29764 11342
rect 30156 10668 30212 10724
rect 29596 10332 29652 10388
rect 30044 10444 30100 10500
rect 29372 9324 29428 9380
rect 29484 9212 29540 9268
rect 29148 9154 29204 9156
rect 29148 9102 29150 9154
rect 29150 9102 29202 9154
rect 29202 9102 29204 9154
rect 29148 9100 29204 9102
rect 29820 9154 29876 9156
rect 29820 9102 29822 9154
rect 29822 9102 29874 9154
rect 29874 9102 29876 9154
rect 29820 9100 29876 9102
rect 30156 10332 30212 10388
rect 30380 14140 30436 14196
rect 30828 16098 30884 16100
rect 30828 16046 30830 16098
rect 30830 16046 30882 16098
rect 30882 16046 30884 16098
rect 30828 16044 30884 16046
rect 31276 16882 31332 16884
rect 31276 16830 31278 16882
rect 31278 16830 31330 16882
rect 31330 16830 31332 16882
rect 31276 16828 31332 16830
rect 31500 17948 31556 18004
rect 32508 19906 32564 19908
rect 32508 19854 32510 19906
rect 32510 19854 32562 19906
rect 32562 19854 32564 19906
rect 32508 19852 32564 19854
rect 32396 19180 32452 19236
rect 32172 18956 32228 19012
rect 32060 16882 32116 16884
rect 32060 16830 32062 16882
rect 32062 16830 32114 16882
rect 32114 16830 32116 16882
rect 32060 16828 32116 16830
rect 31500 16716 31556 16772
rect 31164 15036 31220 15092
rect 32844 19740 32900 19796
rect 33964 23042 34020 23044
rect 33964 22990 33966 23042
rect 33966 22990 34018 23042
rect 34018 22990 34020 23042
rect 33964 22988 34020 22990
rect 33628 21980 33684 22036
rect 33068 21420 33124 21476
rect 33292 21420 33348 21476
rect 33180 20914 33236 20916
rect 33180 20862 33182 20914
rect 33182 20862 33234 20914
rect 33234 20862 33236 20914
rect 33180 20860 33236 20862
rect 32732 16044 32788 16100
rect 32620 15986 32676 15988
rect 32620 15934 32622 15986
rect 32622 15934 32674 15986
rect 32674 15934 32676 15986
rect 32620 15932 32676 15934
rect 31612 15820 31668 15876
rect 31948 15874 32004 15876
rect 31948 15822 31950 15874
rect 31950 15822 32002 15874
rect 32002 15822 32004 15874
rect 31948 15820 32004 15822
rect 30828 14812 30884 14868
rect 30828 14140 30884 14196
rect 30492 11788 30548 11844
rect 30268 9436 30324 9492
rect 29596 8988 29652 9044
rect 30828 11788 30884 11844
rect 30828 11340 30884 11396
rect 32172 15708 32228 15764
rect 32060 15314 32116 15316
rect 32060 15262 32062 15314
rect 32062 15262 32114 15314
rect 32114 15262 32116 15314
rect 32060 15260 32116 15262
rect 31948 15148 32004 15204
rect 31612 14028 31668 14084
rect 31164 13580 31220 13636
rect 31164 12348 31220 12404
rect 30940 10780 30996 10836
rect 30828 10610 30884 10612
rect 30828 10558 30830 10610
rect 30830 10558 30882 10610
rect 30882 10558 30884 10610
rect 30828 10556 30884 10558
rect 30716 10498 30772 10500
rect 30716 10446 30718 10498
rect 30718 10446 30770 10498
rect 30770 10446 30772 10498
rect 30716 10444 30772 10446
rect 30940 10444 30996 10500
rect 31052 12012 31108 12068
rect 32060 13468 32116 13524
rect 32060 12460 32116 12516
rect 31276 12290 31332 12292
rect 31276 12238 31278 12290
rect 31278 12238 31330 12290
rect 31330 12238 31332 12290
rect 31276 12236 31332 12238
rect 31388 11564 31444 11620
rect 31836 12290 31892 12292
rect 31836 12238 31838 12290
rect 31838 12238 31890 12290
rect 31890 12238 31892 12290
rect 31836 12236 31892 12238
rect 31612 12012 31668 12068
rect 31948 11340 32004 11396
rect 30604 9212 30660 9268
rect 30828 9660 30884 9716
rect 31164 9548 31220 9604
rect 30828 9042 30884 9044
rect 30828 8990 30830 9042
rect 30830 8990 30882 9042
rect 30882 8990 30884 9042
rect 30828 8988 30884 8990
rect 29708 8204 29764 8260
rect 29148 8034 29204 8036
rect 29148 7982 29150 8034
rect 29150 7982 29202 8034
rect 29202 7982 29204 8034
rect 29148 7980 29204 7982
rect 28364 6860 28420 6916
rect 28028 6636 28084 6692
rect 27804 6412 27860 6468
rect 27916 6524 27972 6580
rect 27356 6076 27412 6132
rect 27468 5740 27524 5796
rect 27244 5180 27300 5236
rect 26236 3612 26292 3668
rect 27468 5068 27524 5124
rect 27804 5852 27860 5908
rect 28364 6130 28420 6132
rect 28364 6078 28366 6130
rect 28366 6078 28418 6130
rect 28418 6078 28420 6130
rect 28364 6076 28420 6078
rect 28028 5068 28084 5124
rect 28140 5740 28196 5796
rect 28588 6018 28644 6020
rect 28588 5966 28590 6018
rect 28590 5966 28642 6018
rect 28642 5966 28644 6018
rect 28588 5964 28644 5966
rect 28476 5906 28532 5908
rect 28476 5854 28478 5906
rect 28478 5854 28530 5906
rect 28530 5854 28532 5906
rect 28476 5852 28532 5854
rect 28588 3666 28644 3668
rect 28588 3614 28590 3666
rect 28590 3614 28642 3666
rect 28642 3614 28644 3666
rect 28588 3612 28644 3614
rect 29372 8034 29428 8036
rect 29372 7982 29374 8034
rect 29374 7982 29426 8034
rect 29426 7982 29428 8034
rect 29372 7980 29428 7982
rect 29484 7644 29540 7700
rect 29596 8146 29652 8148
rect 29596 8094 29598 8146
rect 29598 8094 29650 8146
rect 29650 8094 29652 8146
rect 29596 8092 29652 8094
rect 29596 7196 29652 7252
rect 28812 6748 28868 6804
rect 29484 6188 29540 6244
rect 29148 5964 29204 6020
rect 29036 5794 29092 5796
rect 29036 5742 29038 5794
rect 29038 5742 29090 5794
rect 29090 5742 29092 5794
rect 29036 5740 29092 5742
rect 29596 6412 29652 6468
rect 30268 8034 30324 8036
rect 30268 7982 30270 8034
rect 30270 7982 30322 8034
rect 30322 7982 30324 8034
rect 30268 7980 30324 7982
rect 30492 8092 30548 8148
rect 30380 7644 30436 7700
rect 30268 7420 30324 7476
rect 29932 6690 29988 6692
rect 29932 6638 29934 6690
rect 29934 6638 29986 6690
rect 29986 6638 29988 6690
rect 29932 6636 29988 6638
rect 30268 6188 30324 6244
rect 30380 7308 30436 7364
rect 30492 6636 30548 6692
rect 30604 6076 30660 6132
rect 30604 5906 30660 5908
rect 30604 5854 30606 5906
rect 30606 5854 30658 5906
rect 30658 5854 30660 5906
rect 30604 5852 30660 5854
rect 31164 9154 31220 9156
rect 31164 9102 31166 9154
rect 31166 9102 31218 9154
rect 31218 9102 31220 9154
rect 31164 9100 31220 9102
rect 31276 8146 31332 8148
rect 31276 8094 31278 8146
rect 31278 8094 31330 8146
rect 31330 8094 31332 8146
rect 31276 8092 31332 8094
rect 30940 7644 30996 7700
rect 31276 7474 31332 7476
rect 31276 7422 31278 7474
rect 31278 7422 31330 7474
rect 31330 7422 31332 7474
rect 31276 7420 31332 7422
rect 32508 14140 32564 14196
rect 32396 14028 32452 14084
rect 32172 11340 32228 11396
rect 32060 10556 32116 10612
rect 31948 10498 32004 10500
rect 31948 10446 31950 10498
rect 31950 10446 32002 10498
rect 32002 10446 32004 10498
rect 31948 10444 32004 10446
rect 32172 10444 32228 10500
rect 31948 9154 32004 9156
rect 31948 9102 31950 9154
rect 31950 9102 32002 9154
rect 32002 9102 32004 9154
rect 31948 9100 32004 9102
rect 31836 9042 31892 9044
rect 31836 8990 31838 9042
rect 31838 8990 31890 9042
rect 31890 8990 31892 9042
rect 31836 8988 31892 8990
rect 33180 19180 33236 19236
rect 33068 19122 33124 19124
rect 33068 19070 33070 19122
rect 33070 19070 33122 19122
rect 33122 19070 33124 19122
rect 33068 19068 33124 19070
rect 32956 18956 33012 19012
rect 33516 18956 33572 19012
rect 32956 18508 33012 18564
rect 33292 17724 33348 17780
rect 33964 21308 34020 21364
rect 34076 21084 34132 21140
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35084 27074 35140 27076
rect 35084 27022 35086 27074
rect 35086 27022 35138 27074
rect 35138 27022 35140 27074
rect 35084 27020 35140 27022
rect 35420 26290 35476 26292
rect 35420 26238 35422 26290
rect 35422 26238 35474 26290
rect 35474 26238 35476 26290
rect 35420 26236 35476 26238
rect 34972 26124 35028 26180
rect 35868 26012 35924 26068
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35980 25676 36036 25732
rect 34972 25506 35028 25508
rect 34972 25454 34974 25506
rect 34974 25454 35026 25506
rect 35026 25454 35028 25506
rect 34972 25452 35028 25454
rect 37212 34690 37268 34692
rect 37212 34638 37214 34690
rect 37214 34638 37266 34690
rect 37266 34638 37268 34690
rect 37212 34636 37268 34638
rect 40348 37154 40404 37156
rect 40348 37102 40350 37154
rect 40350 37102 40402 37154
rect 40402 37102 40404 37154
rect 40348 37100 40404 37102
rect 39340 36482 39396 36484
rect 39340 36430 39342 36482
rect 39342 36430 39394 36482
rect 39394 36430 39396 36482
rect 39340 36428 39396 36430
rect 39676 36482 39732 36484
rect 39676 36430 39678 36482
rect 39678 36430 39730 36482
rect 39730 36430 39732 36482
rect 39676 36428 39732 36430
rect 39228 36316 39284 36372
rect 39564 36092 39620 36148
rect 38892 35810 38948 35812
rect 38892 35758 38894 35810
rect 38894 35758 38946 35810
rect 38946 35758 38948 35810
rect 38892 35756 38948 35758
rect 38780 35308 38836 35364
rect 36988 33234 37044 33236
rect 36988 33182 36990 33234
rect 36990 33182 37042 33234
rect 37042 33182 37044 33234
rect 36988 33180 37044 33182
rect 37996 33516 38052 33572
rect 37324 33458 37380 33460
rect 37324 33406 37326 33458
rect 37326 33406 37378 33458
rect 37378 33406 37380 33458
rect 37324 33404 37380 33406
rect 39004 34076 39060 34132
rect 38668 33292 38724 33348
rect 38780 33740 38836 33796
rect 37212 33122 37268 33124
rect 37212 33070 37214 33122
rect 37214 33070 37266 33122
rect 37266 33070 37268 33122
rect 37212 33068 37268 33070
rect 37436 33122 37492 33124
rect 37436 33070 37438 33122
rect 37438 33070 37490 33122
rect 37490 33070 37492 33122
rect 37436 33068 37492 33070
rect 37100 32396 37156 32452
rect 38108 33122 38164 33124
rect 38108 33070 38110 33122
rect 38110 33070 38162 33122
rect 38162 33070 38164 33122
rect 38108 33068 38164 33070
rect 38332 32844 38388 32900
rect 37884 32396 37940 32452
rect 37548 30492 37604 30548
rect 37996 31836 38052 31892
rect 38220 32450 38276 32452
rect 38220 32398 38222 32450
rect 38222 32398 38274 32450
rect 38274 32398 38276 32450
rect 38220 32396 38276 32398
rect 38220 31554 38276 31556
rect 38220 31502 38222 31554
rect 38222 31502 38274 31554
rect 38274 31502 38276 31554
rect 38220 31500 38276 31502
rect 38556 31948 38612 32004
rect 38668 31836 38724 31892
rect 38780 31500 38836 31556
rect 39116 33852 39172 33908
rect 38668 31388 38724 31444
rect 36988 30156 37044 30212
rect 36316 28812 36372 28868
rect 36428 28924 36484 28980
rect 36540 28700 36596 28756
rect 36988 29036 37044 29092
rect 37100 30380 37156 30436
rect 37884 30380 37940 30436
rect 37324 30268 37380 30324
rect 37212 29426 37268 29428
rect 37212 29374 37214 29426
rect 37214 29374 37266 29426
rect 37266 29374 37268 29426
rect 37212 29372 37268 29374
rect 38332 29820 38388 29876
rect 38556 30268 38612 30324
rect 36764 28364 36820 28420
rect 36876 28924 36932 28980
rect 36428 28140 36484 28196
rect 36428 26124 36484 26180
rect 36092 25452 36148 25508
rect 34860 25340 34916 25396
rect 35420 25394 35476 25396
rect 35420 25342 35422 25394
rect 35422 25342 35474 25394
rect 35474 25342 35476 25394
rect 35420 25340 35476 25342
rect 35196 25282 35252 25284
rect 35196 25230 35198 25282
rect 35198 25230 35250 25282
rect 35250 25230 35252 25282
rect 35196 25228 35252 25230
rect 34748 24780 34804 24836
rect 34972 25116 35028 25172
rect 34748 24610 34804 24612
rect 34748 24558 34750 24610
rect 34750 24558 34802 24610
rect 34802 24558 34804 24610
rect 34748 24556 34804 24558
rect 35084 24722 35140 24724
rect 35084 24670 35086 24722
rect 35086 24670 35138 24722
rect 35138 24670 35140 24722
rect 35084 24668 35140 24670
rect 35868 24610 35924 24612
rect 35868 24558 35870 24610
rect 35870 24558 35922 24610
rect 35922 24558 35924 24610
rect 35868 24556 35924 24558
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35756 23660 35812 23716
rect 35868 23548 35924 23604
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 36540 25282 36596 25284
rect 36540 25230 36542 25282
rect 36542 25230 36594 25282
rect 36594 25230 36596 25282
rect 36540 25228 36596 25230
rect 34860 21474 34916 21476
rect 34860 21422 34862 21474
rect 34862 21422 34914 21474
rect 34914 21422 34916 21474
rect 34860 21420 34916 21422
rect 34524 21084 34580 21140
rect 34188 20690 34244 20692
rect 34188 20638 34190 20690
rect 34190 20638 34242 20690
rect 34242 20638 34244 20690
rect 34188 20636 34244 20638
rect 33964 20524 34020 20580
rect 34076 20130 34132 20132
rect 34076 20078 34078 20130
rect 34078 20078 34130 20130
rect 34130 20078 34132 20130
rect 34076 20076 34132 20078
rect 33628 18508 33684 18564
rect 33852 19292 33908 19348
rect 33852 18450 33908 18452
rect 33852 18398 33854 18450
rect 33854 18398 33906 18450
rect 33906 18398 33908 18450
rect 33852 18396 33908 18398
rect 33628 17554 33684 17556
rect 33628 17502 33630 17554
rect 33630 17502 33682 17554
rect 33682 17502 33684 17554
rect 33628 17500 33684 17502
rect 33068 16940 33124 16996
rect 33068 16492 33124 16548
rect 33068 16044 33124 16100
rect 33180 15538 33236 15540
rect 33180 15486 33182 15538
rect 33182 15486 33234 15538
rect 33234 15486 33236 15538
rect 33180 15484 33236 15486
rect 33852 17724 33908 17780
rect 34412 20412 34468 20468
rect 34636 20300 34692 20356
rect 34636 19404 34692 19460
rect 34300 19292 34356 19348
rect 34972 19122 35028 19124
rect 34972 19070 34974 19122
rect 34974 19070 35026 19122
rect 35026 19070 35028 19122
rect 34972 19068 35028 19070
rect 34524 18956 34580 19012
rect 34188 18844 34244 18900
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35420 20524 35476 20580
rect 35308 20130 35364 20132
rect 35308 20078 35310 20130
rect 35310 20078 35362 20130
rect 35362 20078 35364 20130
rect 35308 20076 35364 20078
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35420 19404 35476 19460
rect 34524 17666 34580 17668
rect 34524 17614 34526 17666
rect 34526 17614 34578 17666
rect 34578 17614 34580 17666
rect 34524 17612 34580 17614
rect 34188 17554 34244 17556
rect 34188 17502 34190 17554
rect 34190 17502 34242 17554
rect 34242 17502 34244 17554
rect 34188 17500 34244 17502
rect 33628 15820 33684 15876
rect 33404 15426 33460 15428
rect 33404 15374 33406 15426
rect 33406 15374 33458 15426
rect 33458 15374 33460 15426
rect 33404 15372 33460 15374
rect 32844 15148 32900 15204
rect 33628 14642 33684 14644
rect 33628 14590 33630 14642
rect 33630 14590 33682 14642
rect 33682 14590 33684 14642
rect 33628 14588 33684 14590
rect 34300 15986 34356 15988
rect 34300 15934 34302 15986
rect 34302 15934 34354 15986
rect 34354 15934 34356 15986
rect 34300 15932 34356 15934
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 34972 17948 35028 18004
rect 35420 16828 35476 16884
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 34860 15596 34916 15652
rect 35308 15932 35364 15988
rect 35420 15596 35476 15652
rect 35756 22092 35812 22148
rect 35868 19010 35924 19012
rect 35868 18958 35870 19010
rect 35870 18958 35922 19010
rect 35922 18958 35924 19010
rect 35868 18956 35924 18958
rect 37100 28642 37156 28644
rect 37100 28590 37102 28642
rect 37102 28590 37154 28642
rect 37154 28590 37156 28642
rect 37100 28588 37156 28590
rect 36988 28530 37044 28532
rect 36988 28478 36990 28530
rect 36990 28478 37042 28530
rect 37042 28478 37044 28530
rect 36988 28476 37044 28478
rect 37212 28418 37268 28420
rect 37212 28366 37214 28418
rect 37214 28366 37266 28418
rect 37266 28366 37268 28418
rect 37212 28364 37268 28366
rect 37212 28140 37268 28196
rect 38108 29036 38164 29092
rect 37436 28924 37492 28980
rect 37436 28700 37492 28756
rect 37436 27020 37492 27076
rect 38780 29148 38836 29204
rect 38556 28812 38612 28868
rect 38220 28364 38276 28420
rect 38444 28140 38500 28196
rect 37212 26572 37268 26628
rect 36988 26460 37044 26516
rect 39340 35922 39396 35924
rect 39340 35870 39342 35922
rect 39342 35870 39394 35922
rect 39394 35870 39396 35922
rect 39340 35868 39396 35870
rect 40124 35756 40180 35812
rect 40348 36204 40404 36260
rect 40348 35196 40404 35252
rect 39676 34130 39732 34132
rect 39676 34078 39678 34130
rect 39678 34078 39730 34130
rect 39730 34078 39732 34130
rect 39676 34076 39732 34078
rect 39340 33346 39396 33348
rect 39340 33294 39342 33346
rect 39342 33294 39394 33346
rect 39394 33294 39396 33346
rect 39340 33292 39396 33294
rect 39340 32396 39396 32452
rect 40124 33628 40180 33684
rect 40236 32620 40292 32676
rect 40348 32732 40404 32788
rect 40012 32508 40068 32564
rect 40012 31948 40068 32004
rect 39340 31890 39396 31892
rect 39340 31838 39342 31890
rect 39342 31838 39394 31890
rect 39394 31838 39396 31890
rect 39340 31836 39396 31838
rect 39340 31500 39396 31556
rect 40908 41804 40964 41860
rect 40684 40572 40740 40628
rect 40796 38892 40852 38948
rect 41132 41970 41188 41972
rect 41132 41918 41134 41970
rect 41134 41918 41186 41970
rect 41186 41918 41188 41970
rect 41132 41916 41188 41918
rect 41468 41916 41524 41972
rect 41132 40796 41188 40852
rect 41468 40348 41524 40404
rect 41804 41858 41860 41860
rect 41804 41806 41806 41858
rect 41806 41806 41858 41858
rect 41858 41806 41860 41858
rect 41804 41804 41860 41806
rect 41692 41692 41748 41748
rect 41804 41132 41860 41188
rect 41020 39058 41076 39060
rect 41020 39006 41022 39058
rect 41022 39006 41074 39058
rect 41074 39006 41076 39058
rect 41020 39004 41076 39006
rect 41580 39900 41636 39956
rect 41468 39004 41524 39060
rect 42140 42140 42196 42196
rect 42812 45666 42868 45668
rect 42812 45614 42814 45666
rect 42814 45614 42866 45666
rect 42866 45614 42868 45666
rect 42812 45612 42868 45614
rect 44604 46114 44660 46116
rect 44604 46062 44606 46114
rect 44606 46062 44658 46114
rect 44658 46062 44660 46114
rect 44604 46060 44660 46062
rect 43260 45500 43316 45556
rect 43148 44492 43204 44548
rect 43036 43820 43092 43876
rect 42700 43484 42756 43540
rect 42476 42812 42532 42868
rect 43260 43372 43316 43428
rect 43708 42866 43764 42868
rect 43708 42814 43710 42866
rect 43710 42814 43762 42866
rect 43762 42814 43764 42866
rect 43708 42812 43764 42814
rect 43148 42476 43204 42532
rect 42588 41916 42644 41972
rect 42476 41186 42532 41188
rect 42476 41134 42478 41186
rect 42478 41134 42530 41186
rect 42530 41134 42532 41186
rect 42476 41132 42532 41134
rect 42588 40796 42644 40852
rect 42364 40124 42420 40180
rect 42028 39452 42084 39508
rect 42476 39900 42532 39956
rect 42700 40236 42756 40292
rect 42812 41692 42868 41748
rect 43372 41916 43428 41972
rect 43484 42028 43540 42084
rect 42924 41244 42980 41300
rect 43372 40572 43428 40628
rect 43484 40460 43540 40516
rect 42588 39452 42644 39508
rect 42028 39058 42084 39060
rect 42028 39006 42030 39058
rect 42030 39006 42082 39058
rect 42082 39006 42084 39058
rect 42028 39004 42084 39006
rect 42252 39228 42308 39284
rect 42476 38946 42532 38948
rect 42476 38894 42478 38946
rect 42478 38894 42530 38946
rect 42530 38894 42532 38946
rect 42476 38892 42532 38894
rect 42588 38780 42644 38836
rect 40796 37938 40852 37940
rect 40796 37886 40798 37938
rect 40798 37886 40850 37938
rect 40850 37886 40852 37938
rect 40796 37884 40852 37886
rect 41916 37938 41972 37940
rect 41916 37886 41918 37938
rect 41918 37886 41970 37938
rect 41970 37886 41972 37938
rect 41916 37884 41972 37886
rect 41132 37772 41188 37828
rect 41804 37772 41860 37828
rect 41132 37378 41188 37380
rect 41132 37326 41134 37378
rect 41134 37326 41186 37378
rect 41186 37326 41188 37378
rect 41132 37324 41188 37326
rect 41132 36092 41188 36148
rect 41468 36258 41524 36260
rect 41468 36206 41470 36258
rect 41470 36206 41522 36258
rect 41522 36206 41524 36258
rect 41468 36204 41524 36206
rect 41356 35980 41412 36036
rect 41244 35586 41300 35588
rect 41244 35534 41246 35586
rect 41246 35534 41298 35586
rect 41298 35534 41300 35586
rect 41244 35532 41300 35534
rect 41916 37100 41972 37156
rect 42140 36482 42196 36484
rect 42140 36430 42142 36482
rect 42142 36430 42194 36482
rect 42194 36430 42196 36482
rect 42140 36428 42196 36430
rect 42700 37100 42756 37156
rect 42364 36370 42420 36372
rect 42364 36318 42366 36370
rect 42366 36318 42418 36370
rect 42418 36318 42420 36370
rect 42364 36316 42420 36318
rect 42476 36258 42532 36260
rect 42476 36206 42478 36258
rect 42478 36206 42530 36258
rect 42530 36206 42532 36258
rect 42476 36204 42532 36206
rect 42140 36092 42196 36148
rect 41692 35698 41748 35700
rect 41692 35646 41694 35698
rect 41694 35646 41746 35698
rect 41746 35646 41748 35698
rect 41692 35644 41748 35646
rect 40908 33628 40964 33684
rect 41468 34130 41524 34132
rect 41468 34078 41470 34130
rect 41470 34078 41522 34130
rect 41522 34078 41524 34130
rect 41468 34076 41524 34078
rect 41356 33404 41412 33460
rect 41916 34860 41972 34916
rect 42476 35980 42532 36036
rect 42588 34690 42644 34692
rect 42588 34638 42590 34690
rect 42590 34638 42642 34690
rect 42642 34638 42644 34690
rect 42588 34636 42644 34638
rect 42812 35868 42868 35924
rect 41692 33740 41748 33796
rect 42252 33458 42308 33460
rect 42252 33406 42254 33458
rect 42254 33406 42306 33458
rect 42306 33406 42308 33458
rect 42252 33404 42308 33406
rect 41580 32844 41636 32900
rect 41916 32956 41972 33012
rect 41468 32732 41524 32788
rect 40908 32674 40964 32676
rect 40908 32622 40910 32674
rect 40910 32622 40962 32674
rect 40962 32622 40964 32674
rect 40908 32620 40964 32622
rect 41132 32562 41188 32564
rect 41132 32510 41134 32562
rect 41134 32510 41186 32562
rect 41186 32510 41188 32562
rect 41132 32508 41188 32510
rect 40572 32396 40628 32452
rect 40348 31164 40404 31220
rect 40124 30380 40180 30436
rect 39788 30268 39844 30324
rect 39228 28812 39284 28868
rect 39564 29372 39620 29428
rect 39004 28364 39060 28420
rect 39340 28028 39396 28084
rect 39900 29820 39956 29876
rect 40012 29538 40068 29540
rect 40012 29486 40014 29538
rect 40014 29486 40066 29538
rect 40066 29486 40068 29538
rect 40012 29484 40068 29486
rect 40236 29372 40292 29428
rect 40460 28812 40516 28868
rect 40124 28028 40180 28084
rect 38108 26572 38164 26628
rect 38668 26514 38724 26516
rect 38668 26462 38670 26514
rect 38670 26462 38722 26514
rect 38722 26462 38724 26514
rect 38668 26460 38724 26462
rect 38220 26402 38276 26404
rect 38220 26350 38222 26402
rect 38222 26350 38274 26402
rect 38274 26350 38276 26402
rect 38220 26348 38276 26350
rect 37548 25452 37604 25508
rect 37100 25116 37156 25172
rect 36988 24556 37044 24612
rect 37436 25282 37492 25284
rect 37436 25230 37438 25282
rect 37438 25230 37490 25282
rect 37490 25230 37492 25282
rect 37436 25228 37492 25230
rect 36092 21980 36148 22036
rect 36988 22092 37044 22148
rect 36428 21756 36484 21812
rect 36316 21644 36372 21700
rect 36204 21532 36260 21588
rect 36316 20802 36372 20804
rect 36316 20750 36318 20802
rect 36318 20750 36370 20802
rect 36370 20750 36372 20802
rect 36316 20748 36372 20750
rect 36988 20802 37044 20804
rect 36988 20750 36990 20802
rect 36990 20750 37042 20802
rect 37042 20750 37044 20802
rect 36988 20748 37044 20750
rect 37772 25116 37828 25172
rect 38444 26290 38500 26292
rect 38444 26238 38446 26290
rect 38446 26238 38498 26290
rect 38498 26238 38500 26290
rect 38444 26236 38500 26238
rect 38892 26402 38948 26404
rect 38892 26350 38894 26402
rect 38894 26350 38946 26402
rect 38946 26350 38948 26402
rect 38892 26348 38948 26350
rect 39004 26290 39060 26292
rect 39004 26238 39006 26290
rect 39006 26238 39058 26290
rect 39058 26238 39060 26290
rect 39004 26236 39060 26238
rect 39452 26178 39508 26180
rect 39452 26126 39454 26178
rect 39454 26126 39506 26178
rect 39506 26126 39508 26178
rect 39452 26124 39508 26126
rect 40012 26178 40068 26180
rect 40012 26126 40014 26178
rect 40014 26126 40066 26178
rect 40066 26126 40068 26178
rect 40012 26124 40068 26126
rect 40012 25676 40068 25732
rect 39228 25618 39284 25620
rect 39228 25566 39230 25618
rect 39230 25566 39282 25618
rect 39282 25566 39284 25618
rect 39228 25564 39284 25566
rect 39788 25282 39844 25284
rect 39788 25230 39790 25282
rect 39790 25230 39842 25282
rect 39842 25230 39844 25282
rect 39788 25228 39844 25230
rect 39116 24892 39172 24948
rect 38780 24722 38836 24724
rect 38780 24670 38782 24722
rect 38782 24670 38834 24722
rect 38834 24670 38836 24722
rect 38780 24668 38836 24670
rect 39676 23660 39732 23716
rect 40236 25228 40292 25284
rect 40348 24834 40404 24836
rect 40348 24782 40350 24834
rect 40350 24782 40402 24834
rect 40402 24782 40404 24834
rect 40348 24780 40404 24782
rect 41020 30716 41076 30772
rect 40796 30210 40852 30212
rect 40796 30158 40798 30210
rect 40798 30158 40850 30210
rect 40850 30158 40852 30210
rect 40796 30156 40852 30158
rect 42252 31836 42308 31892
rect 41580 31500 41636 31556
rect 41468 30156 41524 30212
rect 41356 29484 41412 29540
rect 41244 29426 41300 29428
rect 41244 29374 41246 29426
rect 41246 29374 41298 29426
rect 41298 29374 41300 29426
rect 41244 29372 41300 29374
rect 41020 28082 41076 28084
rect 41020 28030 41022 28082
rect 41022 28030 41074 28082
rect 41074 28030 41076 28082
rect 41020 28028 41076 28030
rect 40796 26124 40852 26180
rect 41020 26124 41076 26180
rect 40908 25228 40964 25284
rect 40124 23714 40180 23716
rect 40124 23662 40126 23714
rect 40126 23662 40178 23714
rect 40178 23662 40180 23714
rect 40124 23660 40180 23662
rect 40012 23548 40068 23604
rect 38556 23436 38612 23492
rect 37436 22204 37492 22260
rect 37100 20524 37156 20580
rect 37212 21756 37268 21812
rect 36092 20130 36148 20132
rect 36092 20078 36094 20130
rect 36094 20078 36146 20130
rect 36146 20078 36148 20130
rect 36092 20076 36148 20078
rect 37884 21756 37940 21812
rect 37324 21698 37380 21700
rect 37324 21646 37326 21698
rect 37326 21646 37378 21698
rect 37378 21646 37380 21698
rect 37324 21644 37380 21646
rect 37660 21644 37716 21700
rect 37772 21474 37828 21476
rect 37772 21422 37774 21474
rect 37774 21422 37826 21474
rect 37826 21422 37828 21474
rect 37772 21420 37828 21422
rect 38220 23100 38276 23156
rect 38108 21644 38164 21700
rect 38444 23042 38500 23044
rect 38444 22990 38446 23042
rect 38446 22990 38498 23042
rect 38498 22990 38500 23042
rect 38444 22988 38500 22990
rect 38332 21644 38388 21700
rect 38444 21756 38500 21812
rect 37884 20524 37940 20580
rect 38444 20300 38500 20356
rect 38892 23154 38948 23156
rect 38892 23102 38894 23154
rect 38894 23102 38946 23154
rect 38946 23102 38948 23154
rect 38892 23100 38948 23102
rect 39004 22988 39060 23044
rect 39228 22930 39284 22932
rect 39228 22878 39230 22930
rect 39230 22878 39282 22930
rect 39282 22878 39284 22930
rect 39228 22876 39284 22878
rect 39004 22204 39060 22260
rect 41244 28700 41300 28756
rect 42252 29484 42308 29540
rect 41692 29314 41748 29316
rect 41692 29262 41694 29314
rect 41694 29262 41746 29314
rect 41746 29262 41748 29314
rect 41692 29260 41748 29262
rect 41356 28588 41412 28644
rect 41468 28812 41524 28868
rect 42364 31724 42420 31780
rect 42700 31554 42756 31556
rect 42700 31502 42702 31554
rect 42702 31502 42754 31554
rect 42754 31502 42756 31554
rect 42700 31500 42756 31502
rect 42140 29148 42196 29204
rect 41916 28530 41972 28532
rect 41916 28478 41918 28530
rect 41918 28478 41970 28530
rect 41970 28478 41972 28530
rect 41916 28476 41972 28478
rect 42252 28924 42308 28980
rect 41804 28140 41860 28196
rect 43260 39004 43316 39060
rect 43036 38668 43092 38724
rect 43260 38834 43316 38836
rect 43260 38782 43262 38834
rect 43262 38782 43314 38834
rect 43314 38782 43316 38834
rect 43260 38780 43316 38782
rect 43148 37772 43204 37828
rect 43260 37212 43316 37268
rect 43036 35980 43092 36036
rect 43148 36876 43204 36932
rect 43148 36428 43204 36484
rect 43484 38108 43540 38164
rect 44268 45724 44324 45780
rect 44156 44828 44212 44884
rect 44380 45612 44436 45668
rect 43932 43708 43988 43764
rect 43932 42364 43988 42420
rect 43820 41804 43876 41860
rect 43820 41132 43876 41188
rect 43708 40348 43764 40404
rect 44044 41746 44100 41748
rect 44044 41694 44046 41746
rect 44046 41694 44098 41746
rect 44098 41694 44100 41746
rect 44044 41692 44100 41694
rect 44268 42530 44324 42532
rect 44268 42478 44270 42530
rect 44270 42478 44322 42530
rect 44322 42478 44324 42530
rect 44268 42476 44324 42478
rect 45388 45612 45444 45668
rect 45276 45276 45332 45332
rect 44828 45218 44884 45220
rect 44828 45166 44830 45218
rect 44830 45166 44882 45218
rect 44882 45166 44884 45218
rect 44828 45164 44884 45166
rect 44940 45106 44996 45108
rect 44940 45054 44942 45106
rect 44942 45054 44994 45106
rect 44994 45054 44996 45106
rect 44940 45052 44996 45054
rect 44828 43820 44884 43876
rect 44492 42924 44548 42980
rect 44940 43538 44996 43540
rect 44940 43486 44942 43538
rect 44942 43486 44994 43538
rect 44994 43486 44996 43538
rect 44940 43484 44996 43486
rect 44828 42812 44884 42868
rect 45164 42812 45220 42868
rect 44268 41692 44324 41748
rect 43932 40572 43988 40628
rect 43820 40290 43876 40292
rect 43820 40238 43822 40290
rect 43822 40238 43874 40290
rect 43874 40238 43876 40290
rect 43820 40236 43876 40238
rect 44156 40908 44212 40964
rect 44380 40684 44436 40740
rect 44492 41244 44548 41300
rect 44828 41970 44884 41972
rect 44828 41918 44830 41970
rect 44830 41918 44882 41970
rect 44882 41918 44884 41970
rect 44828 41916 44884 41918
rect 45276 41858 45332 41860
rect 45276 41806 45278 41858
rect 45278 41806 45330 41858
rect 45330 41806 45332 41858
rect 45276 41804 45332 41806
rect 45052 41692 45108 41748
rect 44940 41580 44996 41636
rect 44940 41074 44996 41076
rect 44940 41022 44942 41074
rect 44942 41022 44994 41074
rect 44994 41022 44996 41074
rect 44940 41020 44996 41022
rect 44604 40908 44660 40964
rect 44940 40402 44996 40404
rect 44940 40350 44942 40402
rect 44942 40350 44994 40402
rect 44994 40350 44996 40402
rect 44940 40348 44996 40350
rect 43708 38108 43764 38164
rect 43596 37772 43652 37828
rect 42924 35644 42980 35700
rect 42924 34860 42980 34916
rect 43036 32956 43092 33012
rect 42812 30492 42868 30548
rect 44380 39452 44436 39508
rect 44044 39004 44100 39060
rect 44156 39228 44212 39284
rect 44044 38162 44100 38164
rect 44044 38110 44046 38162
rect 44046 38110 44098 38162
rect 44098 38110 44100 38162
rect 44044 38108 44100 38110
rect 43932 37154 43988 37156
rect 43932 37102 43934 37154
rect 43934 37102 43986 37154
rect 43986 37102 43988 37154
rect 43932 37100 43988 37102
rect 43820 36316 43876 36372
rect 44828 39506 44884 39508
rect 44828 39454 44830 39506
rect 44830 39454 44882 39506
rect 44882 39454 44884 39506
rect 44828 39452 44884 39454
rect 45052 39116 45108 39172
rect 44828 39058 44884 39060
rect 44828 39006 44830 39058
rect 44830 39006 44882 39058
rect 44882 39006 44884 39058
rect 44828 39004 44884 39006
rect 45276 39228 45332 39284
rect 45836 44546 45892 44548
rect 45836 44494 45838 44546
rect 45838 44494 45890 44546
rect 45890 44494 45892 44546
rect 45836 44492 45892 44494
rect 48412 47068 48468 47124
rect 46508 45778 46564 45780
rect 46508 45726 46510 45778
rect 46510 45726 46562 45778
rect 46562 45726 46564 45778
rect 46508 45724 46564 45726
rect 46732 45500 46788 45556
rect 45948 43596 46004 43652
rect 46844 44828 46900 44884
rect 45612 43484 45668 43540
rect 45500 43148 45556 43204
rect 45500 41916 45556 41972
rect 45836 42978 45892 42980
rect 45836 42926 45838 42978
rect 45838 42926 45890 42978
rect 45890 42926 45892 42978
rect 45836 42924 45892 42926
rect 46620 42476 46676 42532
rect 45500 40460 45556 40516
rect 45388 39004 45444 39060
rect 44828 38780 44884 38836
rect 46284 41804 46340 41860
rect 46284 40796 46340 40852
rect 45948 40460 46004 40516
rect 45836 40402 45892 40404
rect 45836 40350 45838 40402
rect 45838 40350 45890 40402
rect 45890 40350 45892 40402
rect 45836 40348 45892 40350
rect 44828 38220 44884 38276
rect 45500 38780 45556 38836
rect 45164 38220 45220 38276
rect 45052 38108 45108 38164
rect 44492 37436 44548 37492
rect 44940 37154 44996 37156
rect 44940 37102 44942 37154
rect 44942 37102 44994 37154
rect 44994 37102 44996 37154
rect 44940 37100 44996 37102
rect 43820 35980 43876 36036
rect 43596 35868 43652 35924
rect 43596 35698 43652 35700
rect 43596 35646 43598 35698
rect 43598 35646 43650 35698
rect 43650 35646 43652 35698
rect 43596 35644 43652 35646
rect 44604 36316 44660 36372
rect 44268 35980 44324 36036
rect 44044 35532 44100 35588
rect 45164 37938 45220 37940
rect 45164 37886 45166 37938
rect 45166 37886 45218 37938
rect 45218 37886 45220 37938
rect 45164 37884 45220 37886
rect 45164 36258 45220 36260
rect 45164 36206 45166 36258
rect 45166 36206 45218 36258
rect 45218 36206 45220 36258
rect 45164 36204 45220 36206
rect 44492 35532 44548 35588
rect 44268 34802 44324 34804
rect 44268 34750 44270 34802
rect 44270 34750 44322 34802
rect 44322 34750 44324 34802
rect 44268 34748 44324 34750
rect 44380 34636 44436 34692
rect 43372 32956 43428 33012
rect 43708 33180 43764 33236
rect 43820 33122 43876 33124
rect 43820 33070 43822 33122
rect 43822 33070 43874 33122
rect 43874 33070 43876 33122
rect 43820 33068 43876 33070
rect 43372 30604 43428 30660
rect 43260 30156 43316 30212
rect 45724 37100 45780 37156
rect 45388 36988 45444 37044
rect 45500 35980 45556 36036
rect 46508 40626 46564 40628
rect 46508 40574 46510 40626
rect 46510 40574 46562 40626
rect 46562 40574 46564 40626
rect 46508 40572 46564 40574
rect 46396 38332 46452 38388
rect 46060 38220 46116 38276
rect 45388 35196 45444 35252
rect 44940 34690 44996 34692
rect 44940 34638 44942 34690
rect 44942 34638 44994 34690
rect 44994 34638 44996 34690
rect 44940 34636 44996 34638
rect 44828 33234 44884 33236
rect 44828 33182 44830 33234
rect 44830 33182 44882 33234
rect 44882 33182 44884 33234
rect 44828 33180 44884 33182
rect 44380 33068 44436 33124
rect 43932 31500 43988 31556
rect 44716 31836 44772 31892
rect 44380 31612 44436 31668
rect 44828 31554 44884 31556
rect 44828 31502 44830 31554
rect 44830 31502 44882 31554
rect 44882 31502 44884 31554
rect 44828 31500 44884 31502
rect 44940 31388 44996 31444
rect 43932 30770 43988 30772
rect 43932 30718 43934 30770
rect 43934 30718 43986 30770
rect 43986 30718 43988 30770
rect 43932 30716 43988 30718
rect 43596 30492 43652 30548
rect 42700 29314 42756 29316
rect 42700 29262 42702 29314
rect 42702 29262 42754 29314
rect 42754 29262 42756 29314
rect 42700 29260 42756 29262
rect 42588 29202 42644 29204
rect 42588 29150 42590 29202
rect 42590 29150 42642 29202
rect 42642 29150 42644 29202
rect 42588 29148 42644 29150
rect 42700 28812 42756 28868
rect 43372 29484 43428 29540
rect 42812 28588 42868 28644
rect 43260 28642 43316 28644
rect 43260 28590 43262 28642
rect 43262 28590 43314 28642
rect 43314 28590 43316 28642
rect 43260 28588 43316 28590
rect 42364 28028 42420 28084
rect 41244 25116 41300 25172
rect 42140 27186 42196 27188
rect 42140 27134 42142 27186
rect 42142 27134 42194 27186
rect 42194 27134 42196 27186
rect 42140 27132 42196 27134
rect 41244 24780 41300 24836
rect 40572 22876 40628 22932
rect 40796 22428 40852 22484
rect 40460 22258 40516 22260
rect 40460 22206 40462 22258
rect 40462 22206 40514 22258
rect 40514 22206 40516 22258
rect 40460 22204 40516 22206
rect 40124 21868 40180 21924
rect 39788 21474 39844 21476
rect 39788 21422 39790 21474
rect 39790 21422 39842 21474
rect 39842 21422 39844 21474
rect 39788 21420 39844 21422
rect 39228 20914 39284 20916
rect 39228 20862 39230 20914
rect 39230 20862 39282 20914
rect 39282 20862 39284 20914
rect 39228 20860 39284 20862
rect 38780 20130 38836 20132
rect 38780 20078 38782 20130
rect 38782 20078 38834 20130
rect 38834 20078 38836 20130
rect 38780 20076 38836 20078
rect 38556 19964 38612 20020
rect 39004 20018 39060 20020
rect 39004 19966 39006 20018
rect 39006 19966 39058 20018
rect 39058 19966 39060 20018
rect 39004 19964 39060 19966
rect 36540 19404 36596 19460
rect 36652 19068 36708 19124
rect 35644 18732 35700 18788
rect 35868 15596 35924 15652
rect 35756 15484 35812 15540
rect 36652 18620 36708 18676
rect 36988 18396 37044 18452
rect 36316 17612 36372 17668
rect 35980 15484 36036 15540
rect 36092 16882 36148 16884
rect 36092 16830 36094 16882
rect 36094 16830 36146 16882
rect 36146 16830 36148 16882
rect 36092 16828 36148 16830
rect 35644 15372 35700 15428
rect 35980 15202 36036 15204
rect 35980 15150 35982 15202
rect 35982 15150 36034 15202
rect 36034 15150 36036 15202
rect 35980 15148 36036 15150
rect 36540 16882 36596 16884
rect 36540 16830 36542 16882
rect 36542 16830 36594 16882
rect 36594 16830 36596 16882
rect 36540 16828 36596 16830
rect 37100 18956 37156 19012
rect 37660 18508 37716 18564
rect 37996 19292 38052 19348
rect 38892 18674 38948 18676
rect 38892 18622 38894 18674
rect 38894 18622 38946 18674
rect 38946 18622 38948 18674
rect 38892 18620 38948 18622
rect 36988 16828 37044 16884
rect 37100 16940 37156 16996
rect 36316 16156 36372 16212
rect 36428 15314 36484 15316
rect 36428 15262 36430 15314
rect 36430 15262 36482 15314
rect 36482 15262 36484 15314
rect 36428 15260 36484 15262
rect 34188 14530 34244 14532
rect 34188 14478 34190 14530
rect 34190 14478 34242 14530
rect 34242 14478 34244 14530
rect 34188 14476 34244 14478
rect 33292 13692 33348 13748
rect 32508 10444 32564 10500
rect 33180 13468 33236 13524
rect 33180 12572 33236 12628
rect 33068 12460 33124 12516
rect 33180 11788 33236 11844
rect 33964 13746 34020 13748
rect 33964 13694 33966 13746
rect 33966 13694 34018 13746
rect 34018 13694 34020 13746
rect 33964 13692 34020 13694
rect 33516 13074 33572 13076
rect 33516 13022 33518 13074
rect 33518 13022 33570 13074
rect 33570 13022 33572 13074
rect 33516 13020 33572 13022
rect 33404 12962 33460 12964
rect 33404 12910 33406 12962
rect 33406 12910 33458 12962
rect 33458 12910 33460 12962
rect 33404 12908 33460 12910
rect 34188 13132 34244 13188
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 34524 14530 34580 14532
rect 34524 14478 34526 14530
rect 34526 14478 34578 14530
rect 34578 14478 34580 14530
rect 34524 14476 34580 14478
rect 34524 13468 34580 13524
rect 34412 13356 34468 13412
rect 34412 13132 34468 13188
rect 34972 14364 35028 14420
rect 34748 13692 34804 13748
rect 34188 12962 34244 12964
rect 34188 12910 34190 12962
rect 34190 12910 34242 12962
rect 34242 12910 34244 12962
rect 34188 12908 34244 12910
rect 34076 12684 34132 12740
rect 33740 11788 33796 11844
rect 33628 11452 33684 11508
rect 33740 11228 33796 11284
rect 33292 10668 33348 10724
rect 33628 10498 33684 10500
rect 33628 10446 33630 10498
rect 33630 10446 33682 10498
rect 33682 10446 33684 10498
rect 33628 10444 33684 10446
rect 33180 10220 33236 10276
rect 33292 10108 33348 10164
rect 33180 9714 33236 9716
rect 33180 9662 33182 9714
rect 33182 9662 33234 9714
rect 33234 9662 33236 9714
rect 33180 9660 33236 9662
rect 32284 8204 32340 8260
rect 32284 7756 32340 7812
rect 32172 7308 32228 7364
rect 30940 6300 30996 6356
rect 30828 5964 30884 6020
rect 30828 5794 30884 5796
rect 30828 5742 30830 5794
rect 30830 5742 30882 5794
rect 30882 5742 30884 5794
rect 30828 5740 30884 5742
rect 31052 5628 31108 5684
rect 29372 5010 29428 5012
rect 29372 4958 29374 5010
rect 29374 4958 29426 5010
rect 29426 4958 29428 5010
rect 29372 4956 29428 4958
rect 30268 4956 30324 5012
rect 32284 6860 32340 6916
rect 31724 6748 31780 6804
rect 31500 6690 31556 6692
rect 31500 6638 31502 6690
rect 31502 6638 31554 6690
rect 31554 6638 31556 6690
rect 31500 6636 31556 6638
rect 31276 6524 31332 6580
rect 31500 5740 31556 5796
rect 31500 5292 31556 5348
rect 31388 5180 31444 5236
rect 31612 4956 31668 5012
rect 31948 6188 32004 6244
rect 32172 5628 32228 5684
rect 32060 5068 32116 5124
rect 32396 6802 32452 6804
rect 32396 6750 32398 6802
rect 32398 6750 32450 6802
rect 32450 6750 32452 6802
rect 32396 6748 32452 6750
rect 32620 8316 32676 8372
rect 32620 7308 32676 7364
rect 32732 6972 32788 7028
rect 32620 6748 32676 6804
rect 31164 4060 31220 4116
rect 32508 5852 32564 5908
rect 33292 8204 33348 8260
rect 33292 7756 33348 7812
rect 33068 7586 33124 7588
rect 33068 7534 33070 7586
rect 33070 7534 33122 7586
rect 33122 7534 33124 7586
rect 33068 7532 33124 7534
rect 33068 6690 33124 6692
rect 33068 6638 33070 6690
rect 33070 6638 33122 6690
rect 33122 6638 33124 6690
rect 33068 6636 33124 6638
rect 34076 11618 34132 11620
rect 34076 11566 34078 11618
rect 34078 11566 34130 11618
rect 34130 11566 34132 11618
rect 34076 11564 34132 11566
rect 34076 11340 34132 11396
rect 34412 12402 34468 12404
rect 34412 12350 34414 12402
rect 34414 12350 34466 12402
rect 34466 12350 34468 12402
rect 34412 12348 34468 12350
rect 35196 13468 35252 13524
rect 35420 14252 35476 14308
rect 35420 13692 35476 13748
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35084 12962 35140 12964
rect 35084 12910 35086 12962
rect 35086 12910 35138 12962
rect 35138 12910 35140 12962
rect 35084 12908 35140 12910
rect 34748 12684 34804 12740
rect 35980 14588 36036 14644
rect 35868 14140 35924 14196
rect 35756 13132 35812 13188
rect 34860 12460 34916 12516
rect 37324 16492 37380 16548
rect 37212 16380 37268 16436
rect 37324 15538 37380 15540
rect 37324 15486 37326 15538
rect 37326 15486 37378 15538
rect 37378 15486 37380 15538
rect 37324 15484 37380 15486
rect 36540 14476 36596 14532
rect 36316 14418 36372 14420
rect 36316 14366 36318 14418
rect 36318 14366 36370 14418
rect 36370 14366 36372 14418
rect 36316 14364 36372 14366
rect 35980 13020 36036 13076
rect 36092 13692 36148 13748
rect 34636 11676 34692 11732
rect 34524 11394 34580 11396
rect 34524 11342 34526 11394
rect 34526 11342 34578 11394
rect 34578 11342 34580 11394
rect 34524 11340 34580 11342
rect 34188 11282 34244 11284
rect 34188 11230 34190 11282
rect 34190 11230 34242 11282
rect 34242 11230 34244 11282
rect 34188 11228 34244 11230
rect 34076 10892 34132 10948
rect 34524 11004 34580 11060
rect 34860 12178 34916 12180
rect 34860 12126 34862 12178
rect 34862 12126 34914 12178
rect 34914 12126 34916 12178
rect 34860 12124 34916 12126
rect 34972 12012 35028 12068
rect 34860 11900 34916 11956
rect 35532 12178 35588 12180
rect 35532 12126 35534 12178
rect 35534 12126 35586 12178
rect 35586 12126 35588 12178
rect 35532 12124 35588 12126
rect 35644 12012 35700 12068
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 34748 11452 34804 11508
rect 35084 11394 35140 11396
rect 35084 11342 35086 11394
rect 35086 11342 35138 11394
rect 35138 11342 35140 11394
rect 35084 11340 35140 11342
rect 35532 11394 35588 11396
rect 35532 11342 35534 11394
rect 35534 11342 35586 11394
rect 35586 11342 35588 11394
rect 35532 11340 35588 11342
rect 35868 11900 35924 11956
rect 36204 12348 36260 12404
rect 36316 12572 36372 12628
rect 36316 12178 36372 12180
rect 36316 12126 36318 12178
rect 36318 12126 36370 12178
rect 36370 12126 36372 12178
rect 36316 12124 36372 12126
rect 35868 11506 35924 11508
rect 35868 11454 35870 11506
rect 35870 11454 35922 11506
rect 35922 11454 35924 11506
rect 35868 11452 35924 11454
rect 34748 11170 34804 11172
rect 34748 11118 34750 11170
rect 34750 11118 34802 11170
rect 34802 11118 34804 11170
rect 34748 11116 34804 11118
rect 36092 11004 36148 11060
rect 34860 10892 34916 10948
rect 34300 10108 34356 10164
rect 34188 9660 34244 9716
rect 34412 8876 34468 8932
rect 33740 7698 33796 7700
rect 33740 7646 33742 7698
rect 33742 7646 33794 7698
rect 33794 7646 33796 7698
rect 33740 7644 33796 7646
rect 34188 8146 34244 8148
rect 34188 8094 34190 8146
rect 34190 8094 34242 8146
rect 34242 8094 34244 8146
rect 34188 8092 34244 8094
rect 33852 7868 33908 7924
rect 33852 7420 33908 7476
rect 35308 10722 35364 10724
rect 35308 10670 35310 10722
rect 35310 10670 35362 10722
rect 35362 10670 35364 10722
rect 35308 10668 35364 10670
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35308 9938 35364 9940
rect 35308 9886 35310 9938
rect 35310 9886 35362 9938
rect 35362 9886 35364 9938
rect 35308 9884 35364 9886
rect 35308 8988 35364 9044
rect 35420 8930 35476 8932
rect 35420 8878 35422 8930
rect 35422 8878 35474 8930
rect 35474 8878 35476 8930
rect 35420 8876 35476 8878
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 34748 8316 34804 8372
rect 34972 8204 35028 8260
rect 34300 7868 34356 7924
rect 33516 6860 33572 6916
rect 34860 7980 34916 8036
rect 34636 7644 34692 7700
rect 33292 6524 33348 6580
rect 32844 5852 32900 5908
rect 32956 5964 33012 6020
rect 32732 5740 32788 5796
rect 32508 5516 32564 5572
rect 33628 6412 33684 6468
rect 33180 5682 33236 5684
rect 33180 5630 33182 5682
rect 33182 5630 33234 5682
rect 33234 5630 33236 5682
rect 33180 5628 33236 5630
rect 33516 5404 33572 5460
rect 33404 5292 33460 5348
rect 28924 2940 28980 2996
rect 27580 2716 27636 2772
rect 34300 6412 34356 6468
rect 33740 5740 33796 5796
rect 34076 6076 34132 6132
rect 33964 6018 34020 6020
rect 33964 5966 33966 6018
rect 33966 5966 34018 6018
rect 34018 5966 34020 6018
rect 33964 5964 34020 5966
rect 34412 5906 34468 5908
rect 34412 5854 34414 5906
rect 34414 5854 34466 5906
rect 34466 5854 34468 5906
rect 34412 5852 34468 5854
rect 34076 5628 34132 5684
rect 33852 5516 33908 5572
rect 34188 5516 34244 5572
rect 34076 5404 34132 5460
rect 33740 5122 33796 5124
rect 33740 5070 33742 5122
rect 33742 5070 33794 5122
rect 33794 5070 33796 5122
rect 33740 5068 33796 5070
rect 33628 3164 33684 3220
rect 36204 10722 36260 10724
rect 36204 10670 36206 10722
rect 36206 10670 36258 10722
rect 36258 10670 36260 10722
rect 36204 10668 36260 10670
rect 35644 10332 35700 10388
rect 35756 10444 35812 10500
rect 35532 8204 35588 8260
rect 36876 14364 36932 14420
rect 36988 14028 37044 14084
rect 37324 14530 37380 14532
rect 37324 14478 37326 14530
rect 37326 14478 37378 14530
rect 37378 14478 37380 14530
rect 37324 14476 37380 14478
rect 37100 13692 37156 13748
rect 36540 13580 36596 13636
rect 37100 12738 37156 12740
rect 37100 12686 37102 12738
rect 37102 12686 37154 12738
rect 37154 12686 37156 12738
rect 37100 12684 37156 12686
rect 36988 12460 37044 12516
rect 36652 12402 36708 12404
rect 36652 12350 36654 12402
rect 36654 12350 36706 12402
rect 36706 12350 36708 12402
rect 36652 12348 36708 12350
rect 36540 11564 36596 11620
rect 36876 12066 36932 12068
rect 36876 12014 36878 12066
rect 36878 12014 36930 12066
rect 36930 12014 36932 12066
rect 36876 12012 36932 12014
rect 36876 11452 36932 11508
rect 36988 11788 37044 11844
rect 37100 12236 37156 12292
rect 39564 18508 39620 18564
rect 39676 19740 39732 19796
rect 39004 18396 39060 18452
rect 39900 19346 39956 19348
rect 39900 19294 39902 19346
rect 39902 19294 39954 19346
rect 39954 19294 39956 19346
rect 39900 19292 39956 19294
rect 38332 17052 38388 17108
rect 37772 16940 37828 16996
rect 37660 15986 37716 15988
rect 37660 15934 37662 15986
rect 37662 15934 37714 15986
rect 37714 15934 37716 15986
rect 37660 15932 37716 15934
rect 39004 17666 39060 17668
rect 39004 17614 39006 17666
rect 39006 17614 39058 17666
rect 39058 17614 39060 17666
rect 39004 17612 39060 17614
rect 40236 19852 40292 19908
rect 40348 18338 40404 18340
rect 40348 18286 40350 18338
rect 40350 18286 40402 18338
rect 40402 18286 40404 18338
rect 40348 18284 40404 18286
rect 40012 17612 40068 17668
rect 39004 16940 39060 16996
rect 40236 17106 40292 17108
rect 40236 17054 40238 17106
rect 40238 17054 40290 17106
rect 40290 17054 40292 17106
rect 40236 17052 40292 17054
rect 38444 16828 38500 16884
rect 37884 16098 37940 16100
rect 37884 16046 37886 16098
rect 37886 16046 37938 16098
rect 37938 16046 37940 16098
rect 37884 16044 37940 16046
rect 40124 16828 40180 16884
rect 39004 16716 39060 16772
rect 38108 15986 38164 15988
rect 38108 15934 38110 15986
rect 38110 15934 38162 15986
rect 38162 15934 38164 15986
rect 38108 15932 38164 15934
rect 38780 15932 38836 15988
rect 37996 15874 38052 15876
rect 37996 15822 37998 15874
rect 37998 15822 38050 15874
rect 38050 15822 38052 15874
rect 37996 15820 38052 15822
rect 38668 15708 38724 15764
rect 38220 15596 38276 15652
rect 38780 15148 38836 15204
rect 39228 16210 39284 16212
rect 39228 16158 39230 16210
rect 39230 16158 39282 16210
rect 39282 16158 39284 16210
rect 39228 16156 39284 16158
rect 39340 16044 39396 16100
rect 39788 16380 39844 16436
rect 39676 15820 39732 15876
rect 39900 15538 39956 15540
rect 39900 15486 39902 15538
rect 39902 15486 39954 15538
rect 39954 15486 39956 15538
rect 39900 15484 39956 15486
rect 38220 14418 38276 14420
rect 38220 14366 38222 14418
rect 38222 14366 38274 14418
rect 38274 14366 38276 14418
rect 38220 14364 38276 14366
rect 37660 14252 37716 14308
rect 37884 14252 37940 14308
rect 37772 13468 37828 13524
rect 38444 14028 38500 14084
rect 38444 13746 38500 13748
rect 38444 13694 38446 13746
rect 38446 13694 38498 13746
rect 38498 13694 38500 13746
rect 38444 13692 38500 13694
rect 39900 15148 39956 15204
rect 38892 14530 38948 14532
rect 38892 14478 38894 14530
rect 38894 14478 38946 14530
rect 38946 14478 38948 14530
rect 38892 14476 38948 14478
rect 39228 13746 39284 13748
rect 39228 13694 39230 13746
rect 39230 13694 39282 13746
rect 39282 13694 39284 13746
rect 39228 13692 39284 13694
rect 39452 13580 39508 13636
rect 37100 11340 37156 11396
rect 38332 12796 38388 12852
rect 38332 11788 38388 11844
rect 36428 10444 36484 10500
rect 35868 10332 35924 10388
rect 35644 9212 35700 9268
rect 35420 8146 35476 8148
rect 35420 8094 35422 8146
rect 35422 8094 35474 8146
rect 35474 8094 35476 8146
rect 35420 8092 35476 8094
rect 35196 8034 35252 8036
rect 35196 7982 35198 8034
rect 35198 7982 35250 8034
rect 35250 7982 35252 8034
rect 35196 7980 35252 7982
rect 35532 8034 35588 8036
rect 35532 7982 35534 8034
rect 35534 7982 35586 8034
rect 35586 7982 35588 8034
rect 35532 7980 35588 7982
rect 36540 10108 36596 10164
rect 36988 10108 37044 10164
rect 36092 9826 36148 9828
rect 36092 9774 36094 9826
rect 36094 9774 36146 9826
rect 36146 9774 36148 9826
rect 36092 9772 36148 9774
rect 37212 9996 37268 10052
rect 36652 9660 36708 9716
rect 36428 9602 36484 9604
rect 36428 9550 36430 9602
rect 36430 9550 36482 9602
rect 36482 9550 36484 9602
rect 36428 9548 36484 9550
rect 36092 9042 36148 9044
rect 36092 8990 36094 9042
rect 36094 8990 36146 9042
rect 36146 8990 36148 9042
rect 36092 8988 36148 8990
rect 35868 8652 35924 8708
rect 35980 8428 36036 8484
rect 36204 8258 36260 8260
rect 36204 8206 36206 8258
rect 36206 8206 36258 8258
rect 36258 8206 36260 8258
rect 36204 8204 36260 8206
rect 35756 8146 35812 8148
rect 35756 8094 35758 8146
rect 35758 8094 35810 8146
rect 35810 8094 35812 8146
rect 35756 8092 35812 8094
rect 35084 7756 35140 7812
rect 34860 6802 34916 6804
rect 34860 6750 34862 6802
rect 34862 6750 34914 6802
rect 34914 6750 34916 6802
rect 34860 6748 34916 6750
rect 35868 7698 35924 7700
rect 35868 7646 35870 7698
rect 35870 7646 35922 7698
rect 35922 7646 35924 7698
rect 35868 7644 35924 7646
rect 36204 7532 36260 7588
rect 37436 11618 37492 11620
rect 37436 11566 37438 11618
rect 37438 11566 37490 11618
rect 37490 11566 37492 11618
rect 37436 11564 37492 11566
rect 37548 11506 37604 11508
rect 37548 11454 37550 11506
rect 37550 11454 37602 11506
rect 37602 11454 37604 11506
rect 37548 11452 37604 11454
rect 37996 11394 38052 11396
rect 37996 11342 37998 11394
rect 37998 11342 38050 11394
rect 38050 11342 38052 11394
rect 37996 11340 38052 11342
rect 37212 9548 37268 9604
rect 37772 10386 37828 10388
rect 37772 10334 37774 10386
rect 37774 10334 37826 10386
rect 37826 10334 37828 10386
rect 37772 10332 37828 10334
rect 37100 9266 37156 9268
rect 37100 9214 37102 9266
rect 37102 9214 37154 9266
rect 37154 9214 37156 9266
rect 37100 9212 37156 9214
rect 37100 8540 37156 8596
rect 37212 8428 37268 8484
rect 37100 8370 37156 8372
rect 37100 8318 37102 8370
rect 37102 8318 37154 8370
rect 37154 8318 37156 8370
rect 37100 8316 37156 8318
rect 36764 7586 36820 7588
rect 36764 7534 36766 7586
rect 36766 7534 36818 7586
rect 36818 7534 36820 7586
rect 36764 7532 36820 7534
rect 37100 8092 37156 8148
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35644 6972 35700 7028
rect 36428 7196 36484 7252
rect 35980 6748 36036 6804
rect 34860 6300 34916 6356
rect 35196 6412 35252 6468
rect 34748 6188 34804 6244
rect 35756 6578 35812 6580
rect 35756 6526 35758 6578
rect 35758 6526 35810 6578
rect 35810 6526 35812 6578
rect 35756 6524 35812 6526
rect 35756 6188 35812 6244
rect 36988 7196 37044 7252
rect 37436 8034 37492 8036
rect 37436 7982 37438 8034
rect 37438 7982 37490 8034
rect 37490 7982 37492 8034
rect 37436 7980 37492 7982
rect 37100 7420 37156 7476
rect 36876 6748 36932 6804
rect 36316 6690 36372 6692
rect 36316 6638 36318 6690
rect 36318 6638 36370 6690
rect 36370 6638 36372 6690
rect 36316 6636 36372 6638
rect 37212 7586 37268 7588
rect 37212 7534 37214 7586
rect 37214 7534 37266 7586
rect 37266 7534 37268 7586
rect 37212 7532 37268 7534
rect 37660 10108 37716 10164
rect 37996 9826 38052 9828
rect 37996 9774 37998 9826
rect 37998 9774 38050 9826
rect 38050 9774 38052 9826
rect 37996 9772 38052 9774
rect 37772 9436 37828 9492
rect 37772 8258 37828 8260
rect 37772 8206 37774 8258
rect 37774 8206 37826 8258
rect 37826 8206 37828 8258
rect 37772 8204 37828 8206
rect 37996 8258 38052 8260
rect 37996 8206 37998 8258
rect 37998 8206 38050 8258
rect 38050 8206 38052 8258
rect 37996 8204 38052 8206
rect 38556 12796 38612 12852
rect 38444 11004 38500 11060
rect 39564 13244 39620 13300
rect 39676 13468 39732 13524
rect 39004 13020 39060 13076
rect 39004 12348 39060 12404
rect 38332 8540 38388 8596
rect 38556 10108 38612 10164
rect 38668 9660 38724 9716
rect 39228 10444 39284 10500
rect 39788 13020 39844 13076
rect 40236 15484 40292 15540
rect 40236 13746 40292 13748
rect 40236 13694 40238 13746
rect 40238 13694 40290 13746
rect 40290 13694 40292 13746
rect 40236 13692 40292 13694
rect 41916 26178 41972 26180
rect 41916 26126 41918 26178
rect 41918 26126 41970 26178
rect 41970 26126 41972 26178
rect 41916 26124 41972 26126
rect 42140 26178 42196 26180
rect 42140 26126 42142 26178
rect 42142 26126 42194 26178
rect 42194 26126 42196 26178
rect 42140 26124 42196 26126
rect 42140 25788 42196 25844
rect 42140 25452 42196 25508
rect 41580 25282 41636 25284
rect 41580 25230 41582 25282
rect 41582 25230 41634 25282
rect 41634 25230 41636 25282
rect 41580 25228 41636 25230
rect 41356 24668 41412 24724
rect 41244 23772 41300 23828
rect 41132 23548 41188 23604
rect 41132 22482 41188 22484
rect 41132 22430 41134 22482
rect 41134 22430 41186 22482
rect 41186 22430 41188 22482
rect 41132 22428 41188 22430
rect 41020 21868 41076 21924
rect 41916 25116 41972 25172
rect 41356 23660 41412 23716
rect 41580 23548 41636 23604
rect 40908 21474 40964 21476
rect 40908 21422 40910 21474
rect 40910 21422 40962 21474
rect 40962 21422 40964 21474
rect 40908 21420 40964 21422
rect 41916 23548 41972 23604
rect 42364 26402 42420 26404
rect 42364 26350 42366 26402
rect 42366 26350 42418 26402
rect 42418 26350 42420 26402
rect 42364 26348 42420 26350
rect 42812 27132 42868 27188
rect 43260 28252 43316 28308
rect 43260 26348 43316 26404
rect 42252 24722 42308 24724
rect 42252 24670 42254 24722
rect 42254 24670 42306 24722
rect 42306 24670 42308 24722
rect 42252 24668 42308 24670
rect 41692 23042 41748 23044
rect 41692 22990 41694 23042
rect 41694 22990 41746 23042
rect 41746 22990 41748 23042
rect 41692 22988 41748 22990
rect 41916 21868 41972 21924
rect 40908 17612 40964 17668
rect 41804 21362 41860 21364
rect 41804 21310 41806 21362
rect 41806 21310 41858 21362
rect 41858 21310 41860 21362
rect 41804 21308 41860 21310
rect 42476 23714 42532 23716
rect 42476 23662 42478 23714
rect 42478 23662 42530 23714
rect 42530 23662 42532 23714
rect 42476 23660 42532 23662
rect 43484 28700 43540 28756
rect 43596 28924 43652 28980
rect 43932 30268 43988 30324
rect 43820 30156 43876 30212
rect 43708 27132 43764 27188
rect 45948 36258 46004 36260
rect 45948 36206 45950 36258
rect 45950 36206 46002 36258
rect 46002 36206 46004 36258
rect 45948 36204 46004 36206
rect 47068 43596 47124 43652
rect 46956 42140 47012 42196
rect 47404 45666 47460 45668
rect 47404 45614 47406 45666
rect 47406 45614 47458 45666
rect 47458 45614 47460 45666
rect 47404 45612 47460 45614
rect 47404 45218 47460 45220
rect 47404 45166 47406 45218
rect 47406 45166 47458 45218
rect 47458 45166 47460 45218
rect 47404 45164 47460 45166
rect 47740 45052 47796 45108
rect 47404 43426 47460 43428
rect 47404 43374 47406 43426
rect 47406 43374 47458 43426
rect 47458 43374 47460 43426
rect 47404 43372 47460 43374
rect 47516 41916 47572 41972
rect 47068 40402 47124 40404
rect 47068 40350 47070 40402
rect 47070 40350 47122 40402
rect 47122 40350 47124 40402
rect 47068 40348 47124 40350
rect 47404 39116 47460 39172
rect 46956 38332 47012 38388
rect 46844 37938 46900 37940
rect 46844 37886 46846 37938
rect 46846 37886 46898 37938
rect 46898 37886 46900 37938
rect 46844 37884 46900 37886
rect 46732 37826 46788 37828
rect 46732 37774 46734 37826
rect 46734 37774 46786 37826
rect 46786 37774 46788 37826
rect 46732 37772 46788 37774
rect 46396 35868 46452 35924
rect 45276 34636 45332 34692
rect 45164 31836 45220 31892
rect 45724 34748 45780 34804
rect 46172 33234 46228 33236
rect 46172 33182 46174 33234
rect 46174 33182 46226 33234
rect 46226 33182 46228 33234
rect 46172 33180 46228 33182
rect 45836 31836 45892 31892
rect 45276 31724 45332 31780
rect 45612 31666 45668 31668
rect 45612 31614 45614 31666
rect 45614 31614 45666 31666
rect 45666 31614 45668 31666
rect 45612 31612 45668 31614
rect 45612 31388 45668 31444
rect 45052 30994 45108 30996
rect 45052 30942 45054 30994
rect 45054 30942 45106 30994
rect 45106 30942 45108 30994
rect 45052 30940 45108 30942
rect 44940 30156 44996 30212
rect 45164 30268 45220 30324
rect 45836 30940 45892 30996
rect 45612 30210 45668 30212
rect 45612 30158 45614 30210
rect 45614 30158 45666 30210
rect 45666 30158 45668 30210
rect 45612 30156 45668 30158
rect 45052 29932 45108 29988
rect 44044 28812 44100 28868
rect 43932 28754 43988 28756
rect 43932 28702 43934 28754
rect 43934 28702 43986 28754
rect 43986 28702 43988 28754
rect 43932 28700 43988 28702
rect 43484 24444 43540 24500
rect 43148 23772 43204 23828
rect 42700 23548 42756 23604
rect 42812 23660 42868 23716
rect 42252 22482 42308 22484
rect 42252 22430 42254 22482
rect 42254 22430 42306 22482
rect 42306 22430 42308 22482
rect 42252 22428 42308 22430
rect 42252 22092 42308 22148
rect 41692 20636 41748 20692
rect 40908 16882 40964 16884
rect 40908 16830 40910 16882
rect 40910 16830 40962 16882
rect 40962 16830 40964 16882
rect 40908 16828 40964 16830
rect 41020 15372 41076 15428
rect 41132 18396 41188 18452
rect 43148 22764 43204 22820
rect 43372 22540 43428 22596
rect 41580 18284 41636 18340
rect 42028 18338 42084 18340
rect 42028 18286 42030 18338
rect 42030 18286 42082 18338
rect 42082 18286 42084 18338
rect 42028 18284 42084 18286
rect 41916 17666 41972 17668
rect 41916 17614 41918 17666
rect 41918 17614 41970 17666
rect 41970 17614 41972 17666
rect 41916 17612 41972 17614
rect 42812 21308 42868 21364
rect 42700 17948 42756 18004
rect 42924 18956 42980 19012
rect 44492 29260 44548 29316
rect 44492 28028 44548 28084
rect 44268 27186 44324 27188
rect 44268 27134 44270 27186
rect 44270 27134 44322 27186
rect 44322 27134 44324 27186
rect 44268 27132 44324 27134
rect 44716 28812 44772 28868
rect 44940 28642 44996 28644
rect 44940 28590 44942 28642
rect 44942 28590 44994 28642
rect 44994 28590 44996 28642
rect 44940 28588 44996 28590
rect 45388 29484 45444 29540
rect 46620 33068 46676 33124
rect 46732 33292 46788 33348
rect 46172 31500 46228 31556
rect 47404 38108 47460 38164
rect 47628 40348 47684 40404
rect 48076 44210 48132 44212
rect 48076 44158 48078 44210
rect 48078 44158 48130 44210
rect 48130 44158 48132 44210
rect 48076 44156 48132 44158
rect 47964 41804 48020 41860
rect 48188 42642 48244 42644
rect 48188 42590 48190 42642
rect 48190 42590 48242 42642
rect 48242 42590 48244 42642
rect 48188 42588 48244 42590
rect 48412 42588 48468 42644
rect 47852 40514 47908 40516
rect 47852 40462 47854 40514
rect 47854 40462 47906 40514
rect 47906 40462 47908 40514
rect 47852 40460 47908 40462
rect 47628 38050 47684 38052
rect 47628 37998 47630 38050
rect 47630 37998 47682 38050
rect 47682 37998 47684 38050
rect 47628 37996 47684 37998
rect 47404 36876 47460 36932
rect 47740 37436 47796 37492
rect 47740 36988 47796 37044
rect 48076 37660 48132 37716
rect 48300 37212 48356 37268
rect 48188 35586 48244 35588
rect 48188 35534 48190 35586
rect 48190 35534 48242 35586
rect 48242 35534 48244 35586
rect 48188 35532 48244 35534
rect 47180 34972 47236 35028
rect 48188 35026 48244 35028
rect 48188 34974 48190 35026
rect 48190 34974 48242 35026
rect 48242 34974 48244 35026
rect 48188 34972 48244 34974
rect 47852 34636 47908 34692
rect 46172 30940 46228 30996
rect 46060 30156 46116 30212
rect 45836 29372 45892 29428
rect 46060 29484 46116 29540
rect 46396 31106 46452 31108
rect 46396 31054 46398 31106
rect 46398 31054 46450 31106
rect 46450 31054 46452 31106
rect 46396 31052 46452 31054
rect 46620 31388 46676 31444
rect 46396 30434 46452 30436
rect 46396 30382 46398 30434
rect 46398 30382 46450 30434
rect 46450 30382 46452 30434
rect 46396 30380 46452 30382
rect 46508 30268 46564 30324
rect 47852 33346 47908 33348
rect 47852 33294 47854 33346
rect 47854 33294 47906 33346
rect 47906 33294 47908 33346
rect 47852 33292 47908 33294
rect 47516 33234 47572 33236
rect 47516 33182 47518 33234
rect 47518 33182 47570 33234
rect 47570 33182 47572 33234
rect 47516 33180 47572 33182
rect 47180 33068 47236 33124
rect 48076 32284 48132 32340
rect 47404 31106 47460 31108
rect 47404 31054 47406 31106
rect 47406 31054 47458 31106
rect 47458 31054 47460 31106
rect 47404 31052 47460 31054
rect 46956 30716 47012 30772
rect 47628 30604 47684 30660
rect 47628 30380 47684 30436
rect 47068 30210 47124 30212
rect 47068 30158 47070 30210
rect 47070 30158 47122 30210
rect 47122 30158 47124 30210
rect 47068 30156 47124 30158
rect 46284 29484 46340 29540
rect 46620 29484 46676 29540
rect 47068 29426 47124 29428
rect 47068 29374 47070 29426
rect 47070 29374 47122 29426
rect 47122 29374 47124 29426
rect 47068 29372 47124 29374
rect 46172 28812 46228 28868
rect 45276 27580 45332 27636
rect 44380 23772 44436 23828
rect 45052 26348 45108 26404
rect 44940 25564 44996 25620
rect 45052 25506 45108 25508
rect 45052 25454 45054 25506
rect 45054 25454 45106 25506
rect 45106 25454 45108 25506
rect 45052 25452 45108 25454
rect 45276 25340 45332 25396
rect 48076 29986 48132 29988
rect 48076 29934 48078 29986
rect 48078 29934 48130 29986
rect 48130 29934 48132 29986
rect 48076 29932 48132 29934
rect 45836 27858 45892 27860
rect 45836 27806 45838 27858
rect 45838 27806 45890 27858
rect 45890 27806 45892 27858
rect 45836 27804 45892 27806
rect 45500 27634 45556 27636
rect 45500 27582 45502 27634
rect 45502 27582 45554 27634
rect 45554 27582 45556 27634
rect 45500 27580 45556 27582
rect 45164 24668 45220 24724
rect 45052 24050 45108 24052
rect 45052 23998 45054 24050
rect 45054 23998 45106 24050
rect 45106 23998 45108 24050
rect 45052 23996 45108 23998
rect 44828 23660 44884 23716
rect 44940 23266 44996 23268
rect 44940 23214 44942 23266
rect 44942 23214 44994 23266
rect 44994 23214 44996 23266
rect 44940 23212 44996 23214
rect 44156 23100 44212 23156
rect 45500 27356 45556 27412
rect 45836 26684 45892 26740
rect 45612 26402 45668 26404
rect 45612 26350 45614 26402
rect 45614 26350 45666 26402
rect 45666 26350 45668 26402
rect 45612 26348 45668 26350
rect 45836 26236 45892 26292
rect 46396 26684 46452 26740
rect 46508 27132 46564 27188
rect 47516 27804 47572 27860
rect 47068 27634 47124 27636
rect 47068 27582 47070 27634
rect 47070 27582 47122 27634
rect 47122 27582 47124 27634
rect 47068 27580 47124 27582
rect 47068 27132 47124 27188
rect 48188 29314 48244 29316
rect 48188 29262 48190 29314
rect 48190 29262 48242 29314
rect 48242 29262 48244 29314
rect 48188 29260 48244 29262
rect 47852 27356 47908 27412
rect 48188 27356 48244 27412
rect 48188 27186 48244 27188
rect 48188 27134 48190 27186
rect 48190 27134 48242 27186
rect 48242 27134 48244 27186
rect 48188 27132 48244 27134
rect 45836 25676 45892 25732
rect 46508 25676 46564 25732
rect 46060 25228 46116 25284
rect 45948 24722 46004 24724
rect 45948 24670 45950 24722
rect 45950 24670 46002 24722
rect 46002 24670 46004 24722
rect 45948 24668 46004 24670
rect 45612 24498 45668 24500
rect 45612 24446 45614 24498
rect 45614 24446 45666 24498
rect 45666 24446 45668 24498
rect 45612 24444 45668 24446
rect 47404 25788 47460 25844
rect 46732 25116 46788 25172
rect 47628 25788 47684 25844
rect 47516 25564 47572 25620
rect 47404 25506 47460 25508
rect 47404 25454 47406 25506
rect 47406 25454 47458 25506
rect 47458 25454 47460 25506
rect 47404 25452 47460 25454
rect 47180 25340 47236 25396
rect 47292 25282 47348 25284
rect 47292 25230 47294 25282
rect 47294 25230 47346 25282
rect 47346 25230 47348 25282
rect 47292 25228 47348 25230
rect 47628 25116 47684 25172
rect 45276 23100 45332 23156
rect 44268 23042 44324 23044
rect 44268 22990 44270 23042
rect 44270 22990 44322 23042
rect 44322 22990 44324 23042
rect 44268 22988 44324 22990
rect 43820 22764 43876 22820
rect 44156 22540 44212 22596
rect 44044 22146 44100 22148
rect 44044 22094 44046 22146
rect 44046 22094 44098 22146
rect 44098 22094 44100 22146
rect 44044 22092 44100 22094
rect 44044 21420 44100 21476
rect 43932 21308 43988 21364
rect 43932 19964 43988 20020
rect 43708 19346 43764 19348
rect 43708 19294 43710 19346
rect 43710 19294 43762 19346
rect 43762 19294 43764 19346
rect 43708 19292 43764 19294
rect 43036 18284 43092 18340
rect 43036 17724 43092 17780
rect 42028 16828 42084 16884
rect 41244 15708 41300 15764
rect 43148 17500 43204 17556
rect 43036 16492 43092 16548
rect 42924 16098 42980 16100
rect 42924 16046 42926 16098
rect 42926 16046 42978 16098
rect 42978 16046 42980 16098
rect 42924 16044 42980 16046
rect 41916 15874 41972 15876
rect 41916 15822 41918 15874
rect 41918 15822 41970 15874
rect 41970 15822 41972 15874
rect 41916 15820 41972 15822
rect 42476 15820 42532 15876
rect 41692 15372 41748 15428
rect 42812 15314 42868 15316
rect 42812 15262 42814 15314
rect 42814 15262 42866 15314
rect 42866 15262 42868 15314
rect 42812 15260 42868 15262
rect 42140 15202 42196 15204
rect 42140 15150 42142 15202
rect 42142 15150 42194 15202
rect 42194 15150 42196 15202
rect 42140 15148 42196 15150
rect 40908 14476 40964 14532
rect 40908 14306 40964 14308
rect 40908 14254 40910 14306
rect 40910 14254 40962 14306
rect 40962 14254 40964 14306
rect 40908 14252 40964 14254
rect 40572 14028 40628 14084
rect 41020 14028 41076 14084
rect 40908 13468 40964 13524
rect 41020 13244 41076 13300
rect 40684 13074 40740 13076
rect 40684 13022 40686 13074
rect 40686 13022 40738 13074
rect 40738 13022 40740 13074
rect 40684 13020 40740 13022
rect 40460 12908 40516 12964
rect 40348 12572 40404 12628
rect 41692 13020 41748 13076
rect 41468 12572 41524 12628
rect 41132 12066 41188 12068
rect 41132 12014 41134 12066
rect 41134 12014 41186 12066
rect 41186 12014 41188 12066
rect 41132 12012 41188 12014
rect 39676 10444 39732 10500
rect 40572 11676 40628 11732
rect 41132 11676 41188 11732
rect 42812 13356 42868 13412
rect 42812 12908 42868 12964
rect 43148 15484 43204 15540
rect 43148 15148 43204 15204
rect 43820 18450 43876 18452
rect 43820 18398 43822 18450
rect 43822 18398 43874 18450
rect 43874 18398 43876 18450
rect 43820 18396 43876 18398
rect 44380 20914 44436 20916
rect 44380 20862 44382 20914
rect 44382 20862 44434 20914
rect 44434 20862 44436 20914
rect 44380 20860 44436 20862
rect 46396 23212 46452 23268
rect 47180 23266 47236 23268
rect 47180 23214 47182 23266
rect 47182 23214 47234 23266
rect 47234 23214 47236 23266
rect 47180 23212 47236 23214
rect 46732 23154 46788 23156
rect 46732 23102 46734 23154
rect 46734 23102 46786 23154
rect 46786 23102 46788 23154
rect 46732 23100 46788 23102
rect 45724 22540 45780 22596
rect 45276 21196 45332 21252
rect 45388 21532 45444 21588
rect 45948 22764 46004 22820
rect 47516 23212 47572 23268
rect 47404 23042 47460 23044
rect 47404 22990 47406 23042
rect 47406 22990 47458 23042
rect 47458 22990 47460 23042
rect 47404 22988 47460 22990
rect 46620 22316 46676 22372
rect 46396 21644 46452 21700
rect 47180 22370 47236 22372
rect 47180 22318 47182 22370
rect 47182 22318 47234 22370
rect 47234 22318 47236 22370
rect 47180 22316 47236 22318
rect 47964 24722 48020 24724
rect 47964 24670 47966 24722
rect 47966 24670 48018 24722
rect 48018 24670 48020 24722
rect 47964 24668 48020 24670
rect 47964 23996 48020 24052
rect 48188 25788 48244 25844
rect 48412 24668 48468 24724
rect 47852 23212 47908 23268
rect 45052 20188 45108 20244
rect 45052 20018 45108 20020
rect 45052 19966 45054 20018
rect 45054 19966 45106 20018
rect 45106 19966 45108 20018
rect 45052 19964 45108 19966
rect 44604 19906 44660 19908
rect 44604 19854 44606 19906
rect 44606 19854 44658 19906
rect 44658 19854 44660 19906
rect 44604 19852 44660 19854
rect 45276 19852 45332 19908
rect 44604 19292 44660 19348
rect 45052 18844 45108 18900
rect 43372 17500 43428 17556
rect 43596 17612 43652 17668
rect 44044 17778 44100 17780
rect 44044 17726 44046 17778
rect 44046 17726 44098 17778
rect 44098 17726 44100 17778
rect 44044 17724 44100 17726
rect 45500 18562 45556 18564
rect 45500 18510 45502 18562
rect 45502 18510 45554 18562
rect 45554 18510 45556 18562
rect 45500 18508 45556 18510
rect 44716 17666 44772 17668
rect 44716 17614 44718 17666
rect 44718 17614 44770 17666
rect 44770 17614 44772 17666
rect 44716 17612 44772 17614
rect 43932 16716 43988 16772
rect 44156 16882 44212 16884
rect 44156 16830 44158 16882
rect 44158 16830 44210 16882
rect 44210 16830 44212 16882
rect 44156 16828 44212 16830
rect 43708 16044 43764 16100
rect 44044 16044 44100 16100
rect 43484 15538 43540 15540
rect 43484 15486 43486 15538
rect 43486 15486 43538 15538
rect 43538 15486 43540 15538
rect 43484 15484 43540 15486
rect 43932 15538 43988 15540
rect 43932 15486 43934 15538
rect 43934 15486 43986 15538
rect 43986 15486 43988 15538
rect 43932 15484 43988 15486
rect 43708 14476 43764 14532
rect 43260 13916 43316 13972
rect 43148 13074 43204 13076
rect 43148 13022 43150 13074
rect 43150 13022 43202 13074
rect 43202 13022 43204 13074
rect 43148 13020 43204 13022
rect 43036 12796 43092 12852
rect 42364 12066 42420 12068
rect 42364 12014 42366 12066
rect 42366 12014 42418 12066
rect 42418 12014 42420 12066
rect 42364 12012 42420 12014
rect 41468 11506 41524 11508
rect 41468 11454 41470 11506
rect 41470 11454 41522 11506
rect 41522 11454 41524 11506
rect 41468 11452 41524 11454
rect 42364 11452 42420 11508
rect 40236 11394 40292 11396
rect 40236 11342 40238 11394
rect 40238 11342 40290 11394
rect 40290 11342 40292 11394
rect 40236 11340 40292 11342
rect 41132 11394 41188 11396
rect 41132 11342 41134 11394
rect 41134 11342 41186 11394
rect 41186 11342 41188 11394
rect 41132 11340 41188 11342
rect 42028 11394 42084 11396
rect 42028 11342 42030 11394
rect 42030 11342 42082 11394
rect 42082 11342 42084 11394
rect 42028 11340 42084 11342
rect 41020 11228 41076 11284
rect 40012 10610 40068 10612
rect 40012 10558 40014 10610
rect 40014 10558 40066 10610
rect 40066 10558 40068 10610
rect 40012 10556 40068 10558
rect 40124 9884 40180 9940
rect 38444 8316 38500 8372
rect 39340 9212 39396 9268
rect 39900 9212 39956 9268
rect 38668 8034 38724 8036
rect 38668 7982 38670 8034
rect 38670 7982 38722 8034
rect 38722 7982 38724 8034
rect 38668 7980 38724 7982
rect 38556 7868 38612 7924
rect 38108 7474 38164 7476
rect 38108 7422 38110 7474
rect 38110 7422 38162 7474
rect 38162 7422 38164 7474
rect 38108 7420 38164 7422
rect 37884 7308 37940 7364
rect 37212 6860 37268 6916
rect 37772 7250 37828 7252
rect 37772 7198 37774 7250
rect 37774 7198 37826 7250
rect 37826 7198 37828 7250
rect 37772 7196 37828 7198
rect 35980 6076 36036 6132
rect 34972 5628 35028 5684
rect 34636 5234 34692 5236
rect 34636 5182 34638 5234
rect 34638 5182 34690 5234
rect 34690 5182 34692 5234
rect 34636 5180 34692 5182
rect 34748 5122 34804 5124
rect 34748 5070 34750 5122
rect 34750 5070 34802 5122
rect 34802 5070 34804 5122
rect 34748 5068 34804 5070
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35868 5682 35924 5684
rect 35868 5630 35870 5682
rect 35870 5630 35922 5682
rect 35922 5630 35924 5682
rect 35868 5628 35924 5630
rect 36204 6188 36260 6244
rect 36428 6076 36484 6132
rect 37212 6130 37268 6132
rect 37212 6078 37214 6130
rect 37214 6078 37266 6130
rect 37266 6078 37268 6130
rect 37212 6076 37268 6078
rect 36764 5516 36820 5572
rect 35980 4956 36036 5012
rect 34860 4396 34916 4452
rect 36092 4898 36148 4900
rect 36092 4846 36094 4898
rect 36094 4846 36146 4898
rect 36146 4846 36148 4898
rect 36092 4844 36148 4846
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 36316 4226 36372 4228
rect 36316 4174 36318 4226
rect 36318 4174 36370 4226
rect 36370 4174 36372 4226
rect 36316 4172 36372 4174
rect 37772 6748 37828 6804
rect 37436 6466 37492 6468
rect 37436 6414 37438 6466
rect 37438 6414 37490 6466
rect 37490 6414 37492 6466
rect 37436 6412 37492 6414
rect 37324 5516 37380 5572
rect 37212 4956 37268 5012
rect 38332 7362 38388 7364
rect 38332 7310 38334 7362
rect 38334 7310 38386 7362
rect 38386 7310 38388 7362
rect 38332 7308 38388 7310
rect 38220 7196 38276 7252
rect 38108 6914 38164 6916
rect 38108 6862 38110 6914
rect 38110 6862 38162 6914
rect 38162 6862 38164 6914
rect 38108 6860 38164 6862
rect 38892 7698 38948 7700
rect 38892 7646 38894 7698
rect 38894 7646 38946 7698
rect 38946 7646 38948 7698
rect 38892 7644 38948 7646
rect 38668 7474 38724 7476
rect 38668 7422 38670 7474
rect 38670 7422 38722 7474
rect 38722 7422 38724 7474
rect 38668 7420 38724 7422
rect 38892 7308 38948 7364
rect 39788 7980 39844 8036
rect 39676 7868 39732 7924
rect 39228 7644 39284 7700
rect 39116 7586 39172 7588
rect 39116 7534 39118 7586
rect 39118 7534 39170 7586
rect 39170 7534 39172 7586
rect 39116 7532 39172 7534
rect 38780 6860 38836 6916
rect 39340 6972 39396 7028
rect 38892 6748 38948 6804
rect 38556 6578 38612 6580
rect 38556 6526 38558 6578
rect 38558 6526 38610 6578
rect 38610 6526 38612 6578
rect 38556 6524 38612 6526
rect 38780 5516 38836 5572
rect 38444 4844 38500 4900
rect 39004 5404 39060 5460
rect 39564 6412 39620 6468
rect 40012 8092 40068 8148
rect 40124 8316 40180 8372
rect 40908 10444 40964 10500
rect 40348 9772 40404 9828
rect 41692 9996 41748 10052
rect 43932 14476 43988 14532
rect 43484 11788 43540 11844
rect 43036 11506 43092 11508
rect 43036 11454 43038 11506
rect 43038 11454 43090 11506
rect 43090 11454 43092 11506
rect 43036 11452 43092 11454
rect 43484 11506 43540 11508
rect 43484 11454 43486 11506
rect 43486 11454 43538 11506
rect 43538 11454 43540 11506
rect 43484 11452 43540 11454
rect 42476 9996 42532 10052
rect 41020 9714 41076 9716
rect 41020 9662 41022 9714
rect 41022 9662 41074 9714
rect 41074 9662 41076 9714
rect 41020 9660 41076 9662
rect 40460 9100 40516 9156
rect 39788 7420 39844 7476
rect 40236 8034 40292 8036
rect 40236 7982 40238 8034
rect 40238 7982 40290 8034
rect 40290 7982 40292 8034
rect 40236 7980 40292 7982
rect 40236 7698 40292 7700
rect 40236 7646 40238 7698
rect 40238 7646 40290 7698
rect 40290 7646 40292 7698
rect 40236 7644 40292 7646
rect 40348 7532 40404 7588
rect 40796 8316 40852 8372
rect 41020 8258 41076 8260
rect 41020 8206 41022 8258
rect 41022 8206 41074 8258
rect 41074 8206 41076 8258
rect 41020 8204 41076 8206
rect 41020 7868 41076 7924
rect 41916 9772 41972 9828
rect 41244 8204 41300 8260
rect 41356 8428 41412 8484
rect 42476 8876 42532 8932
rect 42252 8316 42308 8372
rect 40908 7644 40964 7700
rect 41244 7644 41300 7700
rect 40124 7084 40180 7140
rect 40124 6748 40180 6804
rect 39788 6578 39844 6580
rect 39788 6526 39790 6578
rect 39790 6526 39842 6578
rect 39842 6526 39844 6578
rect 39788 6524 39844 6526
rect 40236 6466 40292 6468
rect 40236 6414 40238 6466
rect 40238 6414 40290 6466
rect 40290 6414 40292 6466
rect 40236 6412 40292 6414
rect 40348 6188 40404 6244
rect 40908 6300 40964 6356
rect 41020 5964 41076 6020
rect 40908 5740 40964 5796
rect 38892 5010 38948 5012
rect 38892 4958 38894 5010
rect 38894 4958 38946 5010
rect 38946 4958 38948 5010
rect 38892 4956 38948 4958
rect 39116 4508 39172 4564
rect 39788 5404 39844 5460
rect 39676 4114 39732 4116
rect 39676 4062 39678 4114
rect 39678 4062 39730 4114
rect 39730 4062 39732 4114
rect 39676 4060 39732 4062
rect 40124 4562 40180 4564
rect 40124 4510 40126 4562
rect 40126 4510 40178 4562
rect 40178 4510 40180 4562
rect 40124 4508 40180 4510
rect 41020 4508 41076 4564
rect 41244 7084 41300 7140
rect 41580 7644 41636 7700
rect 41468 6972 41524 7028
rect 41916 7980 41972 8036
rect 41804 7474 41860 7476
rect 41804 7422 41806 7474
rect 41806 7422 41858 7474
rect 41858 7422 41860 7474
rect 41804 7420 41860 7422
rect 42140 8258 42196 8260
rect 42140 8206 42142 8258
rect 42142 8206 42194 8258
rect 42194 8206 42196 8258
rect 42140 8204 42196 8206
rect 43148 10722 43204 10724
rect 43148 10670 43150 10722
rect 43150 10670 43202 10722
rect 43202 10670 43204 10722
rect 43148 10668 43204 10670
rect 42812 10050 42868 10052
rect 42812 9998 42814 10050
rect 42814 9998 42866 10050
rect 42866 9998 42868 10050
rect 42812 9996 42868 9998
rect 43036 9826 43092 9828
rect 43036 9774 43038 9826
rect 43038 9774 43090 9826
rect 43090 9774 43092 9826
rect 43036 9772 43092 9774
rect 43484 9212 43540 9268
rect 43260 9100 43316 9156
rect 42812 8540 42868 8596
rect 42812 8258 42868 8260
rect 42812 8206 42814 8258
rect 42814 8206 42866 8258
rect 42866 8206 42868 8258
rect 42812 8204 42868 8206
rect 43148 8146 43204 8148
rect 43148 8094 43150 8146
rect 43150 8094 43202 8146
rect 43202 8094 43204 8146
rect 43148 8092 43204 8094
rect 43260 8034 43316 8036
rect 43260 7982 43262 8034
rect 43262 7982 43314 8034
rect 43314 7982 43316 8034
rect 43260 7980 43316 7982
rect 42812 7868 42868 7924
rect 43372 7868 43428 7924
rect 45164 17554 45220 17556
rect 45164 17502 45166 17554
rect 45166 17502 45218 17554
rect 45218 17502 45220 17554
rect 45164 17500 45220 17502
rect 46396 20242 46452 20244
rect 46396 20190 46398 20242
rect 46398 20190 46450 20242
rect 46450 20190 46452 20242
rect 46396 20188 46452 20190
rect 45836 19964 45892 20020
rect 47180 21644 47236 21700
rect 47852 21698 47908 21700
rect 47852 21646 47854 21698
rect 47854 21646 47906 21698
rect 47906 21646 47908 21698
rect 47852 21644 47908 21646
rect 47068 21474 47124 21476
rect 47068 21422 47070 21474
rect 47070 21422 47122 21474
rect 47122 21422 47124 21474
rect 47068 21420 47124 21422
rect 48076 22988 48132 23044
rect 48076 22204 48132 22260
rect 48076 20860 48132 20916
rect 46844 20018 46900 20020
rect 46844 19966 46846 20018
rect 46846 19966 46898 20018
rect 46898 19966 46900 20018
rect 46844 19964 46900 19966
rect 47068 19740 47124 19796
rect 45836 18508 45892 18564
rect 45948 18284 46004 18340
rect 45388 17666 45444 17668
rect 45388 17614 45390 17666
rect 45390 17614 45442 17666
rect 45442 17614 45444 17666
rect 45388 17612 45444 17614
rect 45612 17554 45668 17556
rect 45612 17502 45614 17554
rect 45614 17502 45666 17554
rect 45666 17502 45668 17554
rect 45612 17500 45668 17502
rect 45276 16828 45332 16884
rect 45052 16044 45108 16100
rect 44380 15260 44436 15316
rect 44716 15260 44772 15316
rect 44268 14476 44324 14532
rect 43820 12962 43876 12964
rect 43820 12910 43822 12962
rect 43822 12910 43874 12962
rect 43874 12910 43876 12962
rect 43820 12908 43876 12910
rect 44156 12402 44212 12404
rect 44156 12350 44158 12402
rect 44158 12350 44210 12402
rect 44210 12350 44212 12402
rect 44156 12348 44212 12350
rect 45388 15260 45444 15316
rect 45500 15148 45556 15204
rect 44380 11788 44436 11844
rect 43820 8930 43876 8932
rect 43820 8878 43822 8930
rect 43822 8878 43874 8930
rect 43874 8878 43876 8930
rect 43820 8876 43876 8878
rect 43820 7980 43876 8036
rect 44268 11004 44324 11060
rect 44156 8258 44212 8260
rect 44156 8206 44158 8258
rect 44158 8206 44210 8258
rect 44210 8206 44212 8258
rect 44156 8204 44212 8206
rect 44156 7644 44212 7700
rect 42476 7532 42532 7588
rect 41692 6412 41748 6468
rect 41356 5964 41412 6020
rect 43708 7474 43764 7476
rect 43708 7422 43710 7474
rect 43710 7422 43762 7474
rect 43762 7422 43764 7474
rect 43708 7420 43764 7422
rect 43260 6972 43316 7028
rect 42140 6578 42196 6580
rect 42140 6526 42142 6578
rect 42142 6526 42194 6578
rect 42194 6526 42196 6578
rect 42140 6524 42196 6526
rect 42476 6412 42532 6468
rect 42140 6188 42196 6244
rect 44492 9548 44548 9604
rect 45836 16716 45892 16772
rect 46956 19292 47012 19348
rect 46284 17554 46340 17556
rect 46284 17502 46286 17554
rect 46286 17502 46338 17554
rect 46338 17502 46340 17554
rect 46284 17500 46340 17502
rect 46060 16828 46116 16884
rect 45948 15372 46004 15428
rect 45836 15148 45892 15204
rect 47180 18284 47236 18340
rect 47068 17554 47124 17556
rect 47068 17502 47070 17554
rect 47070 17502 47122 17554
rect 47122 17502 47124 17554
rect 47068 17500 47124 17502
rect 47516 17554 47572 17556
rect 47516 17502 47518 17554
rect 47518 17502 47570 17554
rect 47570 17502 47572 17554
rect 47516 17500 47572 17502
rect 46396 16716 46452 16772
rect 46956 16492 47012 16548
rect 47516 16882 47572 16884
rect 47516 16830 47518 16882
rect 47518 16830 47570 16882
rect 47570 16830 47572 16882
rect 47516 16828 47572 16830
rect 47740 20018 47796 20020
rect 47740 19966 47742 20018
rect 47742 19966 47794 20018
rect 47794 19966 47796 20018
rect 47740 19964 47796 19966
rect 47852 19794 47908 19796
rect 47852 19742 47854 19794
rect 47854 19742 47906 19794
rect 47906 19742 47908 19794
rect 47852 19740 47908 19742
rect 48188 19346 48244 19348
rect 48188 19294 48190 19346
rect 48190 19294 48242 19346
rect 48242 19294 48244 19346
rect 48188 19292 48244 19294
rect 48076 18450 48132 18452
rect 48076 18398 48078 18450
rect 48078 18398 48130 18450
rect 48130 18398 48132 18450
rect 48076 18396 48132 18398
rect 47964 18284 48020 18340
rect 48076 17500 48132 17556
rect 47628 16492 47684 16548
rect 47404 15426 47460 15428
rect 47404 15374 47406 15426
rect 47406 15374 47458 15426
rect 47458 15374 47460 15426
rect 47404 15372 47460 15374
rect 46284 15260 46340 15316
rect 46844 15314 46900 15316
rect 46844 15262 46846 15314
rect 46846 15262 46898 15314
rect 46898 15262 46900 15314
rect 46844 15260 46900 15262
rect 47964 15314 48020 15316
rect 47964 15262 47966 15314
rect 47966 15262 48018 15314
rect 48018 15262 48020 15314
rect 47964 15260 48020 15262
rect 45612 14700 45668 14756
rect 46060 14418 46116 14420
rect 46060 14366 46062 14418
rect 46062 14366 46114 14418
rect 46114 14366 46116 14418
rect 46060 14364 46116 14366
rect 44940 12402 44996 12404
rect 44940 12350 44942 12402
rect 44942 12350 44994 12402
rect 44994 12350 44996 12402
rect 44940 12348 44996 12350
rect 44940 11282 44996 11284
rect 44940 11230 44942 11282
rect 44942 11230 44994 11282
rect 44994 11230 44996 11282
rect 44940 11228 44996 11230
rect 44828 11004 44884 11060
rect 45276 12348 45332 12404
rect 45164 11340 45220 11396
rect 45724 11564 45780 11620
rect 46956 14364 47012 14420
rect 46956 13746 47012 13748
rect 46956 13694 46958 13746
rect 46958 13694 47010 13746
rect 47010 13694 47012 13746
rect 46956 13692 47012 13694
rect 46284 12572 46340 12628
rect 46844 12460 46900 12516
rect 45948 12012 46004 12068
rect 46732 12124 46788 12180
rect 45276 11228 45332 11284
rect 45164 11170 45220 11172
rect 45164 11118 45166 11170
rect 45166 11118 45218 11170
rect 45218 11118 45220 11170
rect 45164 11116 45220 11118
rect 45500 10668 45556 10724
rect 46060 11116 46116 11172
rect 46396 11618 46452 11620
rect 46396 11566 46398 11618
rect 46398 11566 46450 11618
rect 46450 11566 46452 11618
rect 46396 11564 46452 11566
rect 46508 11394 46564 11396
rect 46508 11342 46510 11394
rect 46510 11342 46562 11394
rect 46562 11342 46564 11394
rect 46508 11340 46564 11342
rect 46396 11282 46452 11284
rect 46396 11230 46398 11282
rect 46398 11230 46450 11282
rect 46450 11230 46452 11282
rect 46396 11228 46452 11230
rect 46844 11282 46900 11284
rect 46844 11230 46846 11282
rect 46846 11230 46898 11282
rect 46898 11230 46900 11282
rect 46844 11228 46900 11230
rect 47628 12572 47684 12628
rect 47516 12012 47572 12068
rect 47852 13746 47908 13748
rect 47852 13694 47854 13746
rect 47854 13694 47906 13746
rect 47906 13694 47908 13746
rect 47852 13692 47908 13694
rect 47852 12850 47908 12852
rect 47852 12798 47854 12850
rect 47854 12798 47906 12850
rect 47906 12798 47908 12850
rect 47852 12796 47908 12798
rect 48188 12572 48244 12628
rect 47852 12124 47908 12180
rect 48188 12066 48244 12068
rect 48188 12014 48190 12066
rect 48190 12014 48242 12066
rect 48242 12014 48244 12066
rect 48188 12012 48244 12014
rect 48300 11452 48356 11508
rect 47628 11394 47684 11396
rect 47628 11342 47630 11394
rect 47630 11342 47682 11394
rect 47682 11342 47684 11394
rect 47628 11340 47684 11342
rect 46956 10556 47012 10612
rect 44940 9602 44996 9604
rect 44940 9550 44942 9602
rect 44942 9550 44994 9602
rect 44994 9550 44996 9602
rect 44940 9548 44996 9550
rect 44492 8204 44548 8260
rect 44940 8034 44996 8036
rect 44940 7982 44942 8034
rect 44942 7982 44994 8034
rect 44994 7982 44996 8034
rect 44940 7980 44996 7982
rect 45052 7698 45108 7700
rect 45052 7646 45054 7698
rect 45054 7646 45106 7698
rect 45106 7646 45108 7698
rect 45052 7644 45108 7646
rect 44492 7532 44548 7588
rect 43708 6300 43764 6356
rect 44380 6412 44436 6468
rect 44940 6578 44996 6580
rect 44940 6526 44942 6578
rect 44942 6526 44994 6578
rect 44994 6526 44996 6578
rect 44940 6524 44996 6526
rect 45388 8258 45444 8260
rect 45388 8206 45390 8258
rect 45390 8206 45442 8258
rect 45442 8206 45444 8258
rect 45388 8204 45444 8206
rect 47852 9042 47908 9044
rect 47852 8990 47854 9042
rect 47854 8990 47906 9042
rect 47906 8990 47908 9042
rect 47852 8988 47908 8990
rect 47404 8316 47460 8372
rect 48188 8370 48244 8372
rect 48188 8318 48190 8370
rect 48190 8318 48242 8370
rect 48242 8318 48244 8370
rect 48188 8316 48244 8318
rect 48188 7644 48244 7700
rect 45276 7420 45332 7476
rect 46956 7474 47012 7476
rect 46956 7422 46958 7474
rect 46958 7422 47010 7474
rect 47010 7422 47012 7474
rect 46956 7420 47012 7422
rect 46956 6690 47012 6692
rect 46956 6638 46958 6690
rect 46958 6638 47010 6690
rect 47010 6638 47012 6690
rect 46956 6636 47012 6638
rect 45164 6524 45220 6580
rect 46060 6578 46116 6580
rect 46060 6526 46062 6578
rect 46062 6526 46114 6578
rect 46114 6526 46116 6578
rect 46060 6524 46116 6526
rect 46172 6466 46228 6468
rect 46172 6414 46174 6466
rect 46174 6414 46226 6466
rect 46226 6414 46228 6466
rect 46172 6412 46228 6414
rect 45388 6300 45444 6356
rect 43932 5794 43988 5796
rect 43932 5742 43934 5794
rect 43934 5742 43986 5794
rect 43986 5742 43988 5794
rect 43932 5740 43988 5742
rect 46060 6018 46116 6020
rect 46060 5966 46062 6018
rect 46062 5966 46114 6018
rect 46114 5966 46116 6018
rect 46060 5964 46116 5966
rect 44492 4956 44548 5012
rect 42588 4898 42644 4900
rect 42588 4846 42590 4898
rect 42590 4846 42642 4898
rect 42642 4846 42644 4898
rect 42588 4844 42644 4846
rect 42588 4508 42644 4564
rect 43708 4844 43764 4900
rect 41916 4060 41972 4116
rect 44156 4898 44212 4900
rect 44156 4846 44158 4898
rect 44158 4846 44210 4898
rect 44210 4846 44212 4898
rect 44156 4844 44212 4846
rect 44940 4898 44996 4900
rect 44940 4846 44942 4898
rect 44942 4846 44994 4898
rect 44994 4846 44996 4898
rect 44940 4844 44996 4846
rect 42588 3612 42644 3668
rect 37884 3500 37940 3556
rect 47516 7420 47572 7476
rect 47180 6524 47236 6580
rect 47852 6690 47908 6692
rect 47852 6638 47854 6690
rect 47854 6638 47906 6690
rect 47906 6638 47908 6690
rect 47852 6636 47908 6638
rect 46620 6300 46676 6356
rect 46956 5964 47012 6020
rect 47068 6300 47124 6356
rect 46956 5122 47012 5124
rect 46956 5070 46958 5122
rect 46958 5070 47010 5122
rect 47010 5070 47012 5122
rect 46956 5068 47012 5070
rect 47628 6466 47684 6468
rect 47628 6414 47630 6466
rect 47630 6414 47682 6466
rect 47682 6414 47684 6466
rect 47628 6412 47684 6414
rect 48188 6412 48244 6468
rect 47852 5122 47908 5124
rect 47852 5070 47854 5122
rect 47854 5070 47906 5122
rect 47906 5070 47908 5122
rect 47852 5068 47908 5070
rect 47628 5010 47684 5012
rect 47628 4958 47630 5010
rect 47630 4958 47682 5010
rect 47682 4958 47684 5010
rect 47628 4956 47684 4958
rect 48188 4956 48244 5012
rect 43820 3666 43876 3668
rect 43820 3614 43822 3666
rect 43822 3614 43874 3666
rect 43874 3614 43876 3666
rect 43820 3612 43876 3614
rect 47628 3554 47684 3556
rect 47628 3502 47630 3554
rect 47630 3502 47682 3554
rect 47682 3502 47684 3554
rect 47628 3500 47684 3502
rect 46956 3442 47012 3444
rect 46956 3390 46958 3442
rect 46958 3390 47010 3442
rect 47010 3390 47012 3442
rect 46956 3388 47012 3390
rect 48076 3388 48132 3444
rect 48188 2716 48244 2772
rect 34412 2604 34468 2660
rect 32284 2268 32340 2324
rect 30380 1484 30436 1540
rect 25788 1260 25844 1316
<< metal3 >>
rect 49200 47124 50000 47152
rect 48402 47068 48412 47124
rect 48468 47068 50000 47124
rect 49200 47040 50000 47068
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 20850 46060 20860 46116
rect 20916 46060 22092 46116
rect 22148 46060 22158 46116
rect 22418 46060 22428 46116
rect 22484 46060 25228 46116
rect 25284 46060 25294 46116
rect 33394 46060 33404 46116
rect 33460 46060 36988 46116
rect 37044 46060 37054 46116
rect 38098 46060 38108 46116
rect 38164 46060 40348 46116
rect 40404 46060 40414 46116
rect 41234 46060 41244 46116
rect 41300 46060 44604 46116
rect 44660 46060 44670 46116
rect 35074 45836 35084 45892
rect 35140 45836 35980 45892
rect 36036 45836 36046 45892
rect 13010 45724 13020 45780
rect 13076 45724 13916 45780
rect 13972 45724 13982 45780
rect 14578 45724 14588 45780
rect 14644 45724 16940 45780
rect 16996 45724 17006 45780
rect 44258 45724 44268 45780
rect 44324 45724 46508 45780
rect 46564 45724 46574 45780
rect 5618 45612 5628 45668
rect 5684 45612 9436 45668
rect 9492 45612 9502 45668
rect 11330 45612 11340 45668
rect 11396 45612 13132 45668
rect 13188 45612 13198 45668
rect 42802 45612 42812 45668
rect 42868 45612 44380 45668
rect 44436 45612 44446 45668
rect 45378 45612 45388 45668
rect 45444 45612 47404 45668
rect 47460 45612 47470 45668
rect 13132 45444 13188 45612
rect 43250 45500 43260 45556
rect 43316 45500 46732 45556
rect 46788 45500 46798 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 7970 45388 7980 45444
rect 8036 45388 8540 45444
rect 8596 45388 9548 45444
rect 9604 45388 10892 45444
rect 10948 45388 10958 45444
rect 13132 45388 13524 45444
rect 27122 45388 27132 45444
rect 27188 45388 30996 45444
rect 13468 45332 13524 45388
rect 30940 45332 30996 45388
rect 13468 45276 14028 45332
rect 14084 45276 14094 45332
rect 30930 45276 30940 45332
rect 30996 45276 45276 45332
rect 45332 45276 45342 45332
rect 14028 45108 14084 45276
rect 44818 45164 44828 45220
rect 44884 45164 47404 45220
rect 47460 45164 47470 45220
rect 14028 45052 14588 45108
rect 14644 45052 17500 45108
rect 17556 45052 17566 45108
rect 26338 45052 26348 45108
rect 26404 45052 27468 45108
rect 27524 45052 27534 45108
rect 44930 45052 44940 45108
rect 44996 45052 47740 45108
rect 47796 45052 47806 45108
rect 18610 44940 18620 44996
rect 18676 44940 21308 44996
rect 21364 44940 21374 44996
rect 21858 44940 21868 44996
rect 21924 44940 26124 44996
rect 26180 44940 26190 44996
rect 29922 44940 29932 44996
rect 29988 44940 31388 44996
rect 31444 44940 32172 44996
rect 32228 44940 33180 44996
rect 33236 44940 36428 44996
rect 36484 44940 36494 44996
rect 39218 44828 39228 44884
rect 39284 44828 40012 44884
rect 40068 44828 40078 44884
rect 44146 44828 44156 44884
rect 44212 44828 46844 44884
rect 46900 44828 46910 44884
rect 38770 44716 38780 44772
rect 38836 44716 39340 44772
rect 39396 44716 40348 44772
rect 40404 44716 40414 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 15362 44492 15372 44548
rect 15428 44492 16156 44548
rect 16212 44492 16222 44548
rect 31826 44492 31836 44548
rect 31892 44492 33740 44548
rect 33796 44492 33806 44548
rect 36530 44492 36540 44548
rect 36596 44492 37212 44548
rect 37268 44492 37278 44548
rect 43138 44492 43148 44548
rect 43204 44492 45836 44548
rect 45892 44492 45902 44548
rect 3266 44380 3276 44436
rect 3332 44380 3342 44436
rect 4722 44380 4732 44436
rect 4788 44380 6188 44436
rect 6244 44380 6254 44436
rect 3276 43764 3332 44380
rect 7746 44268 7756 44324
rect 7812 44268 8428 44324
rect 8484 44268 9660 44324
rect 9716 44268 9726 44324
rect 26898 44268 26908 44324
rect 26964 44268 28364 44324
rect 28420 44268 30492 44324
rect 30548 44268 30558 44324
rect 38210 44268 38220 44324
rect 38276 44268 39788 44324
rect 39844 44268 39854 44324
rect 8194 44156 8204 44212
rect 8260 44156 9548 44212
rect 9604 44156 9614 44212
rect 27122 44156 27132 44212
rect 27188 44156 28252 44212
rect 28308 44156 28318 44212
rect 30258 44156 30268 44212
rect 30324 44156 32284 44212
rect 32340 44156 32350 44212
rect 34850 44156 34860 44212
rect 34916 44156 36316 44212
rect 36372 44156 38108 44212
rect 38164 44156 38174 44212
rect 38322 44156 38332 44212
rect 38388 44156 39900 44212
rect 39956 44156 39966 44212
rect 48038 44156 48076 44212
rect 48132 44156 48142 44212
rect 7746 44044 7756 44100
rect 7812 44044 10892 44100
rect 10948 44044 12684 44100
rect 12740 44044 12750 44100
rect 16818 44044 16828 44100
rect 16884 44044 17612 44100
rect 17668 44044 17948 44100
rect 18004 44044 20076 44100
rect 20132 44044 20524 44100
rect 20580 44044 21084 44100
rect 21140 44044 21868 44100
rect 21924 44044 22316 44100
rect 22372 44044 22382 44100
rect 22978 44044 22988 44100
rect 23044 44044 23054 44100
rect 25218 44044 25228 44100
rect 25284 44044 28028 44100
rect 28084 44044 28094 44100
rect 33954 44044 33964 44100
rect 34020 44044 39340 44100
rect 39396 44044 39406 44100
rect 22988 43988 23044 44044
rect 22988 43932 30828 43988
rect 30884 43932 30894 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 12674 43820 12684 43876
rect 12740 43820 13356 43876
rect 13412 43820 13422 43876
rect 27458 43820 27468 43876
rect 27524 43820 28364 43876
rect 28420 43820 28430 43876
rect 37986 43820 37996 43876
rect 38052 43820 38332 43876
rect 38388 43820 38398 43876
rect 43026 43820 43036 43876
rect 43092 43820 44828 43876
rect 44884 43820 44894 43876
rect 3276 43708 3500 43764
rect 3556 43708 3566 43764
rect 7298 43708 7308 43764
rect 7364 43708 8092 43764
rect 8148 43708 8158 43764
rect 13010 43708 13020 43764
rect 13076 43708 13086 43764
rect 28242 43708 28252 43764
rect 28308 43708 29260 43764
rect 29316 43708 29326 43764
rect 31042 43708 31052 43764
rect 31108 43708 32844 43764
rect 32900 43708 32910 43764
rect 38098 43708 38108 43764
rect 38164 43708 43932 43764
rect 43988 43708 43998 43764
rect 13020 43652 13076 43708
rect 39228 43652 39284 43708
rect 3266 43596 3276 43652
rect 3332 43596 4844 43652
rect 4900 43596 4910 43652
rect 12450 43596 12460 43652
rect 12516 43596 13916 43652
rect 13972 43596 13982 43652
rect 14690 43596 14700 43652
rect 14756 43596 15372 43652
rect 15428 43596 15438 43652
rect 24210 43596 24220 43652
rect 24276 43596 25116 43652
rect 25172 43596 25182 43652
rect 25666 43596 25676 43652
rect 25732 43596 26572 43652
rect 26628 43596 26638 43652
rect 30930 43596 30940 43652
rect 30996 43596 32060 43652
rect 32116 43596 32126 43652
rect 34738 43596 34748 43652
rect 34804 43596 35868 43652
rect 35924 43596 38332 43652
rect 38388 43596 38398 43652
rect 39218 43596 39228 43652
rect 39284 43596 39294 43652
rect 45938 43596 45948 43652
rect 46004 43596 47068 43652
rect 47124 43596 47134 43652
rect 14130 43484 14140 43540
rect 14196 43484 15260 43540
rect 15316 43484 16156 43540
rect 16212 43484 16222 43540
rect 21410 43484 21420 43540
rect 21476 43484 24332 43540
rect 24388 43484 24398 43540
rect 24658 43484 24668 43540
rect 24724 43484 25452 43540
rect 25508 43484 25518 43540
rect 29698 43484 29708 43540
rect 29764 43484 31164 43540
rect 31220 43484 31230 43540
rect 37510 43484 37548 43540
rect 37604 43484 37614 43540
rect 40226 43484 40236 43540
rect 40292 43484 42700 43540
rect 42756 43484 44940 43540
rect 44996 43484 45612 43540
rect 45668 43484 45678 43540
rect 5730 43372 5740 43428
rect 5796 43372 6748 43428
rect 6804 43372 6814 43428
rect 14914 43372 14924 43428
rect 14980 43372 16268 43428
rect 16324 43372 16334 43428
rect 18162 43372 18172 43428
rect 18228 43372 20860 43428
rect 20916 43372 20926 43428
rect 22418 43372 22428 43428
rect 22484 43372 23996 43428
rect 24052 43372 24062 43428
rect 32498 43372 32508 43428
rect 32564 43372 37884 43428
rect 37940 43372 38556 43428
rect 38612 43372 38622 43428
rect 39666 43372 39676 43428
rect 39732 43372 41132 43428
rect 41188 43372 41198 43428
rect 43250 43372 43260 43428
rect 43316 43372 47404 43428
rect 47460 43372 47470 43428
rect 1922 43260 1932 43316
rect 1988 43260 3612 43316
rect 3668 43260 4508 43316
rect 4564 43260 4574 43316
rect 15474 43260 15484 43316
rect 15540 43260 16380 43316
rect 16436 43260 16446 43316
rect 16930 43260 16940 43316
rect 16996 43260 23436 43316
rect 23492 43260 23502 43316
rect 34066 43260 34076 43316
rect 34132 43260 38668 43316
rect 38612 43204 38668 43260
rect 9650 43148 9660 43204
rect 9716 43148 10108 43204
rect 10164 43148 10780 43204
rect 10836 43148 28700 43204
rect 28756 43148 28766 43204
rect 38612 43148 40012 43204
rect 40068 43148 45500 43204
rect 45556 43148 45566 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 11778 43036 11788 43092
rect 11844 43036 13580 43092
rect 13636 43036 30828 43092
rect 30884 43036 30894 43092
rect 32050 43036 32060 43092
rect 32116 43036 34076 43092
rect 34132 43036 34142 43092
rect 37538 43036 37548 43092
rect 37604 43036 39004 43092
rect 39060 43036 39070 43092
rect 4834 42924 4844 42980
rect 4900 42924 6300 42980
rect 6356 42924 6366 42980
rect 6626 42924 6636 42980
rect 6692 42924 15708 42980
rect 15764 42924 15774 42980
rect 17938 42924 17948 42980
rect 18004 42924 18956 42980
rect 19012 42924 19022 42980
rect 30930 42924 30940 42980
rect 30996 42924 35308 42980
rect 35364 42924 35868 42980
rect 35924 42924 35934 42980
rect 37090 42924 37100 42980
rect 37156 42924 37660 42980
rect 37716 42924 40124 42980
rect 40180 42924 40190 42980
rect 44482 42924 44492 42980
rect 44548 42924 45836 42980
rect 45892 42924 45902 42980
rect 3378 42812 3388 42868
rect 3444 42812 3724 42868
rect 3780 42812 3790 42868
rect 23650 42812 23660 42868
rect 23716 42812 29260 42868
rect 29316 42812 30044 42868
rect 30100 42812 30110 42868
rect 33170 42812 33180 42868
rect 33236 42812 33964 42868
rect 34020 42812 34030 42868
rect 38854 42812 38892 42868
rect 38948 42812 38958 42868
rect 41346 42812 41356 42868
rect 41412 42812 42476 42868
rect 42532 42812 42542 42868
rect 43670 42812 43708 42868
rect 43764 42812 43774 42868
rect 44818 42812 44828 42868
rect 44884 42812 45164 42868
rect 45220 42812 45230 42868
rect 8642 42700 8652 42756
rect 8708 42700 9660 42756
rect 9716 42700 9726 42756
rect 13906 42700 13916 42756
rect 13972 42700 14588 42756
rect 14644 42700 15484 42756
rect 15540 42700 15550 42756
rect 20290 42700 20300 42756
rect 20356 42700 21420 42756
rect 21476 42700 21486 42756
rect 26674 42700 26684 42756
rect 26740 42700 27916 42756
rect 27972 42700 27982 42756
rect 29474 42700 29484 42756
rect 29540 42700 31276 42756
rect 31332 42700 31342 42756
rect 32162 42700 32172 42756
rect 32228 42700 34188 42756
rect 34244 42700 34254 42756
rect 3490 42588 3500 42644
rect 3556 42588 4732 42644
rect 4788 42588 5740 42644
rect 5796 42588 5806 42644
rect 6738 42588 6748 42644
rect 6804 42588 10332 42644
rect 10388 42588 10398 42644
rect 12786 42588 12796 42644
rect 12852 42588 14140 42644
rect 14196 42588 14206 42644
rect 25302 42588 25340 42644
rect 25396 42588 25788 42644
rect 25844 42588 25854 42644
rect 26114 42588 26124 42644
rect 26180 42588 26796 42644
rect 26852 42588 26862 42644
rect 34738 42588 34748 42644
rect 34804 42588 37100 42644
rect 37156 42588 37166 42644
rect 40562 42588 40572 42644
rect 40628 42588 48188 42644
rect 48244 42588 48412 42644
rect 48468 42588 48478 42644
rect 1698 42476 1708 42532
rect 1764 42476 2268 42532
rect 2324 42476 3164 42532
rect 3220 42476 6300 42532
rect 6356 42476 6366 42532
rect 7186 42476 7196 42532
rect 7252 42476 7644 42532
rect 7700 42476 7710 42532
rect 12114 42476 12124 42532
rect 12180 42476 13580 42532
rect 13636 42476 13646 42532
rect 16706 42476 16716 42532
rect 16772 42476 16940 42532
rect 16996 42476 17006 42532
rect 17490 42476 17500 42532
rect 17556 42476 19180 42532
rect 19236 42476 21308 42532
rect 21364 42476 21374 42532
rect 21746 42476 21756 42532
rect 21812 42476 22316 42532
rect 22372 42476 25228 42532
rect 25284 42476 25294 42532
rect 29138 42476 29148 42532
rect 29204 42476 29484 42532
rect 29540 42476 30268 42532
rect 30324 42476 30334 42532
rect 39218 42476 39228 42532
rect 39284 42476 40012 42532
rect 40068 42476 43148 42532
rect 43204 42476 43214 42532
rect 44258 42476 44268 42532
rect 44324 42476 46620 42532
rect 46676 42476 46686 42532
rect 2818 42364 2828 42420
rect 2884 42364 6412 42420
rect 6468 42364 9604 42420
rect 33618 42364 33628 42420
rect 33684 42364 43932 42420
rect 43988 42364 43998 42420
rect 9548 42196 9604 42364
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 26226 42252 26236 42308
rect 26292 42252 26684 42308
rect 26740 42252 26750 42308
rect 30034 42252 30044 42308
rect 30100 42252 31836 42308
rect 31892 42252 31902 42308
rect 49200 42196 50000 42224
rect 9538 42140 9548 42196
rect 9604 42140 9614 42196
rect 11666 42140 11676 42196
rect 11732 42140 22876 42196
rect 22932 42140 23324 42196
rect 23380 42140 23390 42196
rect 37202 42140 37212 42196
rect 37268 42140 38948 42196
rect 42130 42140 42140 42196
rect 42196 42140 46956 42196
rect 47012 42140 47022 42196
rect 47180 42140 50000 42196
rect 38892 42084 38948 42140
rect 47180 42084 47236 42140
rect 49200 42112 50000 42140
rect 5730 42028 5740 42084
rect 5796 42028 8764 42084
rect 8820 42028 8830 42084
rect 30706 42028 30716 42084
rect 30772 42028 31500 42084
rect 31556 42028 31566 42084
rect 36418 42028 36428 42084
rect 36484 42028 38332 42084
rect 38388 42028 38668 42084
rect 38724 42028 38734 42084
rect 38882 42028 38892 42084
rect 38948 42028 38958 42084
rect 39778 42028 39788 42084
rect 39844 42028 43484 42084
rect 43540 42028 43550 42084
rect 44930 42028 44940 42084
rect 44996 42028 47236 42084
rect 8530 41916 8540 41972
rect 8596 41916 9660 41972
rect 9716 41916 9726 41972
rect 16818 41916 16828 41972
rect 16884 41916 17500 41972
rect 17556 41916 17566 41972
rect 18386 41916 18396 41972
rect 18452 41916 20524 41972
rect 20580 41916 21420 41972
rect 21476 41916 21486 41972
rect 24658 41916 24668 41972
rect 24724 41916 29260 41972
rect 29316 41916 29326 41972
rect 32498 41916 32508 41972
rect 32564 41916 33628 41972
rect 33684 41916 33694 41972
rect 39890 41916 39900 41972
rect 39956 41916 41132 41972
rect 41188 41916 41198 41972
rect 41458 41916 41468 41972
rect 41524 41916 42588 41972
rect 42644 41916 42654 41972
rect 43362 41916 43372 41972
rect 43428 41916 44828 41972
rect 44884 41916 44894 41972
rect 45490 41916 45500 41972
rect 45556 41916 47516 41972
rect 47572 41916 47582 41972
rect 7298 41804 7308 41860
rect 7364 41804 9436 41860
rect 9492 41804 9502 41860
rect 17378 41804 17388 41860
rect 17444 41804 19068 41860
rect 19124 41804 19404 41860
rect 19460 41804 21532 41860
rect 21588 41804 22204 41860
rect 22260 41804 22270 41860
rect 23202 41804 23212 41860
rect 23268 41804 26908 41860
rect 27906 41804 27916 41860
rect 27972 41804 28812 41860
rect 28868 41804 28878 41860
rect 31154 41804 31164 41860
rect 31220 41804 34412 41860
rect 34468 41804 35532 41860
rect 35588 41804 35598 41860
rect 37202 41804 37212 41860
rect 37268 41804 40460 41860
rect 40516 41804 40526 41860
rect 40898 41804 40908 41860
rect 40964 41804 41804 41860
rect 41860 41804 41870 41860
rect 43698 41804 43708 41860
rect 43764 41804 43820 41860
rect 43876 41804 45276 41860
rect 45332 41804 45342 41860
rect 46274 41804 46284 41860
rect 46340 41804 47964 41860
rect 48020 41804 48030 41860
rect 26852 41748 26908 41804
rect 8082 41692 8092 41748
rect 8148 41692 10108 41748
rect 10164 41692 10174 41748
rect 13458 41692 13468 41748
rect 13524 41692 23772 41748
rect 23828 41692 24332 41748
rect 24388 41692 24398 41748
rect 26852 41692 29036 41748
rect 29092 41692 29932 41748
rect 29988 41692 29998 41748
rect 30594 41692 30604 41748
rect 30660 41692 33068 41748
rect 33124 41692 33134 41748
rect 40338 41692 40348 41748
rect 40404 41692 41692 41748
rect 41748 41692 41758 41748
rect 42802 41692 42812 41748
rect 42868 41692 44044 41748
rect 44100 41692 44268 41748
rect 44324 41692 45052 41748
rect 45108 41692 45118 41748
rect 25554 41580 25564 41636
rect 25620 41580 33404 41636
rect 33460 41580 33740 41636
rect 33796 41580 33806 41636
rect 37426 41580 37436 41636
rect 37492 41580 39452 41636
rect 39508 41580 44940 41636
rect 44996 41580 45006 41636
rect 0 41524 800 41552
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 0 41468 1708 41524
rect 1764 41468 1774 41524
rect 37874 41468 37884 41524
rect 37940 41468 37950 41524
rect 0 41440 800 41468
rect 1362 41356 1372 41412
rect 1428 41356 11564 41412
rect 11620 41356 12460 41412
rect 12516 41356 12526 41412
rect 29250 41356 29260 41412
rect 29316 41356 30156 41412
rect 30212 41356 30222 41412
rect 3826 41244 3836 41300
rect 3892 41244 4620 41300
rect 4676 41244 4686 41300
rect 10658 41244 10668 41300
rect 10724 41244 12012 41300
rect 12068 41244 12684 41300
rect 12740 41244 12750 41300
rect 23986 41244 23996 41300
rect 24052 41244 26908 41300
rect 8306 41132 8316 41188
rect 8372 41132 10220 41188
rect 10276 41132 10286 41188
rect 12338 41132 12348 41188
rect 12404 41132 13468 41188
rect 13524 41132 13534 41188
rect 23874 41020 23884 41076
rect 23940 41020 25844 41076
rect 25788 40964 25844 41020
rect 4722 40908 4732 40964
rect 4788 40908 5852 40964
rect 5908 40908 7084 40964
rect 7140 40908 7150 40964
rect 7746 40908 7756 40964
rect 7812 40908 9772 40964
rect 9828 40908 11676 40964
rect 11732 40908 11742 40964
rect 12226 40908 12236 40964
rect 12292 40908 12302 40964
rect 17490 40908 17500 40964
rect 17556 40908 18396 40964
rect 18452 40908 20524 40964
rect 20580 40908 22316 40964
rect 22372 40908 22382 40964
rect 24098 40908 24108 40964
rect 24164 40908 24892 40964
rect 24948 40908 24958 40964
rect 25778 40908 25788 40964
rect 25844 40908 26124 40964
rect 26180 40908 26190 40964
rect 8306 40796 8316 40852
rect 8372 40796 10668 40852
rect 10724 40796 11564 40852
rect 11620 40796 11630 40852
rect 12236 40740 12292 40908
rect 26852 40852 26908 41244
rect 32386 41132 32396 41188
rect 32452 41132 33068 41188
rect 33124 41132 33134 41188
rect 35186 41132 35196 41188
rect 35252 41132 37436 41188
rect 37492 41132 37502 41188
rect 29138 41020 29148 41076
rect 29204 41020 31948 41076
rect 32004 41020 32014 41076
rect 34290 41020 34300 41076
rect 34356 41020 35980 41076
rect 36036 41020 36046 41076
rect 36418 41020 36428 41076
rect 36484 41020 36876 41076
rect 36932 41020 36942 41076
rect 36306 40908 36316 40964
rect 36372 40908 37548 40964
rect 37604 40908 37614 40964
rect 37884 40852 37940 41468
rect 38658 41356 38668 41412
rect 38724 41356 39116 41412
rect 39172 41356 39182 41412
rect 41804 41244 42924 41300
rect 42980 41244 44492 41300
rect 44548 41244 44558 41300
rect 41804 41188 41860 41244
rect 38882 41132 38892 41188
rect 38948 41132 39004 41188
rect 39060 41132 39070 41188
rect 39666 41132 39676 41188
rect 39732 41132 41804 41188
rect 41860 41132 41870 41188
rect 42466 41132 42476 41188
rect 42532 41132 43820 41188
rect 43876 41132 43886 41188
rect 41234 41020 41244 41076
rect 41300 41020 44940 41076
rect 44996 41020 45006 41076
rect 40002 40908 40012 40964
rect 40068 40908 44156 40964
rect 44212 40908 44604 40964
rect 44660 40908 44670 40964
rect 26852 40796 31948 40852
rect 32004 40796 32014 40852
rect 37884 40796 39228 40852
rect 39284 40796 39294 40852
rect 41122 40796 41132 40852
rect 41188 40796 42588 40852
rect 42644 40796 46284 40852
rect 46340 40796 46350 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 12236 40684 12684 40740
rect 12740 40684 16828 40740
rect 16884 40684 18284 40740
rect 18340 40684 18350 40740
rect 20972 40684 29596 40740
rect 29652 40684 32508 40740
rect 32564 40684 33292 40740
rect 33348 40684 33358 40740
rect 36194 40684 36204 40740
rect 36260 40684 36988 40740
rect 37044 40684 38108 40740
rect 38164 40684 38174 40740
rect 44370 40684 44380 40740
rect 44436 40684 48132 40740
rect 20972 40628 21028 40684
rect 14018 40572 14028 40628
rect 14084 40572 21028 40628
rect 23314 40572 23324 40628
rect 23380 40572 25340 40628
rect 25396 40572 25406 40628
rect 25554 40572 25564 40628
rect 25620 40572 26908 40628
rect 27458 40572 27468 40628
rect 27524 40572 27804 40628
rect 27860 40572 28476 40628
rect 28532 40572 28542 40628
rect 37090 40572 37100 40628
rect 37156 40572 37772 40628
rect 37828 40572 40236 40628
rect 40292 40572 40302 40628
rect 40674 40572 40684 40628
rect 40740 40572 43372 40628
rect 43428 40572 43764 40628
rect 43922 40572 43932 40628
rect 43988 40572 46508 40628
rect 46564 40572 46574 40628
rect 2594 40460 2604 40516
rect 2660 40460 3388 40516
rect 3444 40460 3836 40516
rect 3892 40460 3902 40516
rect 10098 40460 10108 40516
rect 10164 40460 10892 40516
rect 10948 40460 12012 40516
rect 12068 40460 12078 40516
rect 12450 40460 12460 40516
rect 12516 40460 13468 40516
rect 13524 40460 13534 40516
rect 22978 40460 22988 40516
rect 23044 40460 25788 40516
rect 25844 40460 25854 40516
rect 26852 40404 26908 40572
rect 43708 40516 43764 40572
rect 32498 40460 32508 40516
rect 32564 40460 35196 40516
rect 35252 40460 35262 40516
rect 37986 40460 37996 40516
rect 38052 40460 40348 40516
rect 40404 40460 40414 40516
rect 43446 40460 43484 40516
rect 43540 40460 43550 40516
rect 43708 40460 45500 40516
rect 45556 40460 45566 40516
rect 45938 40460 45948 40516
rect 46004 40460 47852 40516
rect 47908 40460 47918 40516
rect 48076 40404 48132 40684
rect 2370 40348 2380 40404
rect 2436 40348 3164 40404
rect 3220 40348 3230 40404
rect 9874 40348 9884 40404
rect 9940 40348 11004 40404
rect 11060 40348 11788 40404
rect 11844 40348 11854 40404
rect 13094 40348 13132 40404
rect 13188 40348 13198 40404
rect 20962 40348 20972 40404
rect 21028 40348 21532 40404
rect 21588 40348 21980 40404
rect 22036 40348 22046 40404
rect 26852 40348 27916 40404
rect 27972 40348 27982 40404
rect 35074 40348 35084 40404
rect 35140 40348 36316 40404
rect 36372 40348 36382 40404
rect 36754 40348 36764 40404
rect 36820 40348 37772 40404
rect 37828 40348 37838 40404
rect 38098 40348 38108 40404
rect 38164 40348 40012 40404
rect 40068 40348 40078 40404
rect 41458 40348 41468 40404
rect 41524 40348 43708 40404
rect 43764 40348 44940 40404
rect 44996 40348 45006 40404
rect 45826 40348 45836 40404
rect 45892 40348 47068 40404
rect 47124 40348 47134 40404
rect 47618 40348 47628 40404
rect 47684 40348 48132 40404
rect 11890 40236 11900 40292
rect 11956 40236 13580 40292
rect 13636 40236 13646 40292
rect 14438 40236 14476 40292
rect 14532 40236 14542 40292
rect 19058 40236 19068 40292
rect 19124 40236 21420 40292
rect 21476 40236 21486 40292
rect 24098 40236 24108 40292
rect 24164 40236 24780 40292
rect 24836 40236 24846 40292
rect 25106 40236 25116 40292
rect 25172 40236 30268 40292
rect 30324 40236 31388 40292
rect 31444 40236 31836 40292
rect 31892 40236 31902 40292
rect 42690 40236 42700 40292
rect 42756 40236 43820 40292
rect 43876 40236 43886 40292
rect 7522 40124 7532 40180
rect 7588 40124 9772 40180
rect 9828 40124 9996 40180
rect 10052 40124 10062 40180
rect 15810 40124 15820 40180
rect 15876 40124 20188 40180
rect 20244 40124 20254 40180
rect 24108 40068 24164 40236
rect 32946 40124 32956 40180
rect 33012 40124 33964 40180
rect 34020 40124 34030 40180
rect 35522 40124 35532 40180
rect 35588 40124 37212 40180
rect 37268 40124 37278 40180
rect 39974 40124 40012 40180
rect 40068 40124 40078 40180
rect 40226 40124 40236 40180
rect 40292 40124 42364 40180
rect 42420 40124 42430 40180
rect 16594 40012 16604 40068
rect 16660 40012 18172 40068
rect 18228 40012 19404 40068
rect 19460 40012 24164 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 30146 39900 30156 39956
rect 30212 39900 33404 39956
rect 33460 39900 33470 39956
rect 37762 39900 37772 39956
rect 37828 39900 38108 39956
rect 38164 39900 41580 39956
rect 41636 39900 42476 39956
rect 42532 39900 42542 39956
rect 20514 39788 20524 39844
rect 20580 39788 21196 39844
rect 21252 39788 22204 39844
rect 22260 39788 23100 39844
rect 23156 39788 23166 39844
rect 28242 39788 28252 39844
rect 28308 39788 29036 39844
rect 29092 39788 29102 39844
rect 36866 39788 36876 39844
rect 36932 39788 37436 39844
rect 37492 39788 38220 39844
rect 38276 39788 38286 39844
rect 9650 39676 9660 39732
rect 9716 39676 10780 39732
rect 10836 39676 10846 39732
rect 17266 39676 17276 39732
rect 17332 39676 19964 39732
rect 20020 39676 20030 39732
rect 22866 39676 22876 39732
rect 22932 39676 26124 39732
rect 26180 39676 26190 39732
rect 27346 39676 27356 39732
rect 27412 39676 29372 39732
rect 29428 39676 32060 39732
rect 32116 39676 33516 39732
rect 33572 39676 35084 39732
rect 35140 39676 35980 39732
rect 36036 39676 36046 39732
rect 13010 39564 13020 39620
rect 13076 39564 13804 39620
rect 13860 39564 13870 39620
rect 20738 39564 20748 39620
rect 20804 39564 22316 39620
rect 22372 39564 22988 39620
rect 23044 39564 23054 39620
rect 30146 39564 30156 39620
rect 30212 39564 31164 39620
rect 31220 39564 31230 39620
rect 31938 39564 31948 39620
rect 32004 39564 34412 39620
rect 34468 39564 35196 39620
rect 35252 39564 35262 39620
rect 8978 39452 8988 39508
rect 9044 39452 9548 39508
rect 9604 39452 9614 39508
rect 10322 39452 10332 39508
rect 10388 39452 11004 39508
rect 11060 39452 11070 39508
rect 15250 39452 15260 39508
rect 15316 39452 22428 39508
rect 22484 39452 22494 39508
rect 22642 39452 22652 39508
rect 22708 39452 24892 39508
rect 24948 39452 24958 39508
rect 26786 39452 26796 39508
rect 26852 39452 28140 39508
rect 28196 39452 28206 39508
rect 29026 39452 29036 39508
rect 29092 39452 32172 39508
rect 32228 39452 33740 39508
rect 33796 39452 33806 39508
rect 42018 39452 42028 39508
rect 42084 39452 42588 39508
rect 42644 39452 42654 39508
rect 44370 39452 44380 39508
rect 44436 39452 44828 39508
rect 44884 39452 44894 39508
rect 1922 39340 1932 39396
rect 1988 39340 3612 39396
rect 3668 39340 5068 39396
rect 5124 39340 5628 39396
rect 5684 39340 8428 39396
rect 8484 39340 9324 39396
rect 9380 39340 9390 39396
rect 9874 39340 9884 39396
rect 9940 39340 11788 39396
rect 11844 39340 11854 39396
rect 15586 39340 15596 39396
rect 15652 39340 17388 39396
rect 17444 39340 17454 39396
rect 19628 39340 28588 39396
rect 28644 39340 29484 39396
rect 29540 39340 29550 39396
rect 34066 39340 34076 39396
rect 34132 39340 37324 39396
rect 37380 39340 37660 39396
rect 37716 39340 37726 39396
rect 10882 39228 10892 39284
rect 10948 39228 14924 39284
rect 14980 39228 14990 39284
rect 19628 39172 19684 39340
rect 42242 39228 42252 39284
rect 42308 39228 44156 39284
rect 44212 39228 45276 39284
rect 45332 39228 45342 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 13906 39116 13916 39172
rect 13972 39116 19684 39172
rect 45042 39116 45052 39172
rect 45108 39116 47404 39172
rect 47460 39116 47470 39172
rect 6962 39004 6972 39060
rect 7028 39004 8092 39060
rect 8148 39004 8540 39060
rect 8596 39004 8606 39060
rect 9202 39004 9212 39060
rect 9268 39004 11116 39060
rect 11172 39004 11182 39060
rect 11554 39004 11564 39060
rect 11620 39004 15932 39060
rect 15988 39004 15998 39060
rect 23202 39004 23212 39060
rect 23268 39004 25004 39060
rect 25060 39004 25070 39060
rect 32274 39004 32284 39060
rect 32340 39004 37884 39060
rect 37940 39004 37950 39060
rect 40002 39004 40012 39060
rect 40068 39004 40348 39060
rect 40404 39004 40414 39060
rect 41010 39004 41020 39060
rect 41076 39004 41468 39060
rect 41524 39004 41534 39060
rect 42018 39004 42028 39060
rect 42084 39004 43260 39060
rect 43316 39004 43326 39060
rect 44034 39004 44044 39060
rect 44100 39004 44828 39060
rect 44884 39004 45388 39060
rect 45444 39004 45454 39060
rect 6850 38892 6860 38948
rect 6916 38892 8316 38948
rect 8372 38892 8652 38948
rect 8708 38892 9660 38948
rect 9716 38892 9726 38948
rect 10966 38892 11004 38948
rect 11060 38892 11070 38948
rect 11218 38892 11228 38948
rect 11284 38892 13580 38948
rect 13636 38892 13646 38948
rect 15026 38892 15036 38948
rect 15092 38892 15260 38948
rect 15316 38892 15326 38948
rect 15474 38892 15484 38948
rect 15540 38892 16380 38948
rect 16436 38892 16446 38948
rect 22418 38892 22428 38948
rect 22484 38892 23660 38948
rect 23716 38892 23726 38948
rect 26852 38892 29148 38948
rect 29204 38892 30044 38948
rect 30100 38892 30110 38948
rect 31266 38892 31276 38948
rect 31332 38892 32508 38948
rect 32564 38892 33404 38948
rect 33460 38892 33470 38948
rect 35634 38892 35644 38948
rect 35700 38892 37212 38948
rect 37268 38892 37278 38948
rect 40786 38892 40796 38948
rect 40852 38892 42476 38948
rect 42532 38892 42542 38948
rect 11228 38836 11284 38892
rect 26852 38836 26908 38892
rect 3154 38780 3164 38836
rect 3220 38780 4172 38836
rect 4228 38780 4508 38836
rect 4564 38780 4844 38836
rect 4900 38780 4910 38836
rect 7522 38780 7532 38836
rect 7588 38780 8204 38836
rect 8260 38780 8270 38836
rect 10098 38780 10108 38836
rect 10164 38780 11284 38836
rect 11442 38780 11452 38836
rect 11508 38780 13020 38836
rect 13076 38780 13086 38836
rect 14018 38780 14028 38836
rect 14084 38780 15204 38836
rect 15148 38724 15204 38780
rect 15372 38780 16044 38836
rect 16100 38780 16110 38836
rect 16930 38780 16940 38836
rect 16996 38780 17724 38836
rect 17780 38780 18844 38836
rect 18900 38780 18910 38836
rect 20066 38780 20076 38836
rect 20132 38780 20748 38836
rect 20804 38780 22204 38836
rect 22260 38780 22876 38836
rect 22932 38780 22942 38836
rect 24658 38780 24668 38836
rect 24724 38780 26908 38836
rect 27794 38780 27804 38836
rect 27860 38780 27870 38836
rect 36876 38780 38780 38836
rect 38836 38780 38846 38836
rect 42578 38780 42588 38836
rect 42644 38780 43260 38836
rect 43316 38780 43326 38836
rect 44818 38780 44828 38836
rect 44884 38780 45500 38836
rect 45556 38780 45566 38836
rect 15372 38724 15428 38780
rect 27804 38724 27860 38780
rect 36876 38724 36932 38780
rect 3378 38668 3388 38724
rect 3444 38668 4396 38724
rect 4452 38668 4956 38724
rect 5012 38668 9548 38724
rect 9604 38668 9614 38724
rect 10546 38668 10556 38724
rect 10612 38668 11564 38724
rect 11620 38668 11630 38724
rect 15148 38668 15428 38724
rect 20402 38668 20412 38724
rect 20468 38668 21420 38724
rect 21476 38668 21486 38724
rect 22306 38668 22316 38724
rect 22372 38668 24108 38724
rect 24164 38668 24174 38724
rect 25228 38668 27860 38724
rect 28354 38668 28364 38724
rect 28420 38668 30324 38724
rect 31826 38668 31836 38724
rect 31892 38668 32732 38724
rect 32788 38668 33180 38724
rect 33236 38668 33246 38724
rect 36866 38668 36876 38724
rect 36932 38668 36942 38724
rect 37202 38668 37212 38724
rect 37268 38668 39004 38724
rect 39060 38668 43036 38724
rect 43092 38668 43102 38724
rect 25228 38612 25284 38668
rect 30268 38612 30324 38668
rect 5170 38556 5180 38612
rect 5236 38556 10780 38612
rect 10836 38556 10846 38612
rect 20290 38556 20300 38612
rect 20356 38556 20972 38612
rect 21028 38556 21038 38612
rect 22978 38556 22988 38612
rect 23044 38556 24668 38612
rect 24724 38556 25228 38612
rect 25284 38556 25294 38612
rect 25442 38556 25452 38612
rect 25508 38556 26012 38612
rect 26068 38556 27132 38612
rect 27188 38556 27198 38612
rect 30268 38556 33852 38612
rect 33908 38556 33918 38612
rect 25228 38500 25284 38556
rect 5842 38444 5852 38500
rect 5908 38444 6636 38500
rect 6692 38444 7644 38500
rect 7700 38444 7710 38500
rect 25228 38444 25676 38500
rect 25732 38444 25742 38500
rect 31938 38444 31948 38500
rect 32004 38444 32396 38500
rect 32452 38444 32462 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 16258 38332 16268 38388
rect 16324 38332 16604 38388
rect 16660 38332 16670 38388
rect 46386 38332 46396 38388
rect 46452 38332 46956 38388
rect 47012 38332 47022 38388
rect 2146 38220 2156 38276
rect 2212 38220 17724 38276
rect 17780 38220 17790 38276
rect 36082 38220 36092 38276
rect 36148 38220 36652 38276
rect 36708 38220 36718 38276
rect 44818 38220 44828 38276
rect 44884 38220 45164 38276
rect 45220 38220 46060 38276
rect 46116 38220 46126 38276
rect 3154 38108 3164 38164
rect 3220 38108 3388 38164
rect 3444 38108 5068 38164
rect 5124 38108 5134 38164
rect 24210 38108 24220 38164
rect 24276 38108 27020 38164
rect 27076 38108 27086 38164
rect 27906 38108 27916 38164
rect 27972 38108 29708 38164
rect 29764 38108 29774 38164
rect 34738 38108 34748 38164
rect 34804 38108 35084 38164
rect 35140 38108 35150 38164
rect 35858 38108 35868 38164
rect 35924 38108 37548 38164
rect 37604 38108 37614 38164
rect 43474 38108 43484 38164
rect 43540 38108 43708 38164
rect 43764 38108 44044 38164
rect 44100 38108 44110 38164
rect 45042 38108 45052 38164
rect 45108 38108 47404 38164
rect 47460 38108 47470 38164
rect 7074 37996 7084 38052
rect 7140 37996 7980 38052
rect 8036 37996 8046 38052
rect 12898 37996 12908 38052
rect 12964 37996 13580 38052
rect 13636 37996 13646 38052
rect 14578 37996 14588 38052
rect 14644 37996 15372 38052
rect 15428 37996 15438 38052
rect 23538 37996 23548 38052
rect 23604 37996 24332 38052
rect 24388 37996 24398 38052
rect 30818 37996 30828 38052
rect 30884 37996 32284 38052
rect 32340 37996 32350 38052
rect 34178 37996 34188 38052
rect 34244 37996 47628 38052
rect 47684 37996 47694 38052
rect 10434 37884 10444 37940
rect 10500 37884 15596 37940
rect 15652 37884 15662 37940
rect 18162 37884 18172 37940
rect 18228 37884 21532 37940
rect 21588 37884 21598 37940
rect 26338 37884 26348 37940
rect 26404 37884 27580 37940
rect 27636 37884 27646 37940
rect 32722 37884 32732 37940
rect 32788 37884 34412 37940
rect 34468 37884 34478 37940
rect 34850 37884 34860 37940
rect 34916 37884 36092 37940
rect 36148 37884 37772 37940
rect 37828 37884 37838 37940
rect 40786 37884 40796 37940
rect 40852 37884 41916 37940
rect 41972 37884 41982 37940
rect 45126 37884 45164 37940
rect 45220 37884 45230 37940
rect 46834 37884 46844 37940
rect 46900 37884 48076 37940
rect 48132 37884 48142 37940
rect 12124 37828 12180 37884
rect 4722 37772 4732 37828
rect 4788 37772 5292 37828
rect 5348 37772 5358 37828
rect 5506 37772 5516 37828
rect 5572 37772 5610 37828
rect 8754 37772 8764 37828
rect 8820 37772 9324 37828
rect 9380 37772 9390 37828
rect 9538 37772 9548 37828
rect 9604 37772 11004 37828
rect 11060 37772 11070 37828
rect 11554 37772 11564 37828
rect 11620 37772 11630 37828
rect 12114 37772 12124 37828
rect 12180 37772 12190 37828
rect 15698 37772 15708 37828
rect 15764 37772 20748 37828
rect 20804 37772 20814 37828
rect 22642 37772 22652 37828
rect 22708 37772 23884 37828
rect 23940 37772 23950 37828
rect 29586 37772 29596 37828
rect 29652 37772 30828 37828
rect 30884 37772 30894 37828
rect 35298 37772 35308 37828
rect 35364 37772 36204 37828
rect 36260 37772 36270 37828
rect 38210 37772 38220 37828
rect 38276 37772 39116 37828
rect 39172 37772 39182 37828
rect 39890 37772 39900 37828
rect 39956 37772 41132 37828
rect 41188 37772 41198 37828
rect 41794 37772 41804 37828
rect 41860 37772 43148 37828
rect 43204 37772 43214 37828
rect 43586 37772 43596 37828
rect 43652 37772 46732 37828
rect 46788 37772 46798 37828
rect 11564 37716 11620 37772
rect 11564 37660 17948 37716
rect 18004 37660 18396 37716
rect 18452 37660 18462 37716
rect 28466 37660 28476 37716
rect 28532 37660 29260 37716
rect 29316 37660 30268 37716
rect 30324 37660 31388 37716
rect 31444 37660 31454 37716
rect 48066 37660 48076 37716
rect 48132 37660 48142 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 9090 37548 9100 37604
rect 9156 37548 9660 37604
rect 9716 37548 12908 37604
rect 12964 37548 12974 37604
rect 23762 37548 23772 37604
rect 23828 37548 29484 37604
rect 29540 37548 30044 37604
rect 30100 37548 31500 37604
rect 31556 37548 31566 37604
rect 37538 37548 37548 37604
rect 37604 37548 38668 37604
rect 38612 37492 38668 37548
rect 48076 37492 48132 37660
rect 1474 37436 1484 37492
rect 1540 37436 3388 37492
rect 3490 37436 3500 37492
rect 3556 37436 4732 37492
rect 4788 37436 4798 37492
rect 5170 37436 5180 37492
rect 5236 37436 7644 37492
rect 7700 37436 7710 37492
rect 9762 37436 9772 37492
rect 9828 37436 10220 37492
rect 10276 37436 10286 37492
rect 13020 37436 18900 37492
rect 31042 37436 31052 37492
rect 31108 37436 33740 37492
rect 33796 37436 33806 37492
rect 35970 37436 35980 37492
rect 36036 37436 37436 37492
rect 37492 37436 38220 37492
rect 38276 37436 38286 37492
rect 38612 37436 41188 37492
rect 44454 37436 44492 37492
rect 44548 37436 44558 37492
rect 47730 37436 47740 37492
rect 47796 37436 48132 37492
rect 3332 37380 3388 37436
rect 13020 37380 13076 37436
rect 3332 37324 8428 37380
rect 8484 37324 8988 37380
rect 9044 37324 9054 37380
rect 10658 37324 10668 37380
rect 10724 37324 11900 37380
rect 11956 37324 11966 37380
rect 13010 37324 13020 37380
rect 13076 37324 13086 37380
rect 4274 37212 4284 37268
rect 4340 37212 5516 37268
rect 5572 37212 5582 37268
rect 5842 37212 5852 37268
rect 5908 37212 6860 37268
rect 6916 37212 6926 37268
rect 10434 37212 10444 37268
rect 10500 37212 11340 37268
rect 11396 37212 11406 37268
rect 12114 37212 12124 37268
rect 12180 37212 12460 37268
rect 12516 37212 12526 37268
rect 14130 37212 14140 37268
rect 14196 37212 17500 37268
rect 17556 37212 17566 37268
rect 18844 37156 18900 37436
rect 41132 37380 41188 37436
rect 28242 37324 28252 37380
rect 28308 37324 29260 37380
rect 29316 37324 29326 37380
rect 34290 37324 34300 37380
rect 34356 37324 35196 37380
rect 35252 37324 35262 37380
rect 36978 37324 36988 37380
rect 37044 37324 38780 37380
rect 38836 37324 39116 37380
rect 39172 37324 39182 37380
rect 41122 37324 41132 37380
rect 41188 37324 41198 37380
rect 49200 37268 50000 37296
rect 26086 37212 26124 37268
rect 26180 37212 26190 37268
rect 30034 37212 30044 37268
rect 30100 37212 31948 37268
rect 32004 37212 32508 37268
rect 32564 37212 33516 37268
rect 33572 37212 33582 37268
rect 36194 37212 36204 37268
rect 36260 37212 37212 37268
rect 37268 37212 37278 37268
rect 43250 37212 43260 37268
rect 43316 37212 48300 37268
rect 48356 37212 50000 37268
rect 49200 37184 50000 37212
rect 2482 37100 2492 37156
rect 2548 37100 5964 37156
rect 6020 37100 6030 37156
rect 15036 37100 16268 37156
rect 16324 37100 16334 37156
rect 18806 37100 18844 37156
rect 18900 37100 18910 37156
rect 40338 37100 40348 37156
rect 40404 37100 41916 37156
rect 41972 37100 41982 37156
rect 42690 37100 42700 37156
rect 42756 37100 43932 37156
rect 43988 37100 43998 37156
rect 44930 37100 44940 37156
rect 44996 37100 45724 37156
rect 45780 37100 45790 37156
rect 15036 37044 15092 37100
rect 2146 36988 2156 37044
rect 2212 36988 5124 37044
rect 5282 36988 5292 37044
rect 5348 36988 6188 37044
rect 6244 36988 10444 37044
rect 10500 36988 10510 37044
rect 15026 36988 15036 37044
rect 15092 36988 15102 37044
rect 16370 36988 16380 37044
rect 16436 36988 17500 37044
rect 17556 36988 17566 37044
rect 18386 36988 18396 37044
rect 18452 36988 18732 37044
rect 18788 36988 18798 37044
rect 19842 36988 19852 37044
rect 19908 36988 20748 37044
rect 20804 36988 20814 37044
rect 43474 36988 43484 37044
rect 43540 36988 45220 37044
rect 45378 36988 45388 37044
rect 45444 36988 47740 37044
rect 47796 36988 47806 37044
rect 5068 36932 5124 36988
rect 45164 36932 45220 36988
rect 5068 36876 5180 36932
rect 5236 36876 5404 36932
rect 5460 36876 5470 36932
rect 25218 36876 25228 36932
rect 25284 36876 26348 36932
rect 26404 36876 26414 36932
rect 43138 36876 43148 36932
rect 43204 36876 44492 36932
rect 44548 36876 44558 36932
rect 45164 36876 47404 36932
rect 47460 36876 47470 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 5282 36764 5292 36820
rect 5348 36764 5516 36820
rect 5572 36764 5582 36820
rect 8530 36764 8540 36820
rect 8596 36764 8876 36820
rect 8932 36764 8942 36820
rect 10322 36764 10332 36820
rect 10388 36764 13132 36820
rect 13188 36764 13198 36820
rect 19058 36764 19068 36820
rect 19124 36764 20188 36820
rect 20244 36764 20254 36820
rect 35634 36764 35644 36820
rect 35700 36764 36316 36820
rect 36372 36764 36382 36820
rect 14354 36652 14364 36708
rect 14420 36652 14700 36708
rect 14756 36652 14766 36708
rect 19394 36652 19404 36708
rect 19460 36652 21308 36708
rect 21364 36652 21374 36708
rect 21746 36652 21756 36708
rect 21812 36652 22764 36708
rect 22820 36652 22830 36708
rect 25890 36652 25900 36708
rect 25956 36652 26796 36708
rect 26852 36652 27580 36708
rect 27636 36652 27646 36708
rect 37090 36652 37100 36708
rect 37156 36652 37996 36708
rect 38052 36652 39732 36708
rect 19170 36540 19180 36596
rect 19236 36540 20412 36596
rect 20468 36540 20478 36596
rect 23762 36540 23772 36596
rect 23828 36540 28924 36596
rect 28980 36540 28990 36596
rect 39676 36484 39732 36652
rect 3938 36428 3948 36484
rect 4004 36428 4396 36484
rect 4452 36428 5068 36484
rect 5124 36428 5134 36484
rect 6178 36428 6188 36484
rect 6244 36428 7196 36484
rect 7252 36428 8204 36484
rect 8260 36428 8270 36484
rect 8754 36428 8764 36484
rect 8820 36428 9212 36484
rect 9268 36428 9278 36484
rect 12002 36428 12012 36484
rect 12068 36428 12460 36484
rect 12516 36428 12526 36484
rect 14802 36428 14812 36484
rect 14868 36428 15036 36484
rect 15092 36428 15102 36484
rect 18834 36428 18844 36484
rect 18900 36428 19964 36484
rect 20020 36428 20030 36484
rect 20738 36428 20748 36484
rect 20804 36428 21532 36484
rect 21588 36428 21598 36484
rect 22754 36428 22764 36484
rect 22820 36428 23996 36484
rect 24052 36428 24062 36484
rect 26562 36428 26572 36484
rect 26628 36428 27356 36484
rect 27412 36428 27422 36484
rect 32946 36428 32956 36484
rect 33012 36428 33628 36484
rect 33684 36428 33694 36484
rect 34738 36428 34748 36484
rect 34804 36428 39340 36484
rect 39396 36428 39406 36484
rect 39666 36428 39676 36484
rect 39732 36428 39742 36484
rect 42130 36428 42140 36484
rect 42196 36428 43148 36484
rect 43204 36428 43214 36484
rect 4834 36316 4844 36372
rect 4900 36316 5852 36372
rect 5908 36316 6636 36372
rect 6692 36316 7420 36372
rect 7476 36316 7486 36372
rect 19618 36316 19628 36372
rect 19684 36316 19740 36372
rect 19796 36316 19806 36372
rect 27010 36316 27020 36372
rect 27076 36316 29148 36372
rect 29204 36316 29214 36372
rect 31042 36316 31052 36372
rect 31108 36316 32396 36372
rect 32452 36316 33180 36372
rect 33236 36316 33246 36372
rect 35074 36316 35084 36372
rect 35140 36316 35756 36372
rect 35812 36316 36988 36372
rect 37044 36316 37054 36372
rect 37874 36316 37884 36372
rect 37940 36316 38556 36372
rect 38612 36316 38622 36372
rect 39218 36316 39228 36372
rect 39284 36316 42364 36372
rect 42420 36316 42430 36372
rect 43810 36316 43820 36372
rect 43876 36316 44604 36372
rect 44660 36316 44670 36372
rect 2482 36204 2492 36260
rect 2548 36204 6412 36260
rect 6468 36204 6478 36260
rect 7494 36204 7532 36260
rect 7588 36204 7598 36260
rect 8194 36204 8204 36260
rect 8260 36204 8652 36260
rect 8708 36204 8718 36260
rect 18162 36204 18172 36260
rect 18228 36204 19068 36260
rect 19124 36204 19134 36260
rect 19506 36204 19516 36260
rect 19572 36204 19852 36260
rect 19908 36204 19918 36260
rect 20178 36204 20188 36260
rect 20244 36204 20636 36260
rect 20692 36204 22204 36260
rect 22260 36204 22652 36260
rect 22708 36204 22718 36260
rect 26786 36204 26796 36260
rect 26852 36204 28588 36260
rect 28644 36204 40348 36260
rect 40404 36204 40414 36260
rect 41458 36204 41468 36260
rect 41524 36204 42476 36260
rect 42532 36204 45164 36260
rect 45220 36204 45948 36260
rect 46004 36204 46014 36260
rect 5058 36092 5068 36148
rect 5124 36092 8092 36148
rect 8148 36092 8158 36148
rect 13234 36092 13244 36148
rect 13300 36092 15148 36148
rect 15204 36092 15484 36148
rect 15540 36092 15550 36148
rect 35970 36092 35980 36148
rect 36036 36092 36540 36148
rect 36596 36092 39564 36148
rect 39620 36092 39630 36148
rect 41122 36092 41132 36148
rect 41188 36092 42140 36148
rect 42196 36092 42206 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 41132 36036 41188 36092
rect 14438 35980 14476 36036
rect 14532 35980 14542 36036
rect 19590 35980 19628 36036
rect 19684 35980 19694 36036
rect 22204 35980 23100 36036
rect 23156 35980 23166 36036
rect 33954 35980 33964 36036
rect 34020 35980 41188 36036
rect 41346 35980 41356 36036
rect 41412 35980 41422 36036
rect 42466 35980 42476 36036
rect 42532 35980 43036 36036
rect 43092 35980 43820 36036
rect 43876 35980 44268 36036
rect 44324 35980 45500 36036
rect 45556 35980 45566 36036
rect 22204 35924 22260 35980
rect 41356 35924 41412 35980
rect 6514 35868 6524 35924
rect 6580 35868 7644 35924
rect 7700 35868 7710 35924
rect 9762 35868 9772 35924
rect 9828 35868 10668 35924
rect 10724 35868 10892 35924
rect 10948 35868 10958 35924
rect 12674 35868 12684 35924
rect 12740 35868 13132 35924
rect 13188 35868 13198 35924
rect 13682 35868 13692 35924
rect 13748 35868 22260 35924
rect 22418 35868 22428 35924
rect 22484 35868 23660 35924
rect 23716 35868 25900 35924
rect 25956 35868 26460 35924
rect 26516 35868 26526 35924
rect 30034 35868 30044 35924
rect 30100 35868 32172 35924
rect 32228 35868 32238 35924
rect 33506 35868 33516 35924
rect 33572 35868 35644 35924
rect 35700 35868 35710 35924
rect 39330 35868 39340 35924
rect 39396 35868 41412 35924
rect 42802 35868 42812 35924
rect 42868 35868 43596 35924
rect 43652 35868 46396 35924
rect 46452 35868 46462 35924
rect 42812 35812 42868 35868
rect 6290 35756 6300 35812
rect 6356 35756 7084 35812
rect 7140 35756 7150 35812
rect 9986 35756 9996 35812
rect 10052 35756 14028 35812
rect 14084 35756 14094 35812
rect 23202 35756 23212 35812
rect 23268 35756 25340 35812
rect 25396 35756 25406 35812
rect 27682 35756 27692 35812
rect 27748 35756 29260 35812
rect 29316 35756 29326 35812
rect 32274 35756 32284 35812
rect 32340 35756 34188 35812
rect 34244 35756 34254 35812
rect 38546 35756 38556 35812
rect 38612 35756 38892 35812
rect 38948 35756 40124 35812
rect 40180 35756 42868 35812
rect 11890 35644 11900 35700
rect 11956 35644 12572 35700
rect 12628 35644 14252 35700
rect 14308 35644 14318 35700
rect 17378 35644 17388 35700
rect 17444 35644 18284 35700
rect 18340 35644 18956 35700
rect 19012 35644 19022 35700
rect 20290 35644 20300 35700
rect 20356 35644 21084 35700
rect 21140 35644 21150 35700
rect 23202 35644 23212 35700
rect 23268 35644 23996 35700
rect 24052 35644 25004 35700
rect 25060 35644 25070 35700
rect 26852 35644 28588 35700
rect 28644 35644 28654 35700
rect 29138 35644 29148 35700
rect 29204 35644 29372 35700
rect 29428 35644 30492 35700
rect 30548 35644 30558 35700
rect 30930 35644 30940 35700
rect 30996 35644 31948 35700
rect 32004 35644 32014 35700
rect 41682 35644 41692 35700
rect 41748 35644 42924 35700
rect 42980 35644 43596 35700
rect 43652 35644 43662 35700
rect 11778 35532 11788 35588
rect 11844 35532 13468 35588
rect 13524 35532 14364 35588
rect 14420 35532 14430 35588
rect 19170 35532 19180 35588
rect 19236 35532 20636 35588
rect 20692 35532 20702 35588
rect 26786 35532 26796 35588
rect 26852 35532 26908 35644
rect 29148 35588 29204 35644
rect 27458 35532 27468 35588
rect 27524 35532 29204 35588
rect 31602 35532 31612 35588
rect 31668 35532 36316 35588
rect 36372 35532 36382 35588
rect 41206 35532 41244 35588
rect 41300 35532 41310 35588
rect 44034 35532 44044 35588
rect 44100 35532 44492 35588
rect 44548 35532 48188 35588
rect 48244 35532 48254 35588
rect 8502 35420 8540 35476
rect 8596 35420 8606 35476
rect 12786 35420 12796 35476
rect 12852 35420 14028 35476
rect 14084 35420 14094 35476
rect 16678 35420 16716 35476
rect 16772 35420 16782 35476
rect 5730 35308 5740 35364
rect 5796 35308 6524 35364
rect 6580 35308 6590 35364
rect 6748 35308 10444 35364
rect 10500 35308 10510 35364
rect 13570 35308 13580 35364
rect 13636 35308 15036 35364
rect 15092 35308 16156 35364
rect 16212 35308 16222 35364
rect 37426 35308 37436 35364
rect 37492 35308 38780 35364
rect 38836 35308 38846 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 6748 35252 6804 35308
rect 34066 35252 34076 35308
rect 34132 35252 34142 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 4844 35196 6804 35252
rect 13794 35196 13804 35252
rect 13860 35196 13870 35252
rect 14354 35196 14364 35252
rect 14420 35196 16604 35252
rect 16660 35196 16670 35252
rect 4844 35140 4900 35196
rect 2258 35084 2268 35140
rect 2324 35084 2716 35140
rect 2772 35084 3724 35140
rect 3780 35084 4900 35140
rect 10994 35084 11004 35140
rect 11060 35084 11900 35140
rect 11956 35084 13244 35140
rect 13300 35084 13310 35140
rect 13804 35028 13860 35196
rect 34076 35140 34132 35252
rect 40338 35196 40348 35252
rect 40404 35196 45388 35252
rect 45444 35196 45454 35252
rect 14130 35084 14140 35140
rect 14196 35084 14812 35140
rect 14868 35084 16268 35140
rect 16324 35084 16334 35140
rect 19478 35084 19516 35140
rect 19572 35084 19582 35140
rect 22316 35084 24668 35140
rect 24724 35084 24734 35140
rect 34076 35084 34636 35140
rect 34692 35084 34702 35140
rect 35298 35084 35308 35140
rect 35364 35084 35644 35140
rect 35700 35084 35710 35140
rect 22316 35028 22372 35084
rect 9874 34972 9884 35028
rect 9940 34972 11116 35028
rect 11172 34972 11182 35028
rect 13804 34972 15372 35028
rect 15428 34972 15438 35028
rect 16380 34972 22316 35028
rect 22372 34972 22382 35028
rect 24322 34972 24332 35028
rect 24388 34972 27244 35028
rect 27300 34972 27310 35028
rect 30146 34972 30156 35028
rect 30212 34972 31276 35028
rect 31332 34972 32732 35028
rect 32788 34972 33292 35028
rect 33348 34972 33358 35028
rect 33842 34972 33852 35028
rect 33908 34972 34188 35028
rect 34244 34972 34254 35028
rect 34962 34972 34972 35028
rect 35028 34972 35980 35028
rect 36036 34972 36046 35028
rect 47170 34972 47180 35028
rect 47236 34972 48188 35028
rect 48244 34972 48254 35028
rect 16380 34916 16436 34972
rect 5170 34860 5180 34916
rect 5236 34860 5628 34916
rect 5684 34860 7196 34916
rect 7252 34860 9996 34916
rect 10052 34860 10062 34916
rect 12562 34860 12572 34916
rect 12628 34860 13916 34916
rect 13972 34860 14700 34916
rect 14756 34860 14766 34916
rect 15092 34860 16436 34916
rect 16594 34860 16604 34916
rect 16660 34860 17276 34916
rect 17332 34860 17342 34916
rect 19618 34860 19628 34916
rect 19684 34860 20076 34916
rect 20132 34860 20142 34916
rect 21410 34860 21420 34916
rect 21476 34860 21980 34916
rect 22036 34860 22046 34916
rect 24098 34860 24108 34916
rect 24164 34860 27580 34916
rect 27636 34860 27646 34916
rect 31378 34860 31388 34916
rect 31444 34860 31948 34916
rect 32004 34860 34300 34916
rect 34356 34860 34366 34916
rect 35186 34860 35196 34916
rect 35252 34860 36204 34916
rect 36260 34860 36270 34916
rect 41906 34860 41916 34916
rect 41972 34860 42924 34916
rect 42980 34860 42990 34916
rect 1810 34748 1820 34804
rect 1876 34748 3052 34804
rect 3108 34748 4172 34804
rect 4228 34748 4238 34804
rect 8194 34748 8204 34804
rect 8260 34748 9772 34804
rect 9828 34748 9838 34804
rect 10322 34748 10332 34804
rect 10388 34748 12012 34804
rect 12068 34748 13804 34804
rect 13860 34748 13870 34804
rect 15092 34692 15148 34860
rect 18498 34748 18508 34804
rect 18564 34748 19964 34804
rect 20020 34748 20030 34804
rect 20178 34748 20188 34804
rect 20244 34748 22204 34804
rect 22260 34748 23548 34804
rect 23604 34748 25116 34804
rect 25172 34748 25182 34804
rect 27346 34748 27356 34804
rect 27412 34748 30940 34804
rect 30996 34748 31276 34804
rect 31332 34748 31724 34804
rect 31780 34748 31790 34804
rect 32386 34748 32396 34804
rect 32452 34748 33404 34804
rect 33460 34748 36428 34804
rect 36484 34748 36494 34804
rect 44258 34748 44268 34804
rect 44324 34748 45724 34804
rect 45780 34748 45790 34804
rect 1698 34636 1708 34692
rect 1764 34636 3388 34692
rect 3444 34636 4620 34692
rect 4676 34636 4686 34692
rect 5142 34636 5180 34692
rect 5236 34636 5246 34692
rect 9090 34636 9100 34692
rect 9156 34636 11116 34692
rect 11172 34636 11182 34692
rect 11666 34636 11676 34692
rect 11732 34636 13132 34692
rect 13188 34636 15148 34692
rect 19628 34636 19852 34692
rect 19908 34636 19918 34692
rect 20626 34636 20636 34692
rect 20692 34636 23100 34692
rect 23156 34636 23166 34692
rect 32834 34636 32844 34692
rect 32900 34636 33516 34692
rect 33572 34636 33582 34692
rect 35242 34636 35252 34692
rect 35308 34636 35644 34692
rect 35700 34636 35710 34692
rect 36306 34636 36316 34692
rect 36372 34636 37212 34692
rect 37268 34636 37278 34692
rect 42578 34636 42588 34692
rect 42644 34636 44380 34692
rect 44436 34636 44446 34692
rect 44930 34636 44940 34692
rect 44996 34636 45276 34692
rect 45332 34636 47852 34692
rect 47908 34636 47918 34692
rect 7410 34524 7420 34580
rect 7476 34524 8540 34580
rect 8596 34524 9436 34580
rect 9492 34524 9502 34580
rect 15250 34524 15260 34580
rect 15316 34524 17612 34580
rect 17668 34524 17678 34580
rect 1922 34412 1932 34468
rect 1988 34412 1998 34468
rect 6038 34412 6076 34468
rect 6132 34412 6142 34468
rect 15026 34412 15036 34468
rect 15092 34412 16044 34468
rect 16100 34412 16110 34468
rect 1932 34020 1988 34412
rect 19628 34356 19684 34636
rect 23846 34524 23884 34580
rect 23940 34524 23950 34580
rect 35410 34524 35420 34580
rect 35476 34524 35868 34580
rect 35924 34524 35934 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 23958 34412 23996 34468
rect 24052 34412 24062 34468
rect 29138 34412 29148 34468
rect 29204 34412 29214 34468
rect 12338 34300 12348 34356
rect 12404 34300 14364 34356
rect 14420 34300 14430 34356
rect 19170 34300 19180 34356
rect 19236 34300 24108 34356
rect 24164 34300 24174 34356
rect 2818 34188 2828 34244
rect 2884 34188 5068 34244
rect 5124 34188 5134 34244
rect 11666 34188 11676 34244
rect 11732 34188 15148 34244
rect 15204 34188 15820 34244
rect 15876 34188 15886 34244
rect 17714 34188 17724 34244
rect 17780 34188 22652 34244
rect 22708 34188 22718 34244
rect 23650 34188 23660 34244
rect 23716 34188 24332 34244
rect 24388 34188 24398 34244
rect 29148 34132 29204 34412
rect 29558 34300 29596 34356
rect 29652 34300 29662 34356
rect 4834 34076 4844 34132
rect 4900 34076 5628 34132
rect 5684 34076 7084 34132
rect 7140 34076 7150 34132
rect 8082 34076 8092 34132
rect 8148 34076 10332 34132
rect 10388 34076 10398 34132
rect 14354 34076 14364 34132
rect 14420 34076 16044 34132
rect 16100 34076 17836 34132
rect 17892 34076 17902 34132
rect 18050 34076 18060 34132
rect 18116 34076 18284 34132
rect 18340 34076 18508 34132
rect 18564 34076 18574 34132
rect 18722 34076 18732 34132
rect 18788 34076 18826 34132
rect 19506 34076 19516 34132
rect 19572 34076 19740 34132
rect 19796 34076 19806 34132
rect 23314 34076 23324 34132
rect 23380 34076 24556 34132
rect 24612 34076 24622 34132
rect 25330 34076 25340 34132
rect 25396 34076 29708 34132
rect 29764 34076 29774 34132
rect 38994 34076 39004 34132
rect 39060 34076 39676 34132
rect 39732 34076 41468 34132
rect 41524 34076 41534 34132
rect 24556 34020 24612 34076
rect 1922 33964 1932 34020
rect 1988 33964 1998 34020
rect 7746 33964 7756 34020
rect 7812 33964 9772 34020
rect 9828 33964 9838 34020
rect 10098 33964 10108 34020
rect 10164 33964 11004 34020
rect 11060 33964 11070 34020
rect 24556 33964 26572 34020
rect 26628 33964 26638 34020
rect 6066 33852 6076 33908
rect 6132 33852 6636 33908
rect 6692 33852 8316 33908
rect 8372 33852 13580 33908
rect 13636 33852 13646 33908
rect 14018 33852 14028 33908
rect 14084 33852 16268 33908
rect 16324 33852 16334 33908
rect 19170 33852 19180 33908
rect 19236 33852 20188 33908
rect 20244 33852 20254 33908
rect 33506 33852 33516 33908
rect 33572 33852 39116 33908
rect 39172 33852 39182 33908
rect 10322 33740 10332 33796
rect 10388 33740 10892 33796
rect 10948 33740 10958 33796
rect 21970 33740 21980 33796
rect 22036 33740 23884 33796
rect 23940 33740 23950 33796
rect 38770 33740 38780 33796
rect 38836 33740 41692 33796
rect 41748 33740 41758 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 2370 33628 2380 33684
rect 2436 33628 4228 33684
rect 5618 33628 5628 33684
rect 5684 33628 12236 33684
rect 12292 33628 14252 33684
rect 14308 33628 15036 33684
rect 15092 33628 15102 33684
rect 21522 33628 21532 33684
rect 21588 33628 23436 33684
rect 23492 33628 23502 33684
rect 24658 33628 24668 33684
rect 24724 33628 25284 33684
rect 26226 33628 26236 33684
rect 26292 33628 30212 33684
rect 40114 33628 40124 33684
rect 40180 33628 40908 33684
rect 40964 33628 40974 33684
rect 2930 33516 2940 33572
rect 2996 33516 3276 33572
rect 3332 33516 3342 33572
rect 4172 33236 4228 33628
rect 25228 33572 25284 33628
rect 30156 33572 30212 33628
rect 5618 33516 5628 33572
rect 5684 33516 6412 33572
rect 6468 33516 6478 33572
rect 8866 33516 8876 33572
rect 8932 33516 14028 33572
rect 14084 33516 14094 33572
rect 15092 33516 20748 33572
rect 20804 33516 20814 33572
rect 25228 33516 27468 33572
rect 27524 33516 27534 33572
rect 30156 33516 32508 33572
rect 32564 33516 32574 33572
rect 37986 33516 37996 33572
rect 38052 33516 39396 33572
rect 15092 33460 15148 33516
rect 7970 33404 7980 33460
rect 8036 33404 9996 33460
rect 10052 33404 10062 33460
rect 13570 33404 13580 33460
rect 13636 33404 15148 33460
rect 20514 33404 20524 33460
rect 20580 33404 22876 33460
rect 22932 33404 23436 33460
rect 23492 33404 23502 33460
rect 35252 33404 35420 33460
rect 35476 33404 35486 33460
rect 35858 33404 35868 33460
rect 35924 33404 37324 33460
rect 37380 33404 37390 33460
rect 35252 33348 35308 33404
rect 39340 33348 39396 33516
rect 41346 33404 41356 33460
rect 41412 33404 42252 33460
rect 42308 33404 42318 33460
rect 8978 33292 8988 33348
rect 9044 33292 10556 33348
rect 10612 33292 11676 33348
rect 11732 33292 11742 33348
rect 12002 33292 12012 33348
rect 12068 33292 17164 33348
rect 17220 33292 18172 33348
rect 18228 33292 18238 33348
rect 19058 33292 19068 33348
rect 19124 33292 20300 33348
rect 20356 33292 20366 33348
rect 32050 33292 32060 33348
rect 32116 33292 35308 33348
rect 36418 33292 36428 33348
rect 36484 33292 38668 33348
rect 38724 33292 38734 33348
rect 39330 33292 39340 33348
rect 39396 33292 39406 33348
rect 46722 33292 46732 33348
rect 46788 33292 47852 33348
rect 47908 33292 47918 33348
rect 1670 33180 1708 33236
rect 1764 33180 1774 33236
rect 4162 33180 4172 33236
rect 4228 33180 7420 33236
rect 7476 33180 7532 33236
rect 7588 33180 13580 33236
rect 13636 33180 13646 33236
rect 14886 33180 14924 33236
rect 14980 33180 14990 33236
rect 24434 33180 24444 33236
rect 24500 33180 25452 33236
rect 25508 33180 25518 33236
rect 31490 33180 31500 33236
rect 31556 33180 35756 33236
rect 35812 33180 35822 33236
rect 36082 33180 36092 33236
rect 36148 33180 36988 33236
rect 37044 33180 37054 33236
rect 43698 33180 43708 33236
rect 43764 33180 44828 33236
rect 44884 33180 44894 33236
rect 46162 33180 46172 33236
rect 46228 33180 47516 33236
rect 47572 33180 47582 33236
rect 35756 33124 35812 33180
rect 2006 33068 2044 33124
rect 2100 33068 2110 33124
rect 8754 33068 8764 33124
rect 8820 33068 11452 33124
rect 11508 33068 11518 33124
rect 13654 33068 13692 33124
rect 13748 33068 13758 33124
rect 20374 33068 20412 33124
rect 20468 33068 20478 33124
rect 26338 33068 26348 33124
rect 26404 33068 29260 33124
rect 29316 33068 29326 33124
rect 35756 33068 37212 33124
rect 37268 33068 37278 33124
rect 37426 33068 37436 33124
rect 37492 33068 38108 33124
rect 38164 33068 38174 33124
rect 43810 33068 43820 33124
rect 43876 33068 44380 33124
rect 44436 33068 44446 33124
rect 46610 33068 46620 33124
rect 46676 33068 47180 33124
rect 47236 33068 47246 33124
rect 2230 32956 2268 33012
rect 2324 32956 2334 33012
rect 3826 32956 3836 33012
rect 3892 32956 4172 33012
rect 4228 32956 4238 33012
rect 25442 32956 25452 33012
rect 25508 32956 26012 33012
rect 26068 32956 26078 33012
rect 33842 32956 33852 33012
rect 33908 32956 41916 33012
rect 41972 32956 43036 33012
rect 43092 32956 43372 33012
rect 43428 32956 43438 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 3154 32844 3164 32900
rect 3220 32844 5628 32900
rect 5684 32844 5694 32900
rect 14018 32844 14028 32900
rect 14084 32844 15932 32900
rect 15988 32844 15998 32900
rect 16482 32844 16492 32900
rect 16548 32844 16716 32900
rect 16772 32844 16782 32900
rect 20514 32844 20524 32900
rect 20580 32844 23436 32900
rect 23492 32844 24444 32900
rect 24500 32844 24510 32900
rect 38322 32844 38332 32900
rect 38388 32844 41580 32900
rect 41636 32844 41646 32900
rect 4918 32732 4956 32788
rect 5012 32732 5022 32788
rect 11218 32732 11228 32788
rect 11284 32732 11900 32788
rect 11956 32732 11966 32788
rect 15362 32732 15372 32788
rect 15428 32732 16156 32788
rect 16212 32732 16222 32788
rect 23426 32732 23436 32788
rect 23492 32732 24108 32788
rect 24164 32732 25452 32788
rect 25508 32732 25518 32788
rect 26646 32732 26684 32788
rect 26740 32732 26750 32788
rect 32498 32732 32508 32788
rect 32564 32732 38668 32788
rect 40338 32732 40348 32788
rect 40404 32732 41468 32788
rect 41524 32732 41534 32788
rect 3042 32620 3052 32676
rect 3108 32620 3388 32676
rect 3444 32620 3836 32676
rect 3892 32620 3902 32676
rect 5058 32620 5068 32676
rect 5124 32620 5964 32676
rect 6020 32620 6030 32676
rect 6962 32620 6972 32676
rect 7028 32620 11004 32676
rect 11060 32620 11070 32676
rect 16706 32620 16716 32676
rect 16772 32620 27916 32676
rect 27972 32620 27982 32676
rect 29586 32620 29596 32676
rect 29652 32620 30716 32676
rect 30772 32620 30782 32676
rect 35074 32620 35084 32676
rect 35140 32620 36428 32676
rect 36484 32620 36494 32676
rect 38612 32564 38668 32732
rect 40226 32620 40236 32676
rect 40292 32620 40908 32676
rect 40964 32620 40974 32676
rect 2818 32508 2828 32564
rect 2884 32508 3388 32564
rect 3332 32452 3388 32508
rect 6188 32508 12684 32564
rect 12740 32508 15260 32564
rect 15316 32508 15326 32564
rect 16370 32508 16380 32564
rect 16436 32508 17500 32564
rect 17556 32508 17566 32564
rect 22082 32508 22092 32564
rect 22148 32508 22428 32564
rect 22484 32508 22494 32564
rect 28690 32508 28700 32564
rect 28756 32508 29148 32564
rect 29204 32508 29214 32564
rect 38612 32508 39844 32564
rect 40002 32508 40012 32564
rect 40068 32508 41132 32564
rect 41188 32508 41198 32564
rect 6188 32452 6244 32508
rect 39788 32452 39844 32508
rect 3332 32396 3948 32452
rect 4004 32396 6244 32452
rect 10882 32396 10892 32452
rect 10948 32396 12572 32452
rect 12628 32396 12638 32452
rect 14914 32396 14924 32452
rect 14980 32396 15148 32452
rect 19394 32396 19404 32452
rect 19460 32396 21644 32452
rect 21700 32396 21710 32452
rect 34178 32396 34188 32452
rect 34244 32396 35980 32452
rect 36036 32396 37100 32452
rect 37156 32396 37166 32452
rect 37874 32396 37884 32452
rect 37940 32396 38220 32452
rect 38276 32396 39340 32452
rect 39396 32396 39406 32452
rect 39788 32396 40572 32452
rect 40628 32396 40638 32452
rect 14466 32284 14476 32340
rect 14532 32284 14924 32340
rect 14980 32284 14990 32340
rect 15092 32228 15148 32396
rect 49200 32340 50000 32368
rect 15586 32284 15596 32340
rect 15652 32284 23324 32340
rect 23380 32284 23390 32340
rect 26674 32284 26684 32340
rect 26740 32284 27020 32340
rect 27076 32284 27086 32340
rect 48066 32284 48076 32340
rect 48132 32284 50000 32340
rect 49200 32256 50000 32284
rect 2034 32172 2044 32228
rect 2100 32172 2604 32228
rect 2660 32172 2670 32228
rect 8390 32172 8428 32228
rect 8484 32172 8494 32228
rect 15092 32172 24892 32228
rect 24948 32172 25676 32228
rect 25732 32172 25742 32228
rect 27458 32172 27468 32228
rect 27524 32172 27804 32228
rect 27860 32172 27870 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 2258 32060 2268 32116
rect 2324 32060 3388 32116
rect 3444 32060 3948 32116
rect 4004 32060 4014 32116
rect 8502 32060 8540 32116
rect 8596 32060 8606 32116
rect 9762 32060 9772 32116
rect 9828 32060 10892 32116
rect 10948 32060 10958 32116
rect 18722 32060 18732 32116
rect 18788 32060 20636 32116
rect 20692 32060 20702 32116
rect 2482 31948 2492 32004
rect 2548 31948 3164 32004
rect 3220 31948 3230 32004
rect 4834 31948 4844 32004
rect 4900 31948 8764 32004
rect 8820 31948 8830 32004
rect 9426 31948 9436 32004
rect 9492 31948 9502 32004
rect 10994 31948 11004 32004
rect 11060 31948 11788 32004
rect 11844 31948 11854 32004
rect 18162 31948 18172 32004
rect 18228 31948 22988 32004
rect 23044 31948 23054 32004
rect 38546 31948 38556 32004
rect 38612 31948 40012 32004
rect 40068 31948 40078 32004
rect 9436 31892 9492 31948
rect 1698 31836 1708 31892
rect 1764 31836 8988 31892
rect 9044 31836 9054 31892
rect 9436 31836 11340 31892
rect 11396 31836 11406 31892
rect 13234 31836 13244 31892
rect 13300 31836 14476 31892
rect 14532 31836 14542 31892
rect 18050 31836 18060 31892
rect 18116 31836 22652 31892
rect 22708 31836 23100 31892
rect 23156 31836 23166 31892
rect 24770 31836 24780 31892
rect 24836 31836 25564 31892
rect 25620 31836 25630 31892
rect 32610 31836 32620 31892
rect 32676 31836 37996 31892
rect 38052 31836 38062 31892
rect 38658 31836 38668 31892
rect 38724 31836 39340 31892
rect 39396 31836 39406 31892
rect 42242 31836 42252 31892
rect 42308 31836 44716 31892
rect 44772 31836 44782 31892
rect 45154 31836 45164 31892
rect 45220 31836 45836 31892
rect 45892 31836 45902 31892
rect 37996 31780 38052 31836
rect 2818 31724 2828 31780
rect 2884 31724 3612 31780
rect 3668 31724 3678 31780
rect 5954 31724 5964 31780
rect 6020 31724 7084 31780
rect 7140 31724 7150 31780
rect 8194 31724 8204 31780
rect 8260 31724 9436 31780
rect 9492 31724 9502 31780
rect 12450 31724 12460 31780
rect 12516 31724 14252 31780
rect 14308 31724 14318 31780
rect 14578 31724 14588 31780
rect 14644 31724 16156 31780
rect 16212 31724 16222 31780
rect 16594 31724 16604 31780
rect 16660 31724 17388 31780
rect 17444 31724 17454 31780
rect 19506 31724 19516 31780
rect 19572 31724 21196 31780
rect 21252 31724 21262 31780
rect 22642 31724 22652 31780
rect 22708 31724 24108 31780
rect 24164 31724 26460 31780
rect 26516 31724 26796 31780
rect 26852 31724 26862 31780
rect 27122 31724 27132 31780
rect 27188 31724 27198 31780
rect 33058 31724 33068 31780
rect 33124 31724 33516 31780
rect 33572 31724 33582 31780
rect 37996 31724 38668 31780
rect 42354 31724 42364 31780
rect 42420 31724 45276 31780
rect 45332 31724 45342 31780
rect 16604 31668 16660 31724
rect 27132 31668 27188 31724
rect 3154 31612 3164 31668
rect 3220 31612 3724 31668
rect 3780 31612 3790 31668
rect 4508 31612 4956 31668
rect 5012 31612 5852 31668
rect 5908 31612 5918 31668
rect 6066 31612 6076 31668
rect 6132 31612 6412 31668
rect 6468 31612 7196 31668
rect 7252 31612 7262 31668
rect 8838 31612 8876 31668
rect 8932 31612 8942 31668
rect 13122 31612 13132 31668
rect 13188 31612 13468 31668
rect 13524 31612 13692 31668
rect 13748 31612 13758 31668
rect 15586 31612 15596 31668
rect 15652 31612 16660 31668
rect 18162 31612 18172 31668
rect 18228 31612 21420 31668
rect 21476 31612 21486 31668
rect 23986 31612 23996 31668
rect 24052 31612 27188 31668
rect 28578 31612 28588 31668
rect 28644 31612 29148 31668
rect 29204 31612 30492 31668
rect 30548 31612 30558 31668
rect 34626 31612 34636 31668
rect 34692 31612 35644 31668
rect 35700 31612 35710 31668
rect 4508 31556 4564 31612
rect 38612 31556 38668 31724
rect 44370 31612 44380 31668
rect 44436 31612 45612 31668
rect 45668 31612 45678 31668
rect 2370 31500 2380 31556
rect 2436 31500 2446 31556
rect 2594 31500 2604 31556
rect 2660 31500 3836 31556
rect 3892 31500 3902 31556
rect 4498 31500 4508 31556
rect 4564 31500 4574 31556
rect 4722 31500 4732 31556
rect 4788 31500 4798 31556
rect 6850 31500 6860 31556
rect 6916 31500 7420 31556
rect 7476 31500 7486 31556
rect 9874 31500 9884 31556
rect 9940 31500 11564 31556
rect 11620 31500 11630 31556
rect 15092 31500 18060 31556
rect 18116 31500 18126 31556
rect 19282 31500 19292 31556
rect 19348 31500 20636 31556
rect 20692 31500 20702 31556
rect 22530 31500 22540 31556
rect 22596 31500 25228 31556
rect 25284 31500 25294 31556
rect 29250 31500 29260 31556
rect 29316 31500 30380 31556
rect 30436 31500 30446 31556
rect 38210 31500 38220 31556
rect 38276 31500 38286 31556
rect 38612 31500 38780 31556
rect 38836 31500 39340 31556
rect 39396 31500 39406 31556
rect 41570 31500 41580 31556
rect 41636 31500 42700 31556
rect 42756 31500 42766 31556
rect 43922 31500 43932 31556
rect 43988 31500 44828 31556
rect 44884 31500 46172 31556
rect 46228 31500 46238 31556
rect 2380 31444 2436 31500
rect 4732 31444 4788 31500
rect 15092 31444 15148 31500
rect 38220 31444 38276 31500
rect 2380 31388 3276 31444
rect 3332 31388 4788 31444
rect 5058 31388 5068 31444
rect 5124 31388 5292 31444
rect 5348 31388 7196 31444
rect 7252 31388 15148 31444
rect 18162 31388 18172 31444
rect 18228 31388 19516 31444
rect 19572 31388 19582 31444
rect 20290 31388 20300 31444
rect 20356 31388 20748 31444
rect 20804 31388 20814 31444
rect 25554 31388 25564 31444
rect 25620 31388 33180 31444
rect 33236 31388 33740 31444
rect 33796 31388 33806 31444
rect 38220 31388 38668 31444
rect 38724 31388 38734 31444
rect 44930 31388 44940 31444
rect 44996 31388 45612 31444
rect 45668 31388 46620 31444
rect 46676 31388 46686 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 3378 31276 3388 31332
rect 3444 31276 4508 31332
rect 4564 31276 4574 31332
rect 7522 31276 7532 31332
rect 7588 31276 10332 31332
rect 10388 31276 10398 31332
rect 11330 31276 11340 31332
rect 11396 31276 13580 31332
rect 13636 31276 13646 31332
rect 22306 31276 22316 31332
rect 22372 31276 22876 31332
rect 22932 31276 22942 31332
rect 28914 31276 28924 31332
rect 28980 31276 38668 31332
rect 38612 31220 38668 31276
rect 2146 31164 2156 31220
rect 2212 31164 4060 31220
rect 4116 31164 4126 31220
rect 6066 31164 6076 31220
rect 6132 31164 6524 31220
rect 6580 31164 6590 31220
rect 7858 31164 7868 31220
rect 7924 31164 10220 31220
rect 10276 31164 10286 31220
rect 17154 31164 17164 31220
rect 17220 31164 23996 31220
rect 24052 31164 24062 31220
rect 30146 31164 30156 31220
rect 30212 31164 31612 31220
rect 31668 31164 31678 31220
rect 31826 31164 31836 31220
rect 31892 31164 34860 31220
rect 34916 31164 34926 31220
rect 38612 31164 40348 31220
rect 40404 31164 40414 31220
rect 4386 31052 4396 31108
rect 4452 31052 6860 31108
rect 6916 31052 6926 31108
rect 8978 31052 8988 31108
rect 9044 31052 9660 31108
rect 9716 31052 12124 31108
rect 12180 31052 13244 31108
rect 13300 31052 13310 31108
rect 14466 31052 14476 31108
rect 14532 31052 16156 31108
rect 16212 31052 16222 31108
rect 22418 31052 22428 31108
rect 22484 31052 22988 31108
rect 23044 31052 23054 31108
rect 30482 31052 30492 31108
rect 30548 31052 33068 31108
rect 33124 31052 33134 31108
rect 34514 31052 34524 31108
rect 34580 31052 35756 31108
rect 35812 31052 35822 31108
rect 46386 31052 46396 31108
rect 46452 31052 47404 31108
rect 47460 31052 47470 31108
rect 46396 30996 46452 31052
rect 5170 30940 5180 30996
rect 5236 30940 5292 30996
rect 5348 30940 5358 30996
rect 6514 30940 6524 30996
rect 6580 30940 6972 30996
rect 7028 30940 8204 30996
rect 8260 30940 8270 30996
rect 14914 30940 14924 30996
rect 14980 30940 15372 30996
rect 15428 30940 15820 30996
rect 15876 30940 18732 30996
rect 18788 30940 19740 30996
rect 19796 30940 28700 30996
rect 28756 30940 28766 30996
rect 30818 30940 30828 30996
rect 30884 30940 33180 30996
rect 33236 30940 33246 30996
rect 34850 30940 34860 30996
rect 34916 30940 35868 30996
rect 35924 30940 35934 30996
rect 45042 30940 45052 30996
rect 45108 30940 45836 30996
rect 45892 30940 45902 30996
rect 46162 30940 46172 30996
rect 46228 30940 46452 30996
rect 17490 30828 17500 30884
rect 17556 30828 18396 30884
rect 18452 30828 20076 30884
rect 20132 30828 20142 30884
rect 22418 30828 22428 30884
rect 22484 30828 25340 30884
rect 25396 30828 25406 30884
rect 27570 30828 27580 30884
rect 27636 30828 28252 30884
rect 28308 30828 28318 30884
rect 31826 30828 31836 30884
rect 31892 30828 33852 30884
rect 33908 30828 33918 30884
rect 6514 30716 6524 30772
rect 6580 30716 8428 30772
rect 8484 30716 8494 30772
rect 9426 30716 9436 30772
rect 9492 30716 11564 30772
rect 11620 30716 13692 30772
rect 13748 30716 13758 30772
rect 16258 30716 16268 30772
rect 16324 30716 17276 30772
rect 17332 30716 17342 30772
rect 17938 30716 17948 30772
rect 18004 30716 18014 30772
rect 21494 30716 21532 30772
rect 21588 30716 21598 30772
rect 23986 30716 23996 30772
rect 24052 30716 24444 30772
rect 24500 30716 24510 30772
rect 26002 30716 26012 30772
rect 26068 30716 26078 30772
rect 30370 30716 30380 30772
rect 30436 30716 31388 30772
rect 31444 30716 33292 30772
rect 33348 30716 33358 30772
rect 41010 30716 41020 30772
rect 41076 30716 43932 30772
rect 43988 30716 46956 30772
rect 47012 30716 47022 30772
rect 17948 30660 18004 30716
rect 26012 30660 26068 30716
rect 12226 30604 12236 30660
rect 12292 30604 18004 30660
rect 18386 30604 18396 30660
rect 18452 30604 21644 30660
rect 21700 30604 21710 30660
rect 24098 30604 24108 30660
rect 24164 30604 25340 30660
rect 25396 30604 26068 30660
rect 43362 30604 43372 30660
rect 43428 30604 47628 30660
rect 47684 30604 47694 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 17938 30492 17948 30548
rect 18004 30492 21868 30548
rect 21924 30492 21934 30548
rect 22316 30492 23772 30548
rect 23828 30492 23838 30548
rect 37538 30492 37548 30548
rect 37604 30492 38668 30548
rect 42802 30492 42812 30548
rect 42868 30492 43596 30548
rect 43652 30492 43662 30548
rect 22316 30436 22372 30492
rect 38612 30436 38668 30492
rect 9538 30380 9548 30436
rect 9604 30380 10332 30436
rect 10388 30380 10398 30436
rect 12898 30380 12908 30436
rect 12964 30380 13468 30436
rect 13524 30380 13534 30436
rect 15250 30380 15260 30436
rect 15316 30380 16940 30436
rect 16996 30380 17006 30436
rect 18498 30380 18508 30436
rect 18564 30380 22372 30436
rect 25862 30380 25900 30436
rect 25956 30380 25966 30436
rect 36418 30380 36428 30436
rect 36484 30380 37100 30436
rect 37156 30380 37884 30436
rect 37940 30380 37950 30436
rect 38612 30380 40124 30436
rect 40180 30380 40190 30436
rect 46386 30380 46396 30436
rect 46452 30380 47628 30436
rect 47684 30380 47694 30436
rect 1922 30268 1932 30324
rect 1988 30268 3724 30324
rect 3780 30268 3790 30324
rect 4946 30268 4956 30324
rect 5012 30268 5068 30324
rect 5124 30268 6076 30324
rect 6132 30268 6142 30324
rect 15138 30268 15148 30324
rect 15204 30268 16604 30324
rect 16660 30268 17836 30324
rect 17892 30268 17902 30324
rect 19058 30268 19068 30324
rect 19124 30268 19628 30324
rect 19684 30268 19852 30324
rect 19908 30268 19918 30324
rect 20290 30268 20300 30324
rect 20356 30268 22652 30324
rect 22708 30268 22718 30324
rect 23762 30268 23772 30324
rect 23828 30268 23996 30324
rect 24052 30268 24062 30324
rect 35746 30268 35756 30324
rect 35812 30268 36092 30324
rect 36148 30268 36158 30324
rect 37314 30268 37324 30324
rect 37380 30268 38556 30324
rect 38612 30268 39788 30324
rect 39844 30268 39854 30324
rect 43922 30268 43932 30324
rect 43988 30268 45164 30324
rect 45220 30268 46508 30324
rect 46564 30268 46574 30324
rect 2930 30156 2940 30212
rect 2996 30156 3388 30212
rect 3444 30156 4284 30212
rect 4340 30156 4350 30212
rect 4834 30156 4844 30212
rect 4900 30156 5852 30212
rect 5908 30156 6636 30212
rect 6692 30156 7084 30212
rect 7140 30156 7150 30212
rect 8866 30156 8876 30212
rect 8932 30156 9212 30212
rect 9268 30156 9278 30212
rect 9650 30156 9660 30212
rect 9716 30156 10556 30212
rect 10612 30156 12460 30212
rect 12516 30156 12526 30212
rect 15922 30156 15932 30212
rect 15988 30156 16268 30212
rect 16324 30156 16334 30212
rect 16482 30156 16492 30212
rect 16548 30156 16586 30212
rect 21270 30156 21308 30212
rect 21364 30156 21374 30212
rect 22306 30156 22316 30212
rect 22372 30156 23548 30212
rect 23604 30156 23614 30212
rect 28690 30156 28700 30212
rect 28756 30156 34188 30212
rect 34244 30156 34254 30212
rect 36978 30156 36988 30212
rect 37044 30156 40796 30212
rect 40852 30156 41468 30212
rect 41524 30156 41534 30212
rect 43250 30156 43260 30212
rect 43316 30156 43820 30212
rect 43876 30156 43886 30212
rect 44930 30156 44940 30212
rect 44996 30156 45612 30212
rect 45668 30156 46060 30212
rect 46116 30156 47068 30212
rect 47124 30156 47134 30212
rect 1820 30044 2044 30100
rect 2100 30044 2268 30100
rect 2324 30044 2334 30100
rect 4050 30044 4060 30100
rect 4116 30044 4172 30100
rect 4228 30044 4238 30100
rect 10994 30044 11004 30100
rect 11060 30044 17500 30100
rect 17556 30044 17566 30100
rect 18806 30044 18844 30100
rect 18900 30044 18910 30100
rect 19068 30044 29260 30100
rect 29316 30044 29326 30100
rect 1820 29876 1876 30044
rect 19068 29988 19124 30044
rect 14130 29932 14140 29988
rect 14196 29932 19124 29988
rect 20850 29932 20860 29988
rect 20916 29932 21532 29988
rect 21588 29932 21598 29988
rect 23202 29932 23212 29988
rect 23268 29932 24220 29988
rect 24276 29932 24286 29988
rect 29586 29932 29596 29988
rect 29652 29932 32060 29988
rect 32116 29932 32126 29988
rect 45042 29932 45052 29988
rect 45108 29932 48076 29988
rect 48132 29932 48142 29988
rect 1810 29820 1820 29876
rect 1876 29820 1886 29876
rect 8866 29820 8876 29876
rect 8932 29820 9772 29876
rect 9828 29820 9838 29876
rect 11890 29820 11900 29876
rect 11956 29820 13244 29876
rect 13300 29820 14812 29876
rect 14868 29820 15820 29876
rect 15876 29820 15886 29876
rect 17378 29820 17388 29876
rect 17444 29820 18732 29876
rect 18788 29820 18798 29876
rect 20626 29820 20636 29876
rect 20692 29820 21308 29876
rect 21364 29820 21374 29876
rect 37212 29820 38332 29876
rect 38388 29820 39900 29876
rect 39956 29820 39966 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 6626 29708 6636 29764
rect 6692 29708 10220 29764
rect 10276 29708 11340 29764
rect 11396 29708 11406 29764
rect 12338 29708 12348 29764
rect 12404 29708 13916 29764
rect 13972 29708 13982 29764
rect 23398 29708 23436 29764
rect 23492 29708 24108 29764
rect 24164 29708 24174 29764
rect 28588 29708 29708 29764
rect 29764 29708 30940 29764
rect 30996 29708 31500 29764
rect 31556 29708 32284 29764
rect 32340 29708 32350 29764
rect 28588 29652 28644 29708
rect 10546 29596 10556 29652
rect 10612 29596 10724 29652
rect 11778 29596 11788 29652
rect 11844 29596 12684 29652
rect 12740 29596 12750 29652
rect 12898 29596 12908 29652
rect 12964 29596 28588 29652
rect 28644 29596 28654 29652
rect 29148 29596 34524 29652
rect 34580 29596 34972 29652
rect 35028 29596 35038 29652
rect 2034 29484 2044 29540
rect 2100 29484 5292 29540
rect 5348 29484 5358 29540
rect 8390 29484 8428 29540
rect 8484 29484 8494 29540
rect 9874 29484 9884 29540
rect 9940 29484 10444 29540
rect 10500 29484 10510 29540
rect 6066 29372 6076 29428
rect 6132 29372 8988 29428
rect 9044 29372 9548 29428
rect 9604 29372 9614 29428
rect 4834 29260 4844 29316
rect 4900 29260 5460 29316
rect 8502 29260 8540 29316
rect 8596 29260 8606 29316
rect 4722 29148 4732 29204
rect 4788 29148 4900 29204
rect 5030 29148 5068 29204
rect 5124 29148 5134 29204
rect 1922 29036 1932 29092
rect 1988 29036 2380 29092
rect 2436 29036 2446 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 4844 28868 4900 29148
rect 5404 29092 5460 29260
rect 10668 29204 10724 29596
rect 29148 29540 29204 29596
rect 13542 29484 13580 29540
rect 13636 29484 13646 29540
rect 17910 29484 17948 29540
rect 18004 29484 18014 29540
rect 20374 29484 20412 29540
rect 20468 29484 20478 29540
rect 27906 29484 27916 29540
rect 27972 29484 29148 29540
rect 29204 29484 29214 29540
rect 30146 29484 30156 29540
rect 30212 29484 30380 29540
rect 30436 29484 31052 29540
rect 31108 29484 31118 29540
rect 37212 29428 37268 29820
rect 40002 29484 40012 29540
rect 40068 29484 41356 29540
rect 41412 29484 41422 29540
rect 42242 29484 42252 29540
rect 42308 29484 43372 29540
rect 43428 29484 45388 29540
rect 45444 29484 45454 29540
rect 46050 29484 46060 29540
rect 46116 29484 46284 29540
rect 46340 29484 46620 29540
rect 46676 29484 46686 29540
rect 12338 29372 12348 29428
rect 12404 29372 17612 29428
rect 17668 29372 17678 29428
rect 17826 29372 17836 29428
rect 17892 29372 18396 29428
rect 18452 29372 18462 29428
rect 18946 29372 18956 29428
rect 19012 29372 20748 29428
rect 20804 29372 20814 29428
rect 21756 29372 27132 29428
rect 27188 29372 27198 29428
rect 27458 29372 27468 29428
rect 27524 29372 28588 29428
rect 28644 29372 28812 29428
rect 28868 29372 28878 29428
rect 30818 29372 30828 29428
rect 30884 29372 31612 29428
rect 31668 29372 33180 29428
rect 33236 29372 33246 29428
rect 33730 29372 33740 29428
rect 33796 29372 37212 29428
rect 37268 29372 37278 29428
rect 39554 29372 39564 29428
rect 39620 29372 40236 29428
rect 40292 29372 41244 29428
rect 41300 29372 41310 29428
rect 45826 29372 45836 29428
rect 45892 29372 47068 29428
rect 47124 29372 47134 29428
rect 21756 29316 21812 29372
rect 19842 29260 19852 29316
rect 19908 29260 20636 29316
rect 20692 29260 20702 29316
rect 21746 29260 21756 29316
rect 21812 29260 21822 29316
rect 25666 29260 25676 29316
rect 25732 29260 26572 29316
rect 26628 29260 28140 29316
rect 28196 29260 28206 29316
rect 31826 29260 31836 29316
rect 31892 29260 38668 29316
rect 41682 29260 41692 29316
rect 41748 29260 42700 29316
rect 42756 29260 42766 29316
rect 44482 29260 44492 29316
rect 44548 29260 48188 29316
rect 48244 29260 48254 29316
rect 38612 29204 38668 29260
rect 5590 29148 5628 29204
rect 5684 29148 5694 29204
rect 10658 29148 10668 29204
rect 10724 29148 10734 29204
rect 19282 29148 19292 29204
rect 19348 29148 20300 29204
rect 20356 29148 21420 29204
rect 21476 29148 23436 29204
rect 23492 29148 27692 29204
rect 27748 29148 27758 29204
rect 38612 29148 38780 29204
rect 38836 29148 42140 29204
rect 42196 29148 42588 29204
rect 42644 29148 42654 29204
rect 5404 29036 10332 29092
rect 10388 29036 11004 29092
rect 11060 29036 11070 29092
rect 19506 29036 19516 29092
rect 19572 29036 20188 29092
rect 20244 29036 21196 29092
rect 21252 29036 21262 29092
rect 23090 29036 23100 29092
rect 23156 29036 24668 29092
rect 24724 29036 24734 29092
rect 36978 29036 36988 29092
rect 37044 29036 38108 29092
rect 38164 29036 38174 29092
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 5842 28924 5852 28980
rect 5908 28924 13692 28980
rect 13748 28924 15484 28980
rect 15540 28924 16940 28980
rect 16996 28924 17006 28980
rect 26198 28924 26236 28980
rect 26292 28924 26302 28980
rect 29922 28924 29932 28980
rect 29988 28924 31388 28980
rect 31444 28924 32844 28980
rect 32900 28924 32910 28980
rect 36418 28924 36428 28980
rect 36484 28924 36876 28980
rect 36932 28924 37436 28980
rect 37492 28924 37502 28980
rect 39228 28924 42252 28980
rect 42308 28924 43596 28980
rect 43652 28924 43662 28980
rect 39228 28868 39284 28924
rect 2482 28812 2492 28868
rect 2548 28812 4508 28868
rect 4564 28812 4900 28868
rect 6066 28812 6076 28868
rect 6132 28812 8540 28868
rect 8596 28812 8606 28868
rect 11218 28812 11228 28868
rect 11284 28812 11676 28868
rect 11732 28812 15932 28868
rect 15988 28812 15998 28868
rect 17836 28812 18172 28868
rect 18228 28812 18238 28868
rect 18386 28812 18396 28868
rect 18452 28812 18508 28868
rect 18564 28812 18574 28868
rect 19058 28812 19068 28868
rect 19124 28812 21644 28868
rect 21700 28812 21710 28868
rect 24210 28812 24220 28868
rect 24276 28812 27580 28868
rect 27636 28812 27646 28868
rect 28130 28812 28140 28868
rect 28196 28812 29484 28868
rect 29540 28812 29550 28868
rect 31042 28812 31052 28868
rect 31108 28812 31948 28868
rect 32004 28812 32014 28868
rect 34738 28812 34748 28868
rect 34804 28812 36316 28868
rect 36372 28812 36382 28868
rect 38546 28812 38556 28868
rect 38612 28812 39228 28868
rect 39284 28812 39294 28868
rect 40450 28812 40460 28868
rect 40516 28812 41468 28868
rect 41524 28812 42700 28868
rect 42756 28812 42766 28868
rect 44034 28812 44044 28868
rect 44100 28812 44716 28868
rect 44772 28812 46172 28868
rect 46228 28812 46238 28868
rect 17836 28756 17892 28812
rect 2146 28700 2156 28756
rect 2212 28700 4956 28756
rect 5012 28700 6300 28756
rect 6356 28700 7084 28756
rect 7140 28700 7150 28756
rect 7298 28700 7308 28756
rect 7364 28700 8092 28756
rect 8148 28700 9212 28756
rect 9268 28700 10556 28756
rect 10612 28700 10622 28756
rect 13570 28700 13580 28756
rect 13636 28700 17892 28756
rect 18050 28700 18060 28756
rect 18116 28700 18620 28756
rect 18676 28700 18686 28756
rect 19954 28700 19964 28756
rect 20020 28700 22764 28756
rect 22820 28700 22830 28756
rect 23986 28700 23996 28756
rect 24052 28700 25340 28756
rect 25396 28700 25406 28756
rect 28466 28700 28476 28756
rect 28532 28700 29876 28756
rect 30370 28700 30380 28756
rect 30436 28700 31612 28756
rect 31668 28700 31678 28756
rect 36530 28700 36540 28756
rect 36596 28700 37436 28756
rect 37492 28700 37502 28756
rect 41234 28700 41244 28756
rect 41300 28700 43484 28756
rect 43540 28700 43932 28756
rect 43988 28700 43998 28756
rect 29820 28644 29876 28700
rect 1698 28588 1708 28644
rect 1764 28588 4284 28644
rect 4340 28588 6076 28644
rect 6132 28588 6142 28644
rect 6300 28588 6524 28644
rect 6580 28588 6590 28644
rect 8540 28588 8988 28644
rect 9044 28588 9054 28644
rect 18386 28588 18396 28644
rect 18452 28588 18844 28644
rect 18900 28588 18910 28644
rect 24098 28588 24108 28644
rect 24164 28588 26684 28644
rect 26740 28588 26750 28644
rect 27122 28588 27132 28644
rect 27188 28588 29372 28644
rect 29428 28588 29438 28644
rect 29810 28588 29820 28644
rect 29876 28588 33068 28644
rect 33124 28588 33134 28644
rect 35858 28588 35868 28644
rect 35924 28588 37100 28644
rect 37156 28588 37166 28644
rect 41346 28588 41356 28644
rect 41412 28588 42812 28644
rect 42868 28588 42878 28644
rect 43250 28588 43260 28644
rect 43316 28588 44940 28644
rect 44996 28588 45006 28644
rect 6300 28532 6356 28588
rect 1810 28476 1820 28532
rect 1876 28476 2604 28532
rect 2660 28476 4508 28532
rect 4564 28476 4574 28532
rect 5058 28476 5068 28532
rect 5124 28476 6356 28532
rect 8540 28420 8596 28588
rect 41916 28532 41972 28588
rect 9874 28476 9884 28532
rect 9940 28476 11116 28532
rect 11172 28476 11182 28532
rect 15250 28476 15260 28532
rect 15316 28476 19404 28532
rect 19460 28476 20076 28532
rect 20132 28476 20142 28532
rect 26226 28476 26236 28532
rect 26292 28476 26908 28532
rect 26964 28476 26974 28532
rect 29250 28476 29260 28532
rect 29316 28476 34412 28532
rect 34468 28476 34478 28532
rect 35298 28476 35308 28532
rect 35364 28476 36988 28532
rect 37044 28476 37054 28532
rect 41906 28476 41916 28532
rect 41972 28476 41982 28532
rect 6962 28364 6972 28420
rect 7028 28364 7038 28420
rect 8530 28364 8540 28420
rect 8596 28364 8606 28420
rect 10658 28364 10668 28420
rect 10724 28364 18060 28420
rect 18116 28364 18126 28420
rect 18722 28364 18732 28420
rect 18788 28364 20356 28420
rect 20514 28364 20524 28420
rect 20580 28364 21084 28420
rect 21140 28364 22204 28420
rect 22260 28364 22270 28420
rect 22418 28364 22428 28420
rect 22484 28364 22522 28420
rect 28354 28364 28364 28420
rect 28420 28364 29148 28420
rect 29204 28364 29214 28420
rect 35746 28364 35756 28420
rect 35812 28364 36764 28420
rect 36820 28364 37212 28420
rect 37268 28364 37278 28420
rect 38210 28364 38220 28420
rect 38276 28364 39004 28420
rect 39060 28364 39070 28420
rect 6972 28308 7028 28364
rect 20300 28308 20356 28364
rect 1586 28252 1596 28308
rect 1652 28252 5180 28308
rect 5236 28252 5246 28308
rect 6972 28252 16492 28308
rect 16548 28252 16558 28308
rect 17938 28252 17948 28308
rect 18004 28252 19180 28308
rect 19236 28252 19246 28308
rect 20300 28252 25340 28308
rect 25396 28252 25406 28308
rect 28914 28252 28924 28308
rect 28980 28252 43260 28308
rect 43316 28252 43326 28308
rect 5180 28084 5236 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 5506 28140 5516 28196
rect 5572 28140 6076 28196
rect 6132 28140 6142 28196
rect 7970 28140 7980 28196
rect 8036 28140 9212 28196
rect 9268 28140 9278 28196
rect 10098 28140 10108 28196
rect 10164 28140 10174 28196
rect 11330 28140 11340 28196
rect 11396 28140 12908 28196
rect 12964 28140 12974 28196
rect 19030 28140 19068 28196
rect 19124 28140 19134 28196
rect 20514 28140 20524 28196
rect 20580 28140 21532 28196
rect 21588 28140 22540 28196
rect 22596 28140 22606 28196
rect 35522 28140 35532 28196
rect 35588 28140 36428 28196
rect 36484 28140 36494 28196
rect 37202 28140 37212 28196
rect 37268 28140 38444 28196
rect 38500 28140 41804 28196
rect 41860 28140 41870 28196
rect 10108 28084 10164 28140
rect 1810 28028 1820 28084
rect 1876 28028 2604 28084
rect 2660 28028 2670 28084
rect 5180 28028 8148 28084
rect 8306 28028 8316 28084
rect 8372 28028 10164 28084
rect 11218 28028 11228 28084
rect 11284 28028 27804 28084
rect 27860 28028 27870 28084
rect 39330 28028 39340 28084
rect 39396 28028 40124 28084
rect 40180 28028 40190 28084
rect 41010 28028 41020 28084
rect 41076 28028 42364 28084
rect 42420 28028 44492 28084
rect 44548 28028 44558 28084
rect 4834 27916 4844 27972
rect 4900 27916 6748 27972
rect 6804 27916 7644 27972
rect 7700 27916 7710 27972
rect 8092 27860 8148 28028
rect 8642 27916 8652 27972
rect 8708 27916 10108 27972
rect 10164 27916 10780 27972
rect 10836 27916 10846 27972
rect 11778 27916 11788 27972
rect 11844 27916 14252 27972
rect 14308 27916 14318 27972
rect 17154 27916 17164 27972
rect 17220 27916 17724 27972
rect 17780 27916 17790 27972
rect 19058 27916 19068 27972
rect 19124 27916 21420 27972
rect 21476 27916 21486 27972
rect 24098 27916 24108 27972
rect 24164 27916 27244 27972
rect 27300 27916 29428 27972
rect 33394 27916 33404 27972
rect 33460 27916 34076 27972
rect 34132 27916 34142 27972
rect 29372 27860 29428 27916
rect 3490 27804 3500 27860
rect 3556 27804 4172 27860
rect 4228 27804 7532 27860
rect 7588 27804 7598 27860
rect 8092 27804 9660 27860
rect 9716 27804 9726 27860
rect 11732 27804 14140 27860
rect 14196 27804 15148 27860
rect 15204 27804 15214 27860
rect 18610 27804 18620 27860
rect 18676 27804 18844 27860
rect 18900 27804 23212 27860
rect 23268 27804 24444 27860
rect 24500 27804 24510 27860
rect 25330 27804 25340 27860
rect 25396 27804 26796 27860
rect 26852 27804 26862 27860
rect 27570 27804 27580 27860
rect 27636 27804 28140 27860
rect 28196 27804 28206 27860
rect 29362 27804 29372 27860
rect 29428 27804 29820 27860
rect 29876 27804 29886 27860
rect 45826 27804 45836 27860
rect 45892 27804 47516 27860
rect 47572 27804 47582 27860
rect 11732 27748 11788 27804
rect 7410 27692 7420 27748
rect 7476 27692 11788 27748
rect 15474 27692 15484 27748
rect 15540 27692 17276 27748
rect 17332 27692 17342 27748
rect 18470 27692 18508 27748
rect 18564 27692 18574 27748
rect 19404 27692 20636 27748
rect 20692 27692 20860 27748
rect 20916 27692 20926 27748
rect 21186 27692 21196 27748
rect 21252 27692 22428 27748
rect 22484 27692 22494 27748
rect 24210 27692 24220 27748
rect 24276 27692 24286 27748
rect 33506 27692 33516 27748
rect 33572 27692 34300 27748
rect 34356 27692 34366 27748
rect 19404 27636 19460 27692
rect 24220 27636 24276 27692
rect 5170 27580 5180 27636
rect 5236 27580 7532 27636
rect 7588 27580 7598 27636
rect 16930 27580 16940 27636
rect 16996 27580 19460 27636
rect 19618 27580 19628 27636
rect 19684 27580 24276 27636
rect 26450 27580 26460 27636
rect 26516 27580 27020 27636
rect 27076 27580 27086 27636
rect 45266 27580 45276 27636
rect 45332 27580 45500 27636
rect 45556 27580 47068 27636
rect 47124 27580 47134 27636
rect 9650 27468 9660 27524
rect 9716 27468 11340 27524
rect 11396 27468 13580 27524
rect 13636 27468 13646 27524
rect 20626 27468 20636 27524
rect 20692 27468 21084 27524
rect 21140 27468 21150 27524
rect 34598 27468 34636 27524
rect 34692 27468 34702 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 49200 27412 50000 27440
rect 13010 27356 13020 27412
rect 13076 27356 13356 27412
rect 13412 27356 13422 27412
rect 22194 27356 22204 27412
rect 22260 27356 28364 27412
rect 28420 27356 28430 27412
rect 45490 27356 45500 27412
rect 45556 27356 47852 27412
rect 47908 27356 47918 27412
rect 48178 27356 48188 27412
rect 48244 27356 50000 27412
rect 49200 27328 50000 27356
rect 20748 27244 23996 27300
rect 24052 27244 24062 27300
rect 20748 27188 20804 27244
rect 5058 27132 5068 27188
rect 5124 27132 6860 27188
rect 6916 27132 6926 27188
rect 12674 27132 12684 27188
rect 12740 27132 17724 27188
rect 17780 27132 17790 27188
rect 18162 27132 18172 27188
rect 18228 27132 19180 27188
rect 19236 27132 20188 27188
rect 20244 27132 20804 27188
rect 23762 27132 23772 27188
rect 23828 27132 25116 27188
rect 25172 27132 27356 27188
rect 27412 27132 29148 27188
rect 29204 27132 29708 27188
rect 29764 27132 29774 27188
rect 32162 27132 32172 27188
rect 32228 27132 33404 27188
rect 33460 27132 33470 27188
rect 42130 27132 42140 27188
rect 42196 27132 42812 27188
rect 42868 27132 42878 27188
rect 43698 27132 43708 27188
rect 43764 27132 44268 27188
rect 44324 27132 46508 27188
rect 46564 27132 46574 27188
rect 47058 27132 47068 27188
rect 47124 27132 48188 27188
rect 48244 27132 48254 27188
rect 5394 27020 5404 27076
rect 5460 27020 6972 27076
rect 7028 27020 8428 27076
rect 8484 27020 8494 27076
rect 10322 27020 10332 27076
rect 10388 27020 12236 27076
rect 12292 27020 12302 27076
rect 13010 27020 13020 27076
rect 13076 27020 17388 27076
rect 17444 27020 17454 27076
rect 18498 27020 18508 27076
rect 18564 27020 18844 27076
rect 18900 27020 18910 27076
rect 20066 27020 20076 27076
rect 20132 27020 21196 27076
rect 21252 27020 21262 27076
rect 22082 27020 22092 27076
rect 22148 27020 23100 27076
rect 23156 27020 25340 27076
rect 25396 27020 25406 27076
rect 27794 27020 27804 27076
rect 27860 27020 28252 27076
rect 28308 27020 28700 27076
rect 28756 27020 29484 27076
rect 29540 27020 29550 27076
rect 31826 27020 31836 27076
rect 31892 27020 31902 27076
rect 35074 27020 35084 27076
rect 35140 27020 37436 27076
rect 37492 27020 37502 27076
rect 20076 26964 20132 27020
rect 31836 26964 31892 27020
rect 5506 26908 5516 26964
rect 5572 26908 5964 26964
rect 6020 26908 7756 26964
rect 7812 26908 7822 26964
rect 12786 26908 12796 26964
rect 12852 26908 15708 26964
rect 15764 26908 15774 26964
rect 16818 26908 16828 26964
rect 16884 26908 20132 26964
rect 26796 26908 30604 26964
rect 30660 26908 31892 26964
rect 26796 26852 26852 26908
rect 3332 26796 17052 26852
rect 17108 26796 17118 26852
rect 20850 26796 20860 26852
rect 20916 26796 21532 26852
rect 21588 26796 21598 26852
rect 22866 26796 22876 26852
rect 22932 26796 26852 26852
rect 27458 26796 27468 26852
rect 27524 26796 31276 26852
rect 31332 26796 31342 26852
rect 3332 26740 3388 26796
rect 1474 26684 1484 26740
rect 1540 26684 3388 26740
rect 6038 26684 6076 26740
rect 6132 26684 6142 26740
rect 14578 26684 14588 26740
rect 14644 26684 15596 26740
rect 15652 26684 15662 26740
rect 15922 26684 15932 26740
rect 15988 26684 16604 26740
rect 16660 26684 16670 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 16146 26572 16156 26628
rect 16212 26572 16492 26628
rect 16548 26572 19068 26628
rect 19124 26572 19134 26628
rect 21532 26516 21588 26796
rect 26562 26684 26572 26740
rect 26628 26684 33964 26740
rect 34020 26684 34030 26740
rect 45826 26684 45836 26740
rect 45892 26684 46396 26740
rect 46452 26684 46462 26740
rect 26898 26572 26908 26628
rect 26964 26572 32844 26628
rect 32900 26572 32910 26628
rect 37202 26572 37212 26628
rect 37268 26572 38108 26628
rect 38164 26572 38668 26628
rect 4834 26460 4844 26516
rect 4900 26460 7196 26516
rect 7252 26460 7262 26516
rect 15810 26460 15820 26516
rect 15876 26460 16380 26516
rect 16436 26460 16446 26516
rect 18386 26460 18396 26516
rect 18452 26460 19404 26516
rect 19460 26460 19470 26516
rect 21532 26460 24332 26516
rect 24388 26460 25900 26516
rect 25956 26460 25966 26516
rect 26646 26460 26684 26516
rect 26740 26460 26750 26516
rect 28578 26460 28588 26516
rect 28644 26460 32060 26516
rect 32116 26460 36988 26516
rect 37044 26460 37054 26516
rect 38612 26460 38668 26572
rect 38724 26460 38734 26516
rect 6290 26348 6300 26404
rect 6356 26348 7308 26404
rect 7364 26348 7374 26404
rect 13346 26348 13356 26404
rect 13412 26348 14252 26404
rect 14308 26348 14318 26404
rect 15138 26348 15148 26404
rect 15204 26348 17500 26404
rect 17556 26348 17566 26404
rect 19506 26348 19516 26404
rect 19572 26348 23324 26404
rect 23380 26348 23390 26404
rect 26226 26348 26236 26404
rect 26292 26348 27468 26404
rect 27524 26348 29148 26404
rect 29204 26348 29214 26404
rect 38210 26348 38220 26404
rect 38276 26348 38892 26404
rect 38948 26348 38958 26404
rect 42354 26348 42364 26404
rect 42420 26348 43260 26404
rect 43316 26348 43326 26404
rect 45042 26348 45052 26404
rect 45108 26348 45612 26404
rect 45668 26348 45678 26404
rect 43260 26292 43316 26348
rect 1698 26236 1708 26292
rect 1764 26236 4620 26292
rect 4676 26236 5852 26292
rect 5908 26236 5918 26292
rect 6076 26236 11564 26292
rect 11620 26236 12348 26292
rect 12404 26236 12414 26292
rect 15092 26236 16156 26292
rect 16212 26236 16222 26292
rect 20514 26236 20524 26292
rect 20580 26236 22316 26292
rect 22372 26236 22382 26292
rect 29698 26236 29708 26292
rect 29764 26236 31836 26292
rect 31892 26236 33628 26292
rect 33684 26236 33694 26292
rect 35410 26236 35420 26292
rect 35476 26236 38444 26292
rect 38500 26236 39004 26292
rect 39060 26236 39070 26292
rect 43260 26236 45836 26292
rect 45892 26236 45902 26292
rect 6076 26180 6132 26236
rect 5730 26124 5740 26180
rect 5796 26124 6132 26180
rect 11330 26124 11340 26180
rect 11396 26124 12012 26180
rect 12068 26124 12460 26180
rect 12516 26124 12526 26180
rect 15092 26068 15148 26236
rect 21074 26124 21084 26180
rect 21140 26124 21420 26180
rect 21476 26124 21486 26180
rect 22082 26124 22092 26180
rect 22148 26124 23772 26180
rect 23828 26124 23838 26180
rect 25778 26124 25788 26180
rect 25844 26124 26572 26180
rect 26628 26124 26638 26180
rect 27234 26124 27244 26180
rect 27300 26124 27580 26180
rect 27636 26124 28028 26180
rect 28084 26124 28094 26180
rect 32834 26124 32844 26180
rect 32900 26124 34076 26180
rect 34132 26124 34142 26180
rect 34962 26124 34972 26180
rect 35028 26124 36428 26180
rect 36484 26124 39452 26180
rect 39508 26124 39518 26180
rect 40002 26124 40012 26180
rect 40068 26124 40796 26180
rect 40852 26124 40862 26180
rect 41010 26124 41020 26180
rect 41076 26124 41916 26180
rect 41972 26124 42140 26180
rect 42196 26124 42206 26180
rect 7074 26012 7084 26068
rect 7140 26012 8204 26068
rect 8260 26012 8270 26068
rect 10658 26012 10668 26068
rect 10724 26012 15148 26068
rect 17266 26012 17276 26068
rect 17332 26012 17836 26068
rect 17892 26012 17902 26068
rect 19142 26012 19180 26068
rect 19236 26012 20076 26068
rect 20132 26012 20142 26068
rect 34524 26012 35868 26068
rect 35924 26012 35934 26068
rect 19180 25956 19236 26012
rect 34524 25956 34580 26012
rect 10546 25900 10556 25956
rect 10612 25900 17332 25956
rect 17938 25900 17948 25956
rect 18004 25900 19236 25956
rect 19394 25900 19404 25956
rect 19460 25900 25004 25956
rect 25060 25900 28588 25956
rect 28644 25900 28654 25956
rect 30930 25900 30940 25956
rect 30996 25900 31836 25956
rect 31892 25900 34524 25956
rect 34580 25900 34590 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 17276 25844 17332 25900
rect 27244 25844 27300 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 13906 25788 13916 25844
rect 13972 25788 17052 25844
rect 17108 25788 17118 25844
rect 17276 25788 19628 25844
rect 19684 25788 19694 25844
rect 20412 25788 22764 25844
rect 22820 25788 23548 25844
rect 23604 25788 23614 25844
rect 27234 25788 27244 25844
rect 27300 25788 27310 25844
rect 27692 25788 31108 25844
rect 42130 25788 42140 25844
rect 42196 25788 47404 25844
rect 47460 25788 47628 25844
rect 47684 25788 48188 25844
rect 48244 25788 48254 25844
rect 20412 25732 20468 25788
rect 27692 25732 27748 25788
rect 10770 25676 10780 25732
rect 10836 25676 12796 25732
rect 12852 25676 14700 25732
rect 14756 25676 18284 25732
rect 18340 25676 18350 25732
rect 19506 25676 19516 25732
rect 19572 25676 20468 25732
rect 20524 25676 21308 25732
rect 21364 25676 21532 25732
rect 21588 25676 21598 25732
rect 27682 25676 27692 25732
rect 27748 25676 27758 25732
rect 29586 25676 29596 25732
rect 29652 25676 30604 25732
rect 30660 25676 30670 25732
rect 20524 25620 20580 25676
rect 31052 25620 31108 25788
rect 34514 25676 34524 25732
rect 34580 25676 35980 25732
rect 36036 25676 40012 25732
rect 40068 25676 40078 25732
rect 45826 25676 45836 25732
rect 45892 25676 46508 25732
rect 46564 25676 46574 25732
rect 2146 25564 2156 25620
rect 2212 25564 4620 25620
rect 4676 25564 4686 25620
rect 12562 25564 12572 25620
rect 12628 25564 13692 25620
rect 13748 25564 13758 25620
rect 14242 25564 14252 25620
rect 14308 25564 20580 25620
rect 20738 25564 20748 25620
rect 20804 25564 21868 25620
rect 21924 25564 21934 25620
rect 27570 25564 27580 25620
rect 27636 25564 30044 25620
rect 30100 25564 30110 25620
rect 31052 25564 39228 25620
rect 39284 25564 39294 25620
rect 44930 25564 44940 25620
rect 44996 25564 47516 25620
rect 47572 25564 47582 25620
rect 6738 25452 6748 25508
rect 6804 25452 8540 25508
rect 8596 25452 8606 25508
rect 17042 25452 17052 25508
rect 17108 25452 19516 25508
rect 19572 25452 19582 25508
rect 19730 25452 19740 25508
rect 19796 25452 26012 25508
rect 26068 25452 26078 25508
rect 26226 25452 26236 25508
rect 26292 25452 26684 25508
rect 26740 25452 29484 25508
rect 29540 25452 29550 25508
rect 34962 25452 34972 25508
rect 35028 25452 36092 25508
rect 36148 25452 36158 25508
rect 37538 25452 37548 25508
rect 37604 25452 42140 25508
rect 42196 25452 42206 25508
rect 45042 25452 45052 25508
rect 45108 25452 47404 25508
rect 47460 25452 47470 25508
rect 5954 25340 5964 25396
rect 6020 25340 9548 25396
rect 9604 25340 10220 25396
rect 10276 25340 10286 25396
rect 11228 25340 13692 25396
rect 13748 25340 19068 25396
rect 19124 25340 20860 25396
rect 20916 25340 20926 25396
rect 26562 25340 26572 25396
rect 26628 25340 27356 25396
rect 27412 25340 27422 25396
rect 27570 25340 27580 25396
rect 27636 25340 28588 25396
rect 28644 25340 28654 25396
rect 31266 25340 31276 25396
rect 31332 25340 31948 25396
rect 32004 25340 32014 25396
rect 32162 25340 32172 25396
rect 32228 25340 33068 25396
rect 33124 25340 33134 25396
rect 34850 25340 34860 25396
rect 34916 25340 35420 25396
rect 35476 25340 35486 25396
rect 45266 25340 45276 25396
rect 45332 25340 47180 25396
rect 47236 25340 47246 25396
rect 5058 25228 5068 25284
rect 5124 25228 5516 25284
rect 5572 25228 7420 25284
rect 7476 25228 7486 25284
rect 1474 25116 1484 25172
rect 1540 25116 2156 25172
rect 2212 25116 2222 25172
rect 11228 25060 11284 25340
rect 14354 25228 14364 25284
rect 14420 25228 15036 25284
rect 15092 25228 18284 25284
rect 18340 25228 18350 25284
rect 18498 25228 18508 25284
rect 18564 25228 19404 25284
rect 19460 25228 19470 25284
rect 19618 25228 19628 25284
rect 19684 25228 19964 25284
rect 20020 25228 20030 25284
rect 20626 25228 20636 25284
rect 20692 25228 21084 25284
rect 21140 25228 21756 25284
rect 21812 25228 21822 25284
rect 22754 25228 22764 25284
rect 22820 25228 23436 25284
rect 23492 25228 23502 25284
rect 23762 25228 23772 25284
rect 23828 25228 26908 25284
rect 26964 25228 28252 25284
rect 28308 25228 28318 25284
rect 29138 25228 29148 25284
rect 29204 25228 31052 25284
rect 31108 25228 31118 25284
rect 34290 25228 34300 25284
rect 34356 25228 35196 25284
rect 35252 25228 35262 25284
rect 36530 25228 36540 25284
rect 36596 25228 37436 25284
rect 37492 25228 37502 25284
rect 39778 25228 39788 25284
rect 39844 25228 40236 25284
rect 40292 25228 40908 25284
rect 40964 25228 41580 25284
rect 41636 25228 41646 25284
rect 46050 25228 46060 25284
rect 46116 25228 47292 25284
rect 47348 25228 47358 25284
rect 15474 25116 15484 25172
rect 15540 25116 16268 25172
rect 16324 25116 16828 25172
rect 16884 25116 17836 25172
rect 17892 25116 17902 25172
rect 20290 25116 20300 25172
rect 20356 25116 20748 25172
rect 20804 25116 20814 25172
rect 25218 25116 25228 25172
rect 25284 25116 27356 25172
rect 27412 25116 27422 25172
rect 33506 25116 33516 25172
rect 33572 25116 34972 25172
rect 35028 25116 35038 25172
rect 37090 25116 37100 25172
rect 37156 25116 37772 25172
rect 37828 25116 37838 25172
rect 41234 25116 41244 25172
rect 41300 25116 41916 25172
rect 41972 25116 41982 25172
rect 46722 25116 46732 25172
rect 46788 25116 47628 25172
rect 47684 25116 47694 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 5394 25004 5404 25060
rect 5460 25004 11284 25060
rect 18274 25004 18284 25060
rect 18340 25004 18620 25060
rect 18676 25004 18686 25060
rect 30482 25004 30492 25060
rect 30548 25004 31276 25060
rect 31332 25004 31342 25060
rect 0 24948 800 24976
rect 0 24892 1596 24948
rect 1652 24892 1662 24948
rect 5058 24892 5068 24948
rect 5124 24892 5292 24948
rect 5348 24892 5358 24948
rect 5618 24892 5628 24948
rect 5684 24892 6412 24948
rect 6468 24892 9548 24948
rect 9604 24892 9614 24948
rect 11778 24892 11788 24948
rect 11844 24892 13020 24948
rect 13076 24892 13086 24948
rect 16818 24892 16828 24948
rect 16884 24892 22204 24948
rect 22260 24892 22270 24948
rect 25890 24892 25900 24948
rect 25956 24892 39116 24948
rect 39172 24892 39182 24948
rect 0 24864 800 24892
rect 2930 24780 2940 24836
rect 2996 24780 3836 24836
rect 3892 24780 6188 24836
rect 6244 24780 6972 24836
rect 7028 24780 7038 24836
rect 13794 24780 13804 24836
rect 13860 24780 14812 24836
rect 14868 24780 14878 24836
rect 17910 24780 17948 24836
rect 18004 24780 18014 24836
rect 18246 24780 18284 24836
rect 18340 24780 18350 24836
rect 18806 24780 18844 24836
rect 18900 24780 18910 24836
rect 33058 24780 33068 24836
rect 33124 24780 34748 24836
rect 34804 24780 34814 24836
rect 40338 24780 40348 24836
rect 40404 24780 41244 24836
rect 41300 24780 41310 24836
rect 2706 24668 2716 24724
rect 2772 24668 3388 24724
rect 3444 24668 3724 24724
rect 3780 24668 8204 24724
rect 8260 24668 8270 24724
rect 12226 24668 12236 24724
rect 12292 24668 14028 24724
rect 14084 24668 14094 24724
rect 14690 24668 14700 24724
rect 14756 24668 17500 24724
rect 17556 24668 20076 24724
rect 20132 24668 20142 24724
rect 22754 24668 22764 24724
rect 22820 24668 23548 24724
rect 23604 24668 23614 24724
rect 25190 24668 25228 24724
rect 25284 24668 25294 24724
rect 30258 24668 30268 24724
rect 30324 24668 30940 24724
rect 30996 24668 31006 24724
rect 32274 24668 32284 24724
rect 32340 24668 35084 24724
rect 35140 24668 35150 24724
rect 38770 24668 38780 24724
rect 38836 24668 41356 24724
rect 41412 24668 42252 24724
rect 42308 24668 42318 24724
rect 45154 24668 45164 24724
rect 45220 24668 45948 24724
rect 46004 24668 46014 24724
rect 47954 24668 47964 24724
rect 48020 24668 48412 24724
rect 48468 24668 48478 24724
rect 14130 24556 14140 24612
rect 14196 24556 14924 24612
rect 14980 24556 14990 24612
rect 18162 24556 18172 24612
rect 18228 24556 28588 24612
rect 28644 24556 28654 24612
rect 33842 24556 33852 24612
rect 33908 24556 34748 24612
rect 34804 24556 34814 24612
rect 35858 24556 35868 24612
rect 35924 24556 36988 24612
rect 37044 24556 37054 24612
rect 13570 24444 13580 24500
rect 13636 24444 18956 24500
rect 19012 24444 19022 24500
rect 43474 24444 43484 24500
rect 43540 24444 45612 24500
rect 45668 24444 45678 24500
rect 14578 24332 14588 24388
rect 14644 24332 19628 24388
rect 19684 24332 19694 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 10546 24220 10556 24276
rect 10612 24220 13804 24276
rect 13860 24220 22540 24276
rect 22596 24220 22606 24276
rect 30930 24220 30940 24276
rect 30996 24220 32172 24276
rect 32228 24220 32238 24276
rect 2818 24108 2828 24164
rect 2884 24108 3164 24164
rect 3220 24108 4284 24164
rect 4340 24108 4350 24164
rect 10882 24108 10892 24164
rect 10948 24108 30828 24164
rect 30884 24108 31388 24164
rect 31444 24108 31724 24164
rect 31780 24108 32732 24164
rect 32788 24108 32798 24164
rect 3042 23996 3052 24052
rect 3108 23996 5068 24052
rect 5124 23996 5134 24052
rect 8306 23996 8316 24052
rect 8372 23996 12012 24052
rect 12068 23996 12078 24052
rect 14130 23996 14140 24052
rect 14196 23996 17164 24052
rect 17220 23996 17230 24052
rect 19058 23996 19068 24052
rect 19124 23996 32508 24052
rect 32564 23996 32574 24052
rect 45042 23996 45052 24052
rect 45108 23996 47964 24052
rect 48020 23996 48030 24052
rect 2594 23884 2604 23940
rect 2660 23884 4508 23940
rect 4564 23884 4574 23940
rect 6066 23884 6076 23940
rect 6132 23884 6860 23940
rect 6916 23884 9660 23940
rect 9716 23884 9726 23940
rect 11890 23884 11900 23940
rect 11956 23884 13468 23940
rect 13524 23884 13534 23940
rect 17490 23884 17500 23940
rect 17556 23884 19740 23940
rect 19796 23884 19806 23940
rect 20514 23884 20524 23940
rect 20580 23884 20860 23940
rect 20916 23884 21420 23940
rect 21476 23884 21486 23940
rect 23090 23884 23100 23940
rect 23156 23884 27916 23940
rect 27972 23884 27982 23940
rect 29586 23884 29596 23940
rect 29652 23884 29932 23940
rect 29988 23884 29998 23940
rect 4274 23772 4284 23828
rect 4340 23772 5516 23828
rect 5572 23772 5582 23828
rect 12114 23772 12124 23828
rect 12180 23772 15596 23828
rect 15652 23772 15662 23828
rect 15922 23772 15932 23828
rect 15988 23772 16380 23828
rect 16436 23772 17612 23828
rect 17668 23772 18620 23828
rect 18676 23772 20636 23828
rect 20692 23772 20702 23828
rect 23426 23772 23436 23828
rect 23492 23772 30156 23828
rect 30212 23772 30222 23828
rect 41234 23772 41244 23828
rect 41300 23772 43148 23828
rect 43204 23772 44380 23828
rect 44436 23772 44446 23828
rect 3154 23660 3164 23716
rect 3220 23660 4844 23716
rect 4900 23660 4910 23716
rect 13010 23660 13020 23716
rect 13076 23660 13468 23716
rect 13524 23660 13534 23716
rect 15092 23660 20188 23716
rect 20244 23660 20254 23716
rect 35746 23660 35756 23716
rect 35812 23660 39676 23716
rect 39732 23660 40124 23716
rect 40180 23660 41356 23716
rect 41412 23660 42476 23716
rect 42532 23660 42542 23716
rect 42802 23660 42812 23716
rect 42868 23660 44828 23716
rect 44884 23660 44894 23716
rect 15092 23492 15148 23660
rect 15698 23548 15708 23604
rect 15764 23548 17612 23604
rect 17668 23548 17678 23604
rect 25330 23548 25340 23604
rect 25396 23548 30268 23604
rect 30324 23548 30334 23604
rect 34514 23548 34524 23604
rect 34580 23548 35868 23604
rect 35924 23548 35934 23604
rect 40002 23548 40012 23604
rect 40068 23548 41132 23604
rect 41188 23548 41198 23604
rect 41570 23548 41580 23604
rect 41636 23548 41916 23604
rect 41972 23548 42700 23604
rect 42756 23548 42766 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 2482 23436 2492 23492
rect 2548 23436 3948 23492
rect 4004 23436 4014 23492
rect 6402 23436 6412 23492
rect 6468 23436 10780 23492
rect 10836 23436 10846 23492
rect 11666 23436 11676 23492
rect 11732 23436 12124 23492
rect 12180 23436 12190 23492
rect 14242 23436 14252 23492
rect 14308 23436 15148 23492
rect 16594 23436 16604 23492
rect 16660 23436 19180 23492
rect 19236 23436 19246 23492
rect 20972 23436 27076 23492
rect 2370 23324 2380 23380
rect 2436 23324 3612 23380
rect 3668 23324 4732 23380
rect 4788 23324 5628 23380
rect 5684 23324 5694 23380
rect 10210 23324 10220 23380
rect 10276 23324 15148 23380
rect 20066 23324 20076 23380
rect 20132 23324 20412 23380
rect 20468 23324 20478 23380
rect 15092 23268 15148 23324
rect 20972 23268 21028 23436
rect 27020 23380 27076 23436
rect 28476 23436 31388 23492
rect 31444 23436 38556 23492
rect 38612 23436 38622 23492
rect 28476 23380 28532 23436
rect 23174 23324 23212 23380
rect 23268 23324 23278 23380
rect 23650 23324 23660 23380
rect 23716 23324 24108 23380
rect 24164 23324 24556 23380
rect 24612 23324 26908 23380
rect 27020 23324 28532 23380
rect 30818 23324 30828 23380
rect 30884 23324 31500 23380
rect 31556 23324 32060 23380
rect 32116 23324 32126 23380
rect 26852 23268 26908 23324
rect 9650 23212 9660 23268
rect 9716 23212 10108 23268
rect 10164 23212 10174 23268
rect 11554 23212 11564 23268
rect 11620 23212 12236 23268
rect 12292 23212 12302 23268
rect 15092 23212 21028 23268
rect 22866 23212 22876 23268
rect 22932 23212 23772 23268
rect 23828 23212 24332 23268
rect 24388 23212 24398 23268
rect 26002 23212 26012 23268
rect 26068 23212 26572 23268
rect 26628 23212 26638 23268
rect 26852 23212 27916 23268
rect 27972 23212 27982 23268
rect 28130 23212 28140 23268
rect 28196 23212 31724 23268
rect 31780 23212 31790 23268
rect 44930 23212 44940 23268
rect 44996 23212 46396 23268
rect 46452 23212 46462 23268
rect 47170 23212 47180 23268
rect 47236 23212 47516 23268
rect 47572 23212 47852 23268
rect 47908 23212 47918 23268
rect 6178 23100 6188 23156
rect 6244 23100 15316 23156
rect 11666 22988 11676 23044
rect 11732 22988 14476 23044
rect 14532 22988 14542 23044
rect 15260 22932 15316 23100
rect 23492 23100 32508 23156
rect 32564 23100 32574 23156
rect 38210 23100 38220 23156
rect 38276 23100 38892 23156
rect 38948 23100 38958 23156
rect 44146 23100 44156 23156
rect 44212 23100 45276 23156
rect 45332 23100 46732 23156
rect 46788 23100 46798 23156
rect 15474 22988 15484 23044
rect 15540 22988 19068 23044
rect 19124 22988 19134 23044
rect 23492 22932 23548 23100
rect 23762 22988 23772 23044
rect 23828 22988 30268 23044
rect 30324 22988 30828 23044
rect 30884 22988 30894 23044
rect 31154 22988 31164 23044
rect 31220 22988 33964 23044
rect 34020 22988 34030 23044
rect 38434 22988 38444 23044
rect 38500 22988 39004 23044
rect 39060 22988 39070 23044
rect 41682 22988 41692 23044
rect 41748 22988 44268 23044
rect 44324 22988 44334 23044
rect 47394 22988 47404 23044
rect 47460 22988 48076 23044
rect 48132 22988 48142 23044
rect 8194 22876 8204 22932
rect 8260 22876 12012 22932
rect 12068 22876 12078 22932
rect 15260 22876 16044 22932
rect 16100 22876 18844 22932
rect 18900 22876 19068 22932
rect 19124 22876 19292 22932
rect 19348 22876 23548 22932
rect 24546 22876 24556 22932
rect 24612 22876 27132 22932
rect 27188 22876 28028 22932
rect 28084 22876 28094 22932
rect 31164 22820 31220 22988
rect 39218 22876 39228 22932
rect 39284 22876 40572 22932
rect 40628 22876 40638 22932
rect 15362 22764 15372 22820
rect 15428 22764 19068 22820
rect 19124 22764 19134 22820
rect 19394 22764 19404 22820
rect 19460 22764 20076 22820
rect 20132 22764 20142 22820
rect 27906 22764 27916 22820
rect 27972 22764 31220 22820
rect 43138 22764 43148 22820
rect 43204 22764 43820 22820
rect 43876 22764 45948 22820
rect 46004 22764 46014 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 10882 22652 10892 22708
rect 10948 22652 12796 22708
rect 12852 22652 12862 22708
rect 16380 22652 20412 22708
rect 20468 22652 20478 22708
rect 27122 22652 27132 22708
rect 27188 22652 28252 22708
rect 28308 22652 28318 22708
rect 29922 22652 29932 22708
rect 29988 22652 32956 22708
rect 33012 22652 33022 22708
rect 16380 22596 16436 22652
rect 12898 22540 12908 22596
rect 12964 22540 15148 22596
rect 15204 22540 16436 22596
rect 16594 22540 16604 22596
rect 16660 22540 16670 22596
rect 19170 22540 19180 22596
rect 19236 22540 19516 22596
rect 19572 22540 19582 22596
rect 22978 22540 22988 22596
rect 23044 22540 31724 22596
rect 31780 22540 31790 22596
rect 43362 22540 43372 22596
rect 43428 22540 44156 22596
rect 44212 22540 45724 22596
rect 45780 22540 45790 22596
rect 3938 22428 3948 22484
rect 4004 22428 6972 22484
rect 7028 22428 7038 22484
rect 16604 22372 16660 22540
rect 49200 22484 50000 22512
rect 18722 22428 18732 22484
rect 18788 22428 19628 22484
rect 19684 22428 19694 22484
rect 25302 22428 25340 22484
rect 25396 22428 25406 22484
rect 40786 22428 40796 22484
rect 40852 22428 41132 22484
rect 41188 22428 42252 22484
rect 42308 22428 42318 22484
rect 48076 22428 50000 22484
rect 11106 22316 11116 22372
rect 11172 22316 13692 22372
rect 13748 22316 16660 22372
rect 18946 22316 18956 22372
rect 19012 22316 20076 22372
rect 20132 22316 20142 22372
rect 25106 22316 25116 22372
rect 25172 22316 25452 22372
rect 25508 22316 28140 22372
rect 28196 22316 28206 22372
rect 46610 22316 46620 22372
rect 46676 22316 47180 22372
rect 47236 22316 47246 22372
rect 48076 22260 48132 22428
rect 49200 22400 50000 22428
rect 15596 22204 22092 22260
rect 22148 22204 22158 22260
rect 25106 22204 25116 22260
rect 25172 22204 25228 22260
rect 25284 22204 25294 22260
rect 37398 22204 37436 22260
rect 37492 22204 37502 22260
rect 38994 22204 39004 22260
rect 39060 22204 40460 22260
rect 40516 22204 40526 22260
rect 48066 22204 48076 22260
rect 48132 22204 48142 22260
rect 15596 22148 15652 22204
rect 1362 22092 1372 22148
rect 1428 22092 3836 22148
rect 3892 22092 3902 22148
rect 12338 22092 12348 22148
rect 12404 22092 15204 22148
rect 15362 22092 15372 22148
rect 15428 22092 15596 22148
rect 15652 22092 15662 22148
rect 16828 22092 20188 22148
rect 20244 22092 20254 22148
rect 23762 22092 23772 22148
rect 23828 22092 24444 22148
rect 24500 22092 25564 22148
rect 25620 22092 25630 22148
rect 27570 22092 27580 22148
rect 27636 22092 28700 22148
rect 28756 22092 28766 22148
rect 31490 22092 31500 22148
rect 31556 22092 35756 22148
rect 35812 22092 36988 22148
rect 37044 22092 37054 22148
rect 42242 22092 42252 22148
rect 42308 22092 44044 22148
rect 44100 22092 44110 22148
rect 12348 22036 12404 22092
rect 15148 22036 15204 22092
rect 16828 22036 16884 22092
rect 1474 21980 1484 22036
rect 1540 21980 12404 22036
rect 12898 21980 12908 22036
rect 12964 21980 14140 22036
rect 14196 21980 14206 22036
rect 15148 21980 16884 22036
rect 32946 21980 32956 22036
rect 33012 21980 33628 22036
rect 33684 21980 36092 22036
rect 36148 21980 36158 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 10210 21868 10220 21924
rect 10276 21868 10444 21924
rect 10500 21868 10510 21924
rect 17378 21868 17388 21924
rect 17444 21868 19292 21924
rect 19348 21868 19358 21924
rect 22754 21868 22764 21924
rect 22820 21868 24332 21924
rect 24388 21868 24892 21924
rect 24948 21868 24958 21924
rect 29698 21868 29708 21924
rect 29764 21868 31276 21924
rect 31332 21868 32284 21924
rect 32340 21868 32350 21924
rect 40114 21868 40124 21924
rect 40180 21868 41020 21924
rect 41076 21868 41916 21924
rect 41972 21868 41982 21924
rect 7410 21756 7420 21812
rect 7476 21756 10780 21812
rect 10836 21756 10846 21812
rect 11666 21756 11676 21812
rect 11732 21756 14924 21812
rect 14980 21756 14990 21812
rect 16706 21756 16716 21812
rect 16772 21756 17500 21812
rect 17556 21756 17566 21812
rect 17938 21756 17948 21812
rect 18004 21756 18732 21812
rect 18788 21756 18798 21812
rect 21410 21756 21420 21812
rect 21476 21756 21868 21812
rect 21924 21756 21934 21812
rect 25218 21756 25228 21812
rect 25284 21756 25340 21812
rect 25396 21756 25406 21812
rect 36418 21756 36428 21812
rect 36484 21756 37212 21812
rect 37268 21756 37884 21812
rect 37940 21756 38444 21812
rect 38500 21756 38510 21812
rect 2034 21644 2044 21700
rect 2100 21644 4396 21700
rect 4452 21644 4732 21700
rect 4788 21644 4798 21700
rect 5170 21644 5180 21700
rect 5236 21644 5852 21700
rect 5908 21644 8204 21700
rect 8260 21644 8270 21700
rect 11106 21644 11116 21700
rect 11172 21644 13244 21700
rect 13300 21644 13310 21700
rect 16594 21644 16604 21700
rect 16660 21644 19404 21700
rect 19460 21644 19470 21700
rect 20178 21644 20188 21700
rect 20244 21644 20300 21700
rect 20356 21644 20524 21700
rect 20580 21644 20590 21700
rect 21186 21644 21196 21700
rect 21252 21644 23660 21700
rect 23716 21644 23726 21700
rect 27906 21644 27916 21700
rect 27972 21644 29036 21700
rect 29092 21644 29102 21700
rect 29250 21644 29260 21700
rect 29316 21644 30492 21700
rect 30548 21644 30558 21700
rect 36306 21644 36316 21700
rect 36372 21644 37324 21700
rect 37380 21644 37390 21700
rect 37650 21644 37660 21700
rect 37716 21644 38108 21700
rect 38164 21644 38332 21700
rect 38388 21644 38398 21700
rect 46386 21644 46396 21700
rect 46452 21644 47180 21700
rect 47236 21644 47246 21700
rect 47842 21644 47852 21700
rect 47908 21644 47918 21700
rect 37660 21588 37716 21644
rect 47852 21588 47908 21644
rect 4610 21532 4620 21588
rect 4676 21532 5068 21588
rect 5124 21532 5292 21588
rect 5348 21532 5358 21588
rect 10658 21532 10668 21588
rect 10724 21532 12012 21588
rect 12068 21532 12078 21588
rect 12226 21532 12236 21588
rect 12292 21532 16492 21588
rect 16548 21532 16558 21588
rect 16706 21532 16716 21588
rect 16772 21532 19740 21588
rect 19796 21532 19806 21588
rect 20066 21532 20076 21588
rect 20132 21532 22540 21588
rect 22596 21532 22606 21588
rect 23538 21532 23548 21588
rect 23604 21532 26012 21588
rect 26068 21532 27692 21588
rect 27748 21532 27758 21588
rect 30594 21532 30604 21588
rect 30660 21532 31052 21588
rect 31108 21532 32508 21588
rect 32564 21532 32574 21588
rect 36194 21532 36204 21588
rect 36260 21532 37716 21588
rect 45378 21532 45388 21588
rect 45444 21532 47908 21588
rect 1922 21420 1932 21476
rect 1988 21420 2268 21476
rect 2324 21420 2334 21476
rect 11106 21420 11116 21476
rect 11172 21420 11182 21476
rect 15362 21420 15372 21476
rect 15428 21420 17500 21476
rect 17556 21420 17566 21476
rect 22754 21420 22764 21476
rect 22820 21420 23884 21476
rect 23940 21420 33068 21476
rect 33124 21420 33292 21476
rect 33348 21420 34020 21476
rect 34850 21420 34860 21476
rect 34916 21420 37772 21476
rect 37828 21420 37838 21476
rect 39778 21420 39788 21476
rect 39844 21420 40908 21476
rect 40964 21420 40974 21476
rect 44034 21420 44044 21476
rect 44100 21420 47068 21476
rect 47124 21420 47134 21476
rect 1138 21308 1148 21364
rect 1204 21308 5740 21364
rect 5796 21308 5806 21364
rect 11116 21252 11172 21420
rect 33964 21364 34020 21420
rect 16482 21308 16492 21364
rect 16548 21308 17836 21364
rect 17892 21308 17902 21364
rect 23314 21308 23324 21364
rect 23380 21308 24556 21364
rect 24612 21308 26684 21364
rect 26740 21308 26750 21364
rect 33954 21308 33964 21364
rect 34020 21308 34030 21364
rect 41794 21308 41804 21364
rect 41860 21308 42812 21364
rect 42868 21308 43932 21364
rect 43988 21308 43998 21364
rect 10770 21196 10780 21252
rect 10836 21196 11172 21252
rect 13010 21196 13020 21252
rect 13076 21196 16940 21252
rect 16996 21196 17948 21252
rect 18004 21196 18014 21252
rect 18172 21196 18956 21252
rect 19012 21196 19022 21252
rect 21410 21196 21420 21252
rect 21476 21196 22204 21252
rect 22260 21196 22270 21252
rect 45266 21196 45276 21252
rect 45332 21196 45342 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 14914 21084 14924 21140
rect 14980 21084 15764 21140
rect 3266 20972 3276 21028
rect 3332 20972 4060 21028
rect 4116 20972 6748 21028
rect 6804 20972 6814 21028
rect 7746 20972 7756 21028
rect 7812 20972 8540 21028
rect 8596 20972 8606 21028
rect 13234 20972 13244 21028
rect 13300 20972 15260 21028
rect 15316 20972 15326 21028
rect 15708 20916 15764 21084
rect 18172 21028 18228 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 19618 21084 19628 21140
rect 19684 21084 22316 21140
rect 22372 21084 22382 21140
rect 25442 21084 25452 21140
rect 25508 21084 34076 21140
rect 34132 21084 34524 21140
rect 34580 21084 34590 21140
rect 45276 21028 45332 21196
rect 15922 20972 15932 21028
rect 15988 20972 18228 21028
rect 18284 20972 20412 21028
rect 20468 20972 20478 21028
rect 29922 20972 29932 21028
rect 29988 20972 45332 21028
rect 18284 20916 18340 20972
rect 2706 20860 2716 20916
rect 2772 20860 3388 20916
rect 5730 20860 5740 20916
rect 5796 20860 9772 20916
rect 9828 20860 9838 20916
rect 15708 20860 15820 20916
rect 15876 20860 18340 20916
rect 18498 20860 18508 20916
rect 18564 20860 19068 20916
rect 19124 20860 19134 20916
rect 19282 20860 19292 20916
rect 19348 20860 19386 20916
rect 21746 20860 21756 20916
rect 21812 20860 25564 20916
rect 25620 20860 25630 20916
rect 28466 20860 28476 20916
rect 28532 20860 29148 20916
rect 29204 20860 29820 20916
rect 29876 20860 29886 20916
rect 33170 20860 33180 20916
rect 33236 20860 39228 20916
rect 39284 20860 39294 20916
rect 44370 20860 44380 20916
rect 44436 20860 48076 20916
rect 48132 20860 48142 20916
rect 3332 20804 3388 20860
rect 3332 20748 6300 20804
rect 6356 20748 6366 20804
rect 12562 20748 12572 20804
rect 12628 20748 12908 20804
rect 12964 20748 12974 20804
rect 18274 20748 18284 20804
rect 18340 20748 18956 20804
rect 19012 20748 19022 20804
rect 21522 20748 21532 20804
rect 21588 20748 23212 20804
rect 23268 20748 23278 20804
rect 23762 20748 23772 20804
rect 23828 20748 25340 20804
rect 25396 20748 25406 20804
rect 28242 20748 28252 20804
rect 28308 20748 29372 20804
rect 29428 20748 29438 20804
rect 30706 20748 30716 20804
rect 30772 20748 32284 20804
rect 32340 20748 32350 20804
rect 36306 20748 36316 20804
rect 36372 20748 36988 20804
rect 37044 20748 37054 20804
rect 6066 20636 6076 20692
rect 6132 20636 7756 20692
rect 7812 20636 7822 20692
rect 11666 20636 11676 20692
rect 11732 20636 15708 20692
rect 15764 20636 15774 20692
rect 16930 20636 16940 20692
rect 16996 20636 19068 20692
rect 19124 20636 19134 20692
rect 19282 20636 19292 20692
rect 19348 20636 19404 20692
rect 19460 20636 22092 20692
rect 22148 20636 22158 20692
rect 24210 20636 24220 20692
rect 24276 20636 28364 20692
rect 28420 20636 28430 20692
rect 30716 20580 30772 20748
rect 34178 20636 34188 20692
rect 34244 20636 41692 20692
rect 41748 20636 41758 20692
rect 6514 20524 6524 20580
rect 6580 20524 8092 20580
rect 8148 20524 10220 20580
rect 10276 20524 10286 20580
rect 10546 20524 10556 20580
rect 10612 20524 13132 20580
rect 13188 20524 14028 20580
rect 14084 20524 14094 20580
rect 18610 20524 18620 20580
rect 18676 20524 20748 20580
rect 20804 20524 20814 20580
rect 24994 20524 25004 20580
rect 25060 20524 27020 20580
rect 27076 20524 27580 20580
rect 27636 20524 27646 20580
rect 27906 20524 27916 20580
rect 27972 20524 30772 20580
rect 31826 20524 31836 20580
rect 31892 20524 33964 20580
rect 34020 20524 34030 20580
rect 35410 20524 35420 20580
rect 35476 20524 37100 20580
rect 37156 20524 37884 20580
rect 37940 20524 37950 20580
rect 7970 20412 7980 20468
rect 8036 20412 9884 20468
rect 9940 20412 11900 20468
rect 11956 20412 11966 20468
rect 14802 20412 14812 20468
rect 14868 20412 15932 20468
rect 15988 20412 15998 20468
rect 17490 20412 17500 20468
rect 17556 20412 19404 20468
rect 19460 20412 19470 20468
rect 26114 20412 26124 20468
rect 26180 20412 30604 20468
rect 30660 20412 31164 20468
rect 31220 20412 34412 20468
rect 34468 20412 34478 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 17490 20300 17500 20356
rect 17556 20300 17724 20356
rect 17780 20300 17790 20356
rect 18358 20300 18396 20356
rect 18452 20300 18462 20356
rect 25554 20300 25564 20356
rect 25620 20300 27692 20356
rect 27748 20300 29036 20356
rect 29092 20300 29102 20356
rect 30930 20300 30940 20356
rect 30996 20300 31836 20356
rect 31892 20300 34636 20356
rect 34692 20300 34702 20356
rect 38434 20300 38444 20356
rect 38500 20300 38668 20356
rect 5282 20188 5292 20244
rect 5348 20188 7420 20244
rect 7476 20188 7486 20244
rect 9986 20188 9996 20244
rect 10052 20188 15484 20244
rect 15540 20188 15550 20244
rect 15698 20188 15708 20244
rect 15764 20188 20188 20244
rect 20244 20188 20254 20244
rect 25078 20188 25116 20244
rect 25172 20188 25182 20244
rect 25442 20188 25452 20244
rect 25508 20188 32116 20244
rect 11554 20076 11564 20132
rect 11620 20076 14252 20132
rect 14308 20076 14318 20132
rect 19142 20076 19180 20132
rect 19236 20076 19246 20132
rect 20738 20076 20748 20132
rect 20804 20076 21644 20132
rect 21700 20076 21710 20132
rect 25330 20076 25340 20132
rect 25396 20076 27916 20132
rect 27972 20076 27982 20132
rect 9874 19964 9884 20020
rect 9940 19964 11228 20020
rect 11284 19964 13468 20020
rect 13524 19964 13534 20020
rect 17602 19964 17612 20020
rect 17668 19964 19292 20020
rect 19348 19964 19358 20020
rect 20178 19964 20188 20020
rect 20244 19964 20636 20020
rect 20692 19964 20702 20020
rect 26786 19964 26796 20020
rect 26852 19964 27132 20020
rect 27188 19964 27468 20020
rect 27524 19964 27534 20020
rect 1026 19852 1036 19908
rect 1092 19852 2156 19908
rect 2212 19852 2222 19908
rect 3826 19852 3836 19908
rect 3892 19852 8092 19908
rect 8148 19852 8158 19908
rect 18162 19852 18172 19908
rect 18228 19852 19068 19908
rect 19124 19852 19292 19908
rect 19348 19852 22204 19908
rect 22260 19852 22270 19908
rect 32060 19796 32116 20188
rect 38612 20132 38668 20300
rect 45042 20188 45052 20244
rect 45108 20188 46396 20244
rect 46452 20188 46462 20244
rect 34066 20076 34076 20132
rect 34132 20076 35308 20132
rect 35364 20076 36092 20132
rect 36148 20076 36158 20132
rect 38612 20076 38780 20132
rect 38836 20076 38846 20132
rect 38546 19964 38556 20020
rect 38612 19964 39004 20020
rect 39060 19964 39070 20020
rect 43922 19964 43932 20020
rect 43988 19964 45052 20020
rect 45108 19964 45118 20020
rect 45826 19964 45836 20020
rect 45892 19964 46844 20020
rect 46900 19964 47740 20020
rect 47796 19964 47806 20020
rect 32498 19852 32508 19908
rect 32564 19852 40236 19908
rect 40292 19852 40302 19908
rect 44594 19852 44604 19908
rect 44660 19852 45276 19908
rect 45332 19852 45342 19908
rect 3042 19740 3052 19796
rect 3108 19740 5292 19796
rect 5348 19740 5358 19796
rect 16818 19740 16828 19796
rect 16884 19740 21532 19796
rect 21588 19740 21598 19796
rect 23538 19740 23548 19796
rect 23604 19740 23884 19796
rect 23940 19740 23950 19796
rect 24322 19740 24332 19796
rect 24388 19740 25340 19796
rect 25396 19740 25406 19796
rect 32050 19740 32060 19796
rect 32116 19740 32126 19796
rect 32508 19684 32564 19852
rect 32834 19740 32844 19796
rect 32900 19740 39676 19796
rect 39732 19740 39742 19796
rect 47058 19740 47068 19796
rect 47124 19740 47852 19796
rect 47908 19740 47918 19796
rect 15586 19628 15596 19684
rect 15652 19628 18620 19684
rect 18676 19628 18686 19684
rect 19254 19628 19292 19684
rect 19348 19628 20860 19684
rect 20916 19628 20926 19684
rect 21410 19628 21420 19684
rect 21476 19628 22540 19684
rect 22596 19628 23100 19684
rect 23156 19628 24444 19684
rect 24500 19628 24510 19684
rect 30818 19628 30828 19684
rect 30884 19628 32564 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 32844 19572 32900 19740
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 4956 19516 7868 19572
rect 7924 19516 7934 19572
rect 17350 19516 17388 19572
rect 17444 19516 18172 19572
rect 18228 19516 19852 19572
rect 19908 19516 23660 19572
rect 23716 19516 23726 19572
rect 23874 19516 23884 19572
rect 23940 19516 29708 19572
rect 29764 19516 29774 19572
rect 31042 19516 31052 19572
rect 31108 19516 32900 19572
rect 4956 19460 5012 19516
rect 29708 19460 29764 19516
rect 1922 19404 1932 19460
rect 1988 19404 3948 19460
rect 4004 19404 5012 19460
rect 6178 19404 6188 19460
rect 6244 19404 7644 19460
rect 7700 19404 17500 19460
rect 17556 19404 17566 19460
rect 17714 19404 17724 19460
rect 17780 19404 18396 19460
rect 18452 19404 18462 19460
rect 19730 19404 19740 19460
rect 19796 19404 20804 19460
rect 23202 19404 23212 19460
rect 23268 19404 24780 19460
rect 24836 19404 26684 19460
rect 26740 19404 26908 19460
rect 29708 19404 31724 19460
rect 31780 19404 34636 19460
rect 34692 19404 35420 19460
rect 35476 19404 36540 19460
rect 36596 19404 36606 19460
rect 20748 19348 20804 19404
rect 1698 19292 1708 19348
rect 1764 19292 2940 19348
rect 2996 19292 3006 19348
rect 4050 19292 4060 19348
rect 4116 19292 5628 19348
rect 5684 19292 5694 19348
rect 17126 19292 17164 19348
rect 17220 19292 17230 19348
rect 19618 19292 19628 19348
rect 19684 19292 20524 19348
rect 20580 19292 20590 19348
rect 20748 19292 24108 19348
rect 24164 19292 24174 19348
rect 26852 19236 26908 19404
rect 27010 19292 27020 19348
rect 27076 19292 28140 19348
rect 28196 19292 28700 19348
rect 28756 19292 30156 19348
rect 30212 19292 31276 19348
rect 31332 19292 33236 19348
rect 33842 19292 33852 19348
rect 33908 19292 34300 19348
rect 34356 19292 34366 19348
rect 37986 19292 37996 19348
rect 38052 19292 39900 19348
rect 39956 19292 39966 19348
rect 43698 19292 43708 19348
rect 43764 19292 44604 19348
rect 44660 19292 44670 19348
rect 46946 19292 46956 19348
rect 47012 19292 48188 19348
rect 48244 19292 48254 19348
rect 33180 19236 33236 19292
rect 8418 19180 8428 19236
rect 8484 19180 10668 19236
rect 10724 19180 11284 19236
rect 16370 19180 16380 19236
rect 16436 19180 17052 19236
rect 17108 19180 18508 19236
rect 18564 19180 18574 19236
rect 19730 19180 19740 19236
rect 19796 19180 20300 19236
rect 20356 19180 20366 19236
rect 21858 19180 21868 19236
rect 21924 19180 22092 19236
rect 22148 19180 22158 19236
rect 22754 19180 22764 19236
rect 22820 19180 23660 19236
rect 23716 19180 25116 19236
rect 25172 19180 25182 19236
rect 26852 19180 27580 19236
rect 27636 19180 27646 19236
rect 29474 19180 29484 19236
rect 29540 19180 30492 19236
rect 30548 19180 31612 19236
rect 31668 19180 32396 19236
rect 32452 19180 32462 19236
rect 33170 19180 33180 19236
rect 33236 19180 38668 19236
rect 11228 19124 11284 19180
rect 6038 19068 6076 19124
rect 6132 19068 6142 19124
rect 7746 19068 7756 19124
rect 7812 19068 9100 19124
rect 9156 19068 9166 19124
rect 11218 19068 11228 19124
rect 11284 19068 11294 19124
rect 11442 19068 11452 19124
rect 11508 19068 12460 19124
rect 12516 19068 12526 19124
rect 21746 19068 21756 19124
rect 21812 19068 23772 19124
rect 23828 19068 23838 19124
rect 31490 19068 31500 19124
rect 31556 19068 33068 19124
rect 33124 19068 33134 19124
rect 34962 19068 34972 19124
rect 35028 19068 36652 19124
rect 36708 19068 36718 19124
rect 38612 19012 38668 19180
rect 2370 18956 2380 19012
rect 2436 18956 6188 19012
rect 6244 18956 6254 19012
rect 16482 18956 16492 19012
rect 16548 18956 18508 19012
rect 18564 18956 20076 19012
rect 20132 18956 20142 19012
rect 21634 18956 21644 19012
rect 21700 18956 22428 19012
rect 22484 18956 22494 19012
rect 32162 18956 32172 19012
rect 32228 18956 32956 19012
rect 33012 18956 33022 19012
rect 33506 18956 33516 19012
rect 33572 18956 34524 19012
rect 34580 18956 35868 19012
rect 35924 18956 37100 19012
rect 37156 18956 37166 19012
rect 38612 18956 42924 19012
rect 42980 18956 42990 19012
rect 1250 18844 1260 18900
rect 1316 18844 5964 18900
rect 6020 18844 6356 18900
rect 12338 18844 12348 18900
rect 12404 18844 17668 18900
rect 18274 18844 18284 18900
rect 18340 18844 18396 18900
rect 18452 18844 18462 18900
rect 20514 18844 20524 18900
rect 20580 18844 22764 18900
rect 22820 18844 22830 18900
rect 26898 18844 26908 18900
rect 26964 18844 27692 18900
rect 27748 18844 27758 18900
rect 30258 18844 30268 18900
rect 30324 18844 34188 18900
rect 34244 18844 34254 18900
rect 45042 18844 45052 18900
rect 45108 18844 45118 18900
rect 6300 18788 6356 18844
rect 17612 18788 17668 18844
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 2706 18732 2716 18788
rect 2772 18732 3388 18788
rect 6300 18732 16828 18788
rect 16884 18732 17388 18788
rect 17444 18732 17454 18788
rect 17602 18732 17612 18788
rect 17668 18732 17706 18788
rect 20738 18732 20748 18788
rect 20804 18732 20860 18788
rect 20916 18732 23436 18788
rect 23492 18732 23502 18788
rect 23650 18732 23660 18788
rect 23716 18732 35644 18788
rect 35700 18732 35710 18788
rect 3332 18564 3388 18732
rect 6402 18620 6412 18676
rect 6468 18620 7084 18676
rect 7140 18620 7150 18676
rect 14550 18620 14588 18676
rect 14644 18620 14654 18676
rect 17378 18620 17388 18676
rect 17444 18620 18060 18676
rect 18116 18620 18126 18676
rect 23874 18620 23884 18676
rect 23940 18620 25116 18676
rect 25172 18620 25182 18676
rect 36642 18620 36652 18676
rect 36708 18620 38892 18676
rect 38948 18620 38958 18676
rect 3332 18508 6356 18564
rect 10770 18508 10780 18564
rect 10836 18508 11452 18564
rect 11508 18508 11518 18564
rect 15138 18508 15148 18564
rect 15204 18508 17948 18564
rect 18004 18508 21868 18564
rect 21924 18508 21934 18564
rect 22082 18508 22092 18564
rect 22148 18508 23996 18564
rect 24052 18508 24062 18564
rect 24434 18508 24444 18564
rect 24500 18508 29932 18564
rect 29988 18508 29998 18564
rect 31938 18508 31948 18564
rect 32004 18508 32956 18564
rect 33012 18508 33628 18564
rect 33684 18508 33694 18564
rect 37426 18508 37436 18564
rect 37492 18508 37660 18564
rect 37716 18508 39564 18564
rect 39620 18508 39630 18564
rect 6300 18452 6356 18508
rect 45052 18452 45108 18844
rect 45490 18508 45500 18564
rect 45556 18508 45836 18564
rect 45892 18508 45902 18564
rect 2034 18396 2044 18452
rect 2100 18396 2492 18452
rect 2548 18396 4284 18452
rect 4340 18396 5516 18452
rect 5572 18396 5582 18452
rect 6290 18396 6300 18452
rect 6356 18396 6366 18452
rect 6962 18396 6972 18452
rect 7028 18396 7644 18452
rect 7700 18396 7710 18452
rect 10182 18396 10220 18452
rect 10276 18396 10286 18452
rect 11778 18396 11788 18452
rect 11844 18396 14588 18452
rect 14644 18396 14654 18452
rect 15092 18396 17388 18452
rect 17444 18396 17454 18452
rect 18172 18396 20300 18452
rect 20356 18396 20366 18452
rect 23314 18396 23324 18452
rect 23380 18396 29596 18452
rect 29652 18396 31388 18452
rect 31444 18396 31454 18452
rect 33842 18396 33852 18452
rect 33908 18396 36988 18452
rect 37044 18396 37054 18452
rect 38994 18396 39004 18452
rect 39060 18396 41132 18452
rect 41188 18396 43820 18452
rect 43876 18396 43886 18452
rect 45052 18396 48076 18452
rect 48132 18396 48142 18452
rect 15092 18340 15148 18396
rect 18172 18340 18228 18396
rect 3826 18284 3836 18340
rect 3892 18284 7196 18340
rect 7252 18284 7262 18340
rect 10994 18284 11004 18340
rect 11060 18284 11340 18340
rect 11396 18284 12796 18340
rect 12852 18284 12862 18340
rect 13346 18284 13356 18340
rect 13412 18284 15148 18340
rect 16930 18284 16940 18340
rect 16996 18284 17612 18340
rect 17668 18284 17724 18340
rect 17780 18284 18228 18340
rect 18386 18284 18396 18340
rect 18452 18284 19404 18340
rect 19460 18284 19470 18340
rect 19730 18284 19740 18340
rect 19796 18284 21532 18340
rect 21588 18284 21598 18340
rect 23650 18284 23660 18340
rect 23716 18284 23726 18340
rect 24658 18284 24668 18340
rect 24724 18284 26012 18340
rect 26068 18284 26078 18340
rect 23660 18228 23716 18284
rect 29596 18228 29652 18396
rect 40338 18284 40348 18340
rect 40404 18284 41580 18340
rect 41636 18284 41646 18340
rect 42018 18284 42028 18340
rect 42084 18284 43036 18340
rect 43092 18284 43102 18340
rect 45938 18284 45948 18340
rect 46004 18284 47180 18340
rect 47236 18284 47964 18340
rect 48020 18284 48030 18340
rect 5730 18172 5740 18228
rect 5796 18172 8428 18228
rect 8484 18172 9660 18228
rect 9716 18172 12572 18228
rect 12628 18172 12638 18228
rect 17378 18172 17388 18228
rect 17444 18172 18060 18228
rect 18116 18172 22764 18228
rect 22820 18172 22830 18228
rect 23538 18172 23548 18228
rect 23604 18172 23716 18228
rect 23846 18172 23884 18228
rect 23940 18172 23950 18228
rect 29250 18172 29260 18228
rect 29316 18172 29652 18228
rect 1810 18060 1820 18116
rect 1876 18060 2828 18116
rect 2884 18060 3500 18116
rect 3556 18060 3566 18116
rect 4946 18060 4956 18116
rect 5012 18060 6524 18116
rect 6580 18060 6590 18116
rect 14578 18060 14588 18116
rect 14644 18060 22540 18116
rect 22596 18060 23100 18116
rect 23156 18060 23166 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 5170 17948 5180 18004
rect 5236 17948 5852 18004
rect 5908 17948 5918 18004
rect 7522 17948 7532 18004
rect 7588 17948 8092 18004
rect 8148 17948 8158 18004
rect 17378 17948 17388 18004
rect 17444 17948 20748 18004
rect 20804 17948 20814 18004
rect 24210 17948 24220 18004
rect 24276 17948 24780 18004
rect 24836 17948 31500 18004
rect 31556 17948 34972 18004
rect 35028 17948 35038 18004
rect 38612 17948 42700 18004
rect 42756 17948 42766 18004
rect 38612 17892 38668 17948
rect 2930 17836 2940 17892
rect 2996 17836 4396 17892
rect 4452 17836 4462 17892
rect 4834 17836 4844 17892
rect 4900 17836 10220 17892
rect 10276 17836 10286 17892
rect 10892 17836 12236 17892
rect 12292 17836 13244 17892
rect 13300 17836 13310 17892
rect 19842 17836 19852 17892
rect 19908 17836 20412 17892
rect 20468 17836 20478 17892
rect 20626 17836 20636 17892
rect 20692 17836 21980 17892
rect 22036 17836 22046 17892
rect 26852 17836 29148 17892
rect 29204 17836 38668 17892
rect 10892 17780 10948 17836
rect 26852 17780 26908 17836
rect 3332 17724 10948 17780
rect 11666 17724 11676 17780
rect 11732 17724 14140 17780
rect 14196 17724 14206 17780
rect 14354 17724 14364 17780
rect 14420 17724 16156 17780
rect 16212 17724 18284 17780
rect 18340 17724 18350 17780
rect 20132 17724 26908 17780
rect 31154 17724 31164 17780
rect 31220 17724 33292 17780
rect 33348 17724 33852 17780
rect 33908 17724 33918 17780
rect 43026 17724 43036 17780
rect 43092 17724 44044 17780
rect 44100 17724 44110 17780
rect 3266 17388 3276 17444
rect 3332 17388 3388 17724
rect 3938 17612 3948 17668
rect 4004 17612 4844 17668
rect 4900 17612 4910 17668
rect 5506 17612 5516 17668
rect 5572 17612 8204 17668
rect 8260 17612 8270 17668
rect 11778 17612 11788 17668
rect 11844 17612 14924 17668
rect 14980 17612 14990 17668
rect 18162 17612 18172 17668
rect 18228 17612 19628 17668
rect 19684 17612 19694 17668
rect 20132 17556 20188 17724
rect 22754 17612 22764 17668
rect 22820 17612 23436 17668
rect 23492 17612 23502 17668
rect 24658 17612 24668 17668
rect 24724 17612 25900 17668
rect 25956 17612 25966 17668
rect 34514 17612 34524 17668
rect 34580 17612 36316 17668
rect 36372 17612 36382 17668
rect 38994 17612 39004 17668
rect 39060 17612 40012 17668
rect 40068 17612 40908 17668
rect 40964 17612 41916 17668
rect 41972 17612 41982 17668
rect 43586 17612 43596 17668
rect 43652 17612 44716 17668
rect 44772 17612 44782 17668
rect 44940 17612 45388 17668
rect 45444 17612 45454 17668
rect 44940 17556 44996 17612
rect 49200 17556 50000 17584
rect 5394 17500 5404 17556
rect 5460 17500 6300 17556
rect 6356 17500 6366 17556
rect 7746 17500 7756 17556
rect 7812 17500 8988 17556
rect 9044 17500 9054 17556
rect 10098 17500 10108 17556
rect 10164 17500 12572 17556
rect 12628 17500 12638 17556
rect 14690 17500 14700 17556
rect 14756 17500 16716 17556
rect 16772 17500 16782 17556
rect 18508 17500 20188 17556
rect 23426 17500 23436 17556
rect 23492 17500 24108 17556
rect 24164 17500 24174 17556
rect 28326 17500 28364 17556
rect 28420 17500 28430 17556
rect 33618 17500 33628 17556
rect 33684 17500 34188 17556
rect 34244 17500 34254 17556
rect 43138 17500 43148 17556
rect 43204 17500 43372 17556
rect 43428 17500 44996 17556
rect 45154 17500 45164 17556
rect 45220 17500 45612 17556
rect 45668 17500 45678 17556
rect 46274 17500 46284 17556
rect 46340 17500 47068 17556
rect 47124 17500 47134 17556
rect 47506 17500 47516 17556
rect 47572 17500 47582 17556
rect 48066 17500 48076 17556
rect 48132 17500 50000 17556
rect 7186 17388 7196 17444
rect 7252 17388 7644 17444
rect 7700 17388 7710 17444
rect 7858 17388 7868 17444
rect 7924 17388 12124 17444
rect 12180 17388 12190 17444
rect 18508 17332 18564 17500
rect 47516 17444 47572 17500
rect 49200 17472 50000 17500
rect 19506 17388 19516 17444
rect 19572 17388 20076 17444
rect 20132 17388 20142 17444
rect 20626 17388 20636 17444
rect 20692 17388 24556 17444
rect 24612 17388 25116 17444
rect 25172 17388 25182 17444
rect 25778 17388 25788 17444
rect 25844 17388 47572 17444
rect 7298 17276 7308 17332
rect 7364 17276 10108 17332
rect 10164 17276 10174 17332
rect 13468 17276 18564 17332
rect 26002 17276 26012 17332
rect 26068 17276 28924 17332
rect 28980 17276 28990 17332
rect 13468 17220 13524 17276
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 1474 17164 1484 17220
rect 1540 17164 3724 17220
rect 3780 17164 3790 17220
rect 4946 17164 4956 17220
rect 5012 17164 7420 17220
rect 7476 17164 7486 17220
rect 10108 17164 13468 17220
rect 13524 17164 13534 17220
rect 13794 17164 13804 17220
rect 13860 17164 14700 17220
rect 14756 17164 14766 17220
rect 18834 17164 18844 17220
rect 18900 17164 19628 17220
rect 19684 17164 19694 17220
rect 20178 17164 20188 17220
rect 20244 17164 22484 17220
rect 24658 17164 24668 17220
rect 24724 17164 27132 17220
rect 27188 17164 27198 17220
rect 10108 17108 10164 17164
rect 22428 17108 22484 17164
rect 2268 17052 4004 17108
rect 2268 16884 2324 17052
rect 3948 16996 4004 17052
rect 5628 17052 10108 17108
rect 10164 17052 10174 17108
rect 11442 17052 11452 17108
rect 11508 17052 17276 17108
rect 17332 17052 17342 17108
rect 17490 17052 17500 17108
rect 17556 17052 17948 17108
rect 18004 17052 18284 17108
rect 18340 17052 18620 17108
rect 18676 17052 18686 17108
rect 19058 17052 19068 17108
rect 19124 17052 20412 17108
rect 20468 17052 20478 17108
rect 22418 17052 22428 17108
rect 22484 17052 22494 17108
rect 22754 17052 22764 17108
rect 22820 17052 24332 17108
rect 24388 17052 24398 17108
rect 24770 17052 24780 17108
rect 24836 17052 26348 17108
rect 26404 17052 27692 17108
rect 27748 17052 27758 17108
rect 38322 17052 38332 17108
rect 38388 17052 40236 17108
rect 40292 17052 40302 17108
rect 5628 16996 5684 17052
rect 3154 16940 3164 16996
rect 3220 16940 3612 16996
rect 3668 16940 3678 16996
rect 3948 16940 5684 16996
rect 5740 16940 7196 16996
rect 7252 16940 7262 16996
rect 9996 16940 14364 16996
rect 14420 16940 14430 16996
rect 14802 16940 14812 16996
rect 14868 16940 16044 16996
rect 16100 16940 20076 16996
rect 20132 16940 20636 16996
rect 20692 16940 28812 16996
rect 28868 16940 33068 16996
rect 33124 16940 37100 16996
rect 37156 16940 37772 16996
rect 37828 16940 39004 16996
rect 39060 16940 39070 16996
rect 5740 16884 5796 16940
rect 2258 16828 2268 16884
rect 2324 16828 2334 16884
rect 2594 16828 2604 16884
rect 2660 16828 3500 16884
rect 3556 16828 3566 16884
rect 3826 16828 3836 16884
rect 3892 16828 4060 16884
rect 4116 16828 4126 16884
rect 4946 16828 4956 16884
rect 5012 16828 5068 16884
rect 5124 16828 5134 16884
rect 5730 16828 5740 16884
rect 5796 16828 5806 16884
rect 6626 16828 6636 16884
rect 6692 16828 8428 16884
rect 8484 16828 8494 16884
rect 9996 16772 10052 16940
rect 11218 16828 11228 16884
rect 11284 16828 13804 16884
rect 13860 16828 15372 16884
rect 15428 16828 16156 16884
rect 16212 16828 16222 16884
rect 18050 16828 18060 16884
rect 18116 16828 18396 16884
rect 18452 16828 18462 16884
rect 22530 16828 22540 16884
rect 22596 16828 22988 16884
rect 23044 16828 23054 16884
rect 23762 16828 23772 16884
rect 23828 16828 24780 16884
rect 24836 16828 24846 16884
rect 25750 16828 25788 16884
rect 25844 16828 25854 16884
rect 26562 16828 26572 16884
rect 26628 16828 26908 16884
rect 26964 16828 28476 16884
rect 28532 16828 28542 16884
rect 28690 16828 28700 16884
rect 28756 16828 28924 16884
rect 28980 16828 30044 16884
rect 30100 16828 30110 16884
rect 31266 16828 31276 16884
rect 31332 16828 32060 16884
rect 32116 16828 32126 16884
rect 35410 16828 35420 16884
rect 35476 16828 36092 16884
rect 36148 16828 36158 16884
rect 36530 16828 36540 16884
rect 36596 16828 36988 16884
rect 37044 16828 38444 16884
rect 38500 16828 38510 16884
rect 40114 16828 40124 16884
rect 40180 16828 40908 16884
rect 40964 16828 42028 16884
rect 42084 16828 44156 16884
rect 44212 16828 45276 16884
rect 45332 16828 45342 16884
rect 46050 16828 46060 16884
rect 46116 16828 47516 16884
rect 47572 16828 47582 16884
rect 3154 16716 3164 16772
rect 3220 16716 10052 16772
rect 13122 16716 13132 16772
rect 13188 16716 14588 16772
rect 14644 16716 14654 16772
rect 15698 16716 15708 16772
rect 15764 16716 17500 16772
rect 17556 16716 17566 16772
rect 25218 16716 25228 16772
rect 25284 16716 27468 16772
rect 27524 16716 27534 16772
rect 28578 16716 28588 16772
rect 28644 16716 29148 16772
rect 29204 16716 29214 16772
rect 30370 16716 30380 16772
rect 30436 16716 31500 16772
rect 31556 16716 31566 16772
rect 38994 16716 39004 16772
rect 39060 16716 43932 16772
rect 43988 16716 43998 16772
rect 45826 16716 45836 16772
rect 45892 16716 46396 16772
rect 46452 16716 46462 16772
rect 4050 16604 4060 16660
rect 4116 16604 6076 16660
rect 6132 16604 6142 16660
rect 8642 16604 8652 16660
rect 8708 16604 10332 16660
rect 10388 16604 10398 16660
rect 23538 16604 23548 16660
rect 23604 16604 24108 16660
rect 24164 16604 27132 16660
rect 27188 16604 27916 16660
rect 27972 16604 28364 16660
rect 28420 16604 28430 16660
rect 4918 16492 4956 16548
rect 5012 16492 5022 16548
rect 18274 16492 18284 16548
rect 18340 16492 33068 16548
rect 33124 16492 33134 16548
rect 37314 16492 37324 16548
rect 37380 16492 43036 16548
rect 43092 16492 43102 16548
rect 46946 16492 46956 16548
rect 47012 16492 47628 16548
rect 47684 16492 47694 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 4844 16380 14700 16436
rect 14756 16380 14766 16436
rect 17462 16380 17500 16436
rect 17556 16380 17566 16436
rect 21410 16380 21420 16436
rect 21476 16380 23100 16436
rect 23156 16380 23166 16436
rect 26674 16380 26684 16436
rect 26740 16380 27580 16436
rect 27636 16380 27646 16436
rect 37202 16380 37212 16436
rect 37268 16380 39788 16436
rect 39844 16380 39854 16436
rect 4844 16324 4900 16380
rect 4050 16268 4060 16324
rect 4116 16268 4900 16324
rect 12450 16268 12460 16324
rect 12516 16268 14140 16324
rect 14196 16268 14206 16324
rect 16482 16268 16492 16324
rect 16548 16268 18732 16324
rect 18788 16268 18798 16324
rect 23314 16268 23324 16324
rect 23380 16268 26796 16324
rect 26852 16268 26862 16324
rect 3266 16156 3276 16212
rect 3332 16156 6076 16212
rect 6132 16156 6142 16212
rect 7186 16156 7196 16212
rect 7252 16156 16436 16212
rect 16594 16156 16604 16212
rect 16660 16156 22764 16212
rect 22820 16156 23884 16212
rect 23940 16156 23950 16212
rect 36306 16156 36316 16212
rect 36372 16156 39228 16212
rect 39284 16156 39294 16212
rect 16380 16100 16436 16156
rect 4386 16044 4396 16100
rect 4452 16044 5068 16100
rect 5124 16044 5134 16100
rect 6626 16044 6636 16100
rect 6692 16044 7308 16100
rect 7364 16044 7374 16100
rect 10322 16044 10332 16100
rect 10388 16044 11900 16100
rect 11956 16044 11966 16100
rect 16380 16044 19404 16100
rect 19460 16044 19470 16100
rect 20402 16044 20412 16100
rect 20468 16044 24220 16100
rect 24276 16044 24286 16100
rect 25218 16044 25228 16100
rect 25284 16044 25564 16100
rect 25620 16044 30268 16100
rect 30324 16044 30334 16100
rect 30818 16044 30828 16100
rect 30884 16044 32732 16100
rect 32788 16044 32798 16100
rect 33058 16044 33068 16100
rect 33124 16044 37716 16100
rect 37874 16044 37884 16100
rect 37940 16044 39340 16100
rect 39396 16044 39406 16100
rect 42914 16044 42924 16100
rect 42980 16044 43708 16100
rect 43764 16044 43774 16100
rect 44034 16044 44044 16100
rect 44100 16044 45052 16100
rect 45108 16044 45118 16100
rect 37660 15988 37716 16044
rect 3938 15932 3948 15988
rect 4004 15932 4284 15988
rect 4340 15932 4844 15988
rect 4900 15932 4910 15988
rect 5618 15932 5628 15988
rect 5684 15932 6300 15988
rect 6356 15932 6366 15988
rect 6738 15932 6748 15988
rect 6804 15932 7644 15988
rect 7700 15932 7710 15988
rect 10434 15932 10444 15988
rect 10500 15932 13580 15988
rect 13636 15932 13646 15988
rect 16706 15932 16716 15988
rect 16772 15932 17612 15988
rect 17668 15932 20524 15988
rect 20580 15932 20590 15988
rect 20738 15932 20748 15988
rect 20804 15932 20842 15988
rect 21746 15932 21756 15988
rect 21812 15932 22876 15988
rect 22932 15932 22942 15988
rect 24322 15932 24332 15988
rect 24388 15932 25340 15988
rect 25396 15932 25900 15988
rect 25956 15932 25966 15988
rect 29362 15932 29372 15988
rect 29428 15932 32620 15988
rect 32676 15932 32686 15988
rect 34290 15932 34300 15988
rect 34356 15932 35308 15988
rect 35364 15932 35374 15988
rect 37650 15932 37660 15988
rect 37716 15932 37726 15988
rect 38098 15932 38108 15988
rect 38164 15932 38780 15988
rect 38836 15932 38846 15988
rect 2706 15820 2716 15876
rect 2772 15820 3388 15876
rect 4946 15820 4956 15876
rect 5012 15820 5022 15876
rect 6150 15820 6188 15876
rect 6244 15820 6860 15876
rect 6916 15820 12348 15876
rect 12404 15820 12414 15876
rect 19730 15820 19740 15876
rect 19796 15820 24892 15876
rect 24948 15820 24958 15876
rect 27906 15820 27916 15876
rect 27972 15820 31612 15876
rect 31668 15820 31678 15876
rect 31938 15820 31948 15876
rect 32004 15820 33628 15876
rect 33684 15820 33694 15876
rect 3332 15652 3388 15820
rect 4956 15764 5012 15820
rect 37660 15764 37716 15932
rect 37986 15820 37996 15876
rect 38052 15820 39676 15876
rect 39732 15820 39742 15876
rect 41244 15820 41916 15876
rect 41972 15820 42476 15876
rect 42532 15820 42542 15876
rect 41244 15764 41300 15820
rect 4956 15708 7868 15764
rect 7924 15708 7934 15764
rect 12348 15708 15036 15764
rect 15092 15708 15102 15764
rect 21410 15708 21420 15764
rect 21476 15708 22428 15764
rect 22484 15708 22494 15764
rect 23762 15708 23772 15764
rect 23828 15708 24668 15764
rect 24724 15708 24734 15764
rect 28578 15708 28588 15764
rect 28644 15708 32172 15764
rect 32228 15708 32238 15764
rect 37660 15708 38668 15764
rect 38724 15708 38734 15764
rect 41234 15708 41244 15764
rect 41300 15708 41310 15764
rect 12348 15652 12404 15708
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 3332 15596 3500 15652
rect 3556 15596 9884 15652
rect 9940 15596 9950 15652
rect 12338 15596 12348 15652
rect 12404 15596 12414 15652
rect 12674 15596 12684 15652
rect 12740 15596 17052 15652
rect 17108 15596 17118 15652
rect 18246 15596 18284 15652
rect 18340 15596 18350 15652
rect 24332 15596 34860 15652
rect 34916 15596 34926 15652
rect 35410 15596 35420 15652
rect 35476 15596 35868 15652
rect 35924 15596 38220 15652
rect 38276 15596 38286 15652
rect 24332 15540 24388 15596
rect 3938 15484 3948 15540
rect 4004 15484 4620 15540
rect 4676 15484 5292 15540
rect 5348 15484 8596 15540
rect 13234 15484 13244 15540
rect 13300 15484 16268 15540
rect 16324 15484 16334 15540
rect 17490 15484 17500 15540
rect 17556 15484 17566 15540
rect 19058 15484 19068 15540
rect 19124 15484 20748 15540
rect 20804 15484 20814 15540
rect 24322 15484 24332 15540
rect 24388 15484 24398 15540
rect 27234 15484 27244 15540
rect 27300 15484 33180 15540
rect 33236 15484 35756 15540
rect 35812 15484 35822 15540
rect 35970 15484 35980 15540
rect 36036 15484 37324 15540
rect 37380 15484 37390 15540
rect 39890 15484 39900 15540
rect 39956 15484 40236 15540
rect 40292 15484 40302 15540
rect 43138 15484 43148 15540
rect 43204 15484 43484 15540
rect 43540 15484 43932 15540
rect 43988 15484 43998 15540
rect 8540 15428 8596 15484
rect 17500 15428 17556 15484
rect 24332 15428 24388 15484
rect 5506 15372 5516 15428
rect 5572 15372 7420 15428
rect 7476 15372 8316 15428
rect 8372 15372 8382 15428
rect 8540 15372 17556 15428
rect 19628 15372 24388 15428
rect 27346 15372 27356 15428
rect 27412 15372 33404 15428
rect 33460 15372 35644 15428
rect 35700 15372 35710 15428
rect 41010 15372 41020 15428
rect 41076 15372 41692 15428
rect 41748 15372 41758 15428
rect 45938 15372 45948 15428
rect 46004 15372 47404 15428
rect 47460 15372 47470 15428
rect 6374 15260 6412 15316
rect 6468 15260 6478 15316
rect 7858 15260 7868 15316
rect 7924 15260 8764 15316
rect 8820 15260 8830 15316
rect 13906 15260 13916 15316
rect 13972 15260 15820 15316
rect 15876 15260 15886 15316
rect 17042 15260 17052 15316
rect 17108 15260 19404 15316
rect 19460 15260 19470 15316
rect 19628 15204 19684 15372
rect 20850 15260 20860 15316
rect 20916 15260 25340 15316
rect 25396 15260 25406 15316
rect 27458 15260 27468 15316
rect 27524 15260 28364 15316
rect 28420 15260 32060 15316
rect 32116 15260 36428 15316
rect 36484 15260 36494 15316
rect 42802 15260 42812 15316
rect 42868 15260 44380 15316
rect 44436 15260 44716 15316
rect 44772 15260 44782 15316
rect 45378 15260 45388 15316
rect 45444 15260 46284 15316
rect 46340 15260 46844 15316
rect 46900 15260 47964 15316
rect 48020 15260 48030 15316
rect 1026 15148 1036 15204
rect 1092 15148 6300 15204
rect 6356 15148 7196 15204
rect 7252 15148 7262 15204
rect 7970 15148 7980 15204
rect 8036 15148 8988 15204
rect 9044 15148 9940 15204
rect 11778 15148 11788 15204
rect 11844 15148 13468 15204
rect 13524 15148 13534 15204
rect 15922 15148 15932 15204
rect 15988 15148 16492 15204
rect 16548 15148 17164 15204
rect 17220 15148 19684 15204
rect 21868 15148 24444 15204
rect 24500 15148 25228 15204
rect 25284 15148 25294 15204
rect 31938 15148 31948 15204
rect 32004 15148 32844 15204
rect 32900 15148 35980 15204
rect 36036 15148 36046 15204
rect 38770 15148 38780 15204
rect 38836 15148 39900 15204
rect 39956 15148 39966 15204
rect 42130 15148 42140 15204
rect 42196 15148 43148 15204
rect 43204 15148 45500 15204
rect 45556 15148 45836 15204
rect 45892 15148 45902 15204
rect 9884 15092 9940 15148
rect 21868 15092 21924 15148
rect 2818 15036 2828 15092
rect 2884 15036 8596 15092
rect 9874 15036 9884 15092
rect 9940 15036 9950 15092
rect 17938 15036 17948 15092
rect 18004 15036 20972 15092
rect 21028 15036 21756 15092
rect 21812 15036 21924 15092
rect 30482 15036 30492 15092
rect 30548 15036 31164 15092
rect 31220 15036 31230 15092
rect 8540 14980 8596 15036
rect 5394 14924 5404 14980
rect 5460 14924 6300 14980
rect 6356 14924 6366 14980
rect 8540 14924 10220 14980
rect 10276 14924 10668 14980
rect 10724 14924 10734 14980
rect 12562 14924 12572 14980
rect 12628 14924 15148 14980
rect 21634 14924 21644 14980
rect 21700 14924 22316 14980
rect 22372 14924 22382 14980
rect 27122 14924 27132 14980
rect 27188 14924 28700 14980
rect 28756 14924 28766 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 5282 14812 5292 14868
rect 5348 14812 6524 14868
rect 6580 14812 6590 14868
rect 11554 14812 11564 14868
rect 11620 14812 12684 14868
rect 12740 14812 12750 14868
rect 15092 14756 15148 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 19618 14812 19628 14868
rect 19684 14812 26012 14868
rect 26068 14812 26078 14868
rect 26450 14812 26460 14868
rect 26516 14812 28140 14868
rect 28196 14812 28206 14868
rect 28578 14812 28588 14868
rect 28644 14812 30156 14868
rect 30212 14812 30828 14868
rect 30884 14812 30894 14868
rect 4162 14700 4172 14756
rect 4228 14700 5516 14756
rect 5572 14700 5582 14756
rect 5954 14700 5964 14756
rect 6020 14700 8316 14756
rect 8372 14700 8382 14756
rect 9212 14700 9996 14756
rect 10052 14700 10444 14756
rect 10500 14700 10510 14756
rect 10882 14700 10892 14756
rect 10948 14700 11900 14756
rect 11956 14700 11966 14756
rect 12226 14700 12236 14756
rect 12292 14700 12852 14756
rect 15092 14700 16492 14756
rect 16548 14700 16558 14756
rect 19618 14700 19628 14756
rect 19684 14700 23884 14756
rect 23940 14700 23950 14756
rect 27570 14700 27580 14756
rect 27636 14700 28644 14756
rect 29698 14700 29708 14756
rect 29764 14700 30380 14756
rect 30436 14700 30446 14756
rect 30604 14700 45612 14756
rect 45668 14700 45678 14756
rect 9212 14644 9268 14700
rect 12796 14644 12852 14700
rect 28588 14644 28644 14700
rect 30604 14644 30660 14700
rect 4834 14588 4844 14644
rect 4900 14588 6076 14644
rect 6132 14588 6142 14644
rect 7532 14588 9268 14644
rect 9426 14588 9436 14644
rect 9492 14588 11228 14644
rect 11284 14588 11294 14644
rect 12796 14588 18396 14644
rect 18452 14588 18462 14644
rect 20738 14588 20748 14644
rect 20804 14588 22092 14644
rect 22148 14588 22158 14644
rect 22316 14588 28028 14644
rect 28084 14588 28364 14644
rect 28420 14588 28430 14644
rect 28578 14588 28588 14644
rect 28644 14588 30660 14644
rect 33618 14588 33628 14644
rect 33684 14588 35980 14644
rect 36036 14588 36046 14644
rect 7532 14532 7588 14588
rect 22316 14532 22372 14588
rect 5058 14476 5068 14532
rect 5124 14476 7588 14532
rect 7746 14476 7756 14532
rect 7812 14476 9212 14532
rect 9268 14476 9278 14532
rect 11106 14476 11116 14532
rect 11172 14476 12572 14532
rect 12628 14476 12638 14532
rect 16594 14476 16604 14532
rect 16660 14476 18508 14532
rect 18564 14476 18574 14532
rect 18844 14476 21196 14532
rect 21252 14476 22372 14532
rect 24882 14476 24892 14532
rect 24948 14476 25452 14532
rect 25508 14476 25518 14532
rect 25778 14476 25788 14532
rect 25844 14476 27692 14532
rect 27748 14476 27758 14532
rect 28130 14476 28140 14532
rect 28196 14476 34188 14532
rect 34244 14476 34254 14532
rect 34514 14476 34524 14532
rect 34580 14476 36540 14532
rect 36596 14476 36606 14532
rect 37314 14476 37324 14532
rect 37380 14476 38892 14532
rect 38948 14476 38958 14532
rect 40898 14476 40908 14532
rect 40964 14476 43708 14532
rect 43764 14476 43774 14532
rect 43922 14476 43932 14532
rect 43988 14476 44268 14532
rect 44324 14476 44334 14532
rect 1362 14364 1372 14420
rect 1428 14364 2716 14420
rect 2772 14364 2782 14420
rect 4806 14364 4844 14420
rect 4900 14364 4910 14420
rect 5394 14364 5404 14420
rect 5460 14364 5964 14420
rect 6020 14364 6030 14420
rect 6402 14364 6412 14420
rect 6468 14364 6636 14420
rect 6692 14364 6702 14420
rect 8194 14364 8204 14420
rect 8260 14364 9100 14420
rect 9156 14364 9772 14420
rect 9828 14364 9838 14420
rect 12786 14364 12796 14420
rect 12852 14364 14252 14420
rect 14308 14364 14318 14420
rect 17714 14364 17724 14420
rect 17780 14364 18620 14420
rect 18676 14364 18686 14420
rect 18844 14308 18900 14476
rect 21718 14364 21756 14420
rect 21812 14364 21822 14420
rect 23090 14364 23100 14420
rect 23156 14364 23436 14420
rect 23492 14364 27860 14420
rect 34962 14364 34972 14420
rect 35028 14364 36316 14420
rect 36372 14364 36876 14420
rect 36932 14364 38220 14420
rect 38276 14364 38286 14420
rect 46050 14364 46060 14420
rect 46116 14364 46956 14420
rect 47012 14364 47022 14420
rect 4162 14252 4172 14308
rect 4228 14252 5740 14308
rect 5796 14252 5806 14308
rect 6066 14252 6076 14308
rect 6132 14252 6524 14308
rect 6580 14252 7980 14308
rect 8036 14252 8046 14308
rect 12114 14252 12124 14308
rect 12180 14252 12908 14308
rect 12964 14252 14812 14308
rect 14868 14252 14878 14308
rect 15092 14252 15316 14308
rect 16482 14252 16492 14308
rect 16548 14252 18900 14308
rect 20290 14252 20300 14308
rect 20356 14252 23884 14308
rect 23940 14252 23950 14308
rect 25106 14252 25116 14308
rect 25172 14252 26348 14308
rect 26404 14252 26684 14308
rect 26740 14252 26750 14308
rect 15092 14196 15148 14252
rect 7858 14140 7868 14196
rect 7924 14140 14476 14196
rect 14532 14140 15148 14196
rect 15260 14196 15316 14252
rect 27804 14196 27860 14364
rect 35410 14252 35420 14308
rect 35476 14252 37660 14308
rect 37716 14252 37726 14308
rect 37874 14252 37884 14308
rect 37940 14252 40908 14308
rect 40964 14252 40974 14308
rect 15260 14140 16604 14196
rect 16660 14140 18620 14196
rect 18676 14140 19628 14196
rect 19684 14140 19694 14196
rect 22092 14140 25956 14196
rect 26562 14140 26572 14196
rect 26628 14140 27580 14196
rect 27636 14140 27646 14196
rect 27804 14140 29372 14196
rect 29428 14140 30380 14196
rect 30436 14140 30828 14196
rect 30884 14140 30894 14196
rect 32498 14140 32508 14196
rect 32564 14140 35868 14196
rect 35924 14140 35934 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 22092 14084 22148 14140
rect 25900 14084 25956 14140
rect 7494 14028 7532 14084
rect 7588 14028 12236 14084
rect 12292 14028 12302 14084
rect 13766 14028 13804 14084
rect 13860 14028 17780 14084
rect 20402 14028 20412 14084
rect 20468 14028 21196 14084
rect 21252 14028 21262 14084
rect 22082 14028 22092 14084
rect 22148 14028 22158 14084
rect 1474 13916 1484 13972
rect 1540 13916 2268 13972
rect 2324 13916 2334 13972
rect 7970 13916 7980 13972
rect 8036 13916 8484 13972
rect 8642 13916 8652 13972
rect 8708 13916 9100 13972
rect 9156 13916 9166 13972
rect 15250 13916 15260 13972
rect 15316 13916 15708 13972
rect 15764 13916 16940 13972
rect 16996 13916 17006 13972
rect 8428 13748 8484 13916
rect 17724 13860 17780 14028
rect 19730 13916 19740 13972
rect 19796 13916 20748 13972
rect 20804 13916 20814 13972
rect 22530 13916 22540 13972
rect 22596 13916 23324 13972
rect 23380 13916 23390 13972
rect 23492 13860 23548 14084
rect 23604 14028 25676 14084
rect 25732 14028 25742 14084
rect 25900 14028 31612 14084
rect 31668 14028 32396 14084
rect 32452 14028 36988 14084
rect 37044 14028 37054 14084
rect 38434 14028 38444 14084
rect 38500 14028 40572 14084
rect 40628 14028 41020 14084
rect 41076 14028 41086 14084
rect 25106 13916 25116 13972
rect 25172 13916 26124 13972
rect 26180 13916 26190 13972
rect 28690 13916 28700 13972
rect 28756 13916 29372 13972
rect 29428 13916 29438 13972
rect 30034 13916 30044 13972
rect 30100 13916 30110 13972
rect 38612 13916 43260 13972
rect 43316 13916 43326 13972
rect 30044 13860 30100 13916
rect 38612 13860 38668 13916
rect 10182 13804 10220 13860
rect 10276 13804 14308 13860
rect 16258 13804 16268 13860
rect 16324 13804 17276 13860
rect 17332 13804 17500 13860
rect 17556 13804 17566 13860
rect 17724 13804 23548 13860
rect 23650 13804 23660 13860
rect 23716 13804 26908 13860
rect 26964 13804 26974 13860
rect 27570 13804 27580 13860
rect 27636 13804 30100 13860
rect 30940 13804 38668 13860
rect 3154 13692 3164 13748
rect 3220 13692 5068 13748
rect 5124 13692 5134 13748
rect 8418 13692 8428 13748
rect 8484 13692 8494 13748
rect 10658 13692 10668 13748
rect 10724 13692 13916 13748
rect 13972 13692 13982 13748
rect 14252 13636 14308 13804
rect 30940 13748 30996 13804
rect 15362 13692 15372 13748
rect 15428 13692 16492 13748
rect 16548 13692 16558 13748
rect 17714 13692 17724 13748
rect 17780 13692 19404 13748
rect 19460 13692 19470 13748
rect 21522 13692 21532 13748
rect 21588 13692 22876 13748
rect 22932 13692 23212 13748
rect 23268 13692 23278 13748
rect 23538 13692 23548 13748
rect 23604 13692 24108 13748
rect 24164 13692 25004 13748
rect 25060 13692 27468 13748
rect 27524 13692 30996 13748
rect 33282 13692 33292 13748
rect 33348 13692 33964 13748
rect 34020 13692 34030 13748
rect 34738 13692 34748 13748
rect 34804 13692 35420 13748
rect 35476 13692 35486 13748
rect 36082 13692 36092 13748
rect 36148 13692 37100 13748
rect 37156 13692 38444 13748
rect 38500 13692 38510 13748
rect 38602 13692 38612 13748
rect 38668 13692 39228 13748
rect 39284 13692 40236 13748
rect 40292 13692 40302 13748
rect 46946 13692 46956 13748
rect 47012 13692 47852 13748
rect 47908 13692 47918 13748
rect 3602 13580 3612 13636
rect 3668 13580 10892 13636
rect 10948 13580 11116 13636
rect 11172 13580 11182 13636
rect 11330 13580 11340 13636
rect 11396 13580 12124 13636
rect 12180 13580 12190 13636
rect 14252 13580 14364 13636
rect 14420 13580 15036 13636
rect 15092 13580 22092 13636
rect 22148 13580 22316 13636
rect 22372 13580 22382 13636
rect 25526 13580 25564 13636
rect 25620 13580 25630 13636
rect 25778 13580 25788 13636
rect 25844 13580 27020 13636
rect 27076 13580 27086 13636
rect 31126 13580 31164 13636
rect 31220 13580 31230 13636
rect 36530 13580 36540 13636
rect 36596 13580 39452 13636
rect 39508 13580 39518 13636
rect 4610 13468 4620 13524
rect 4676 13468 5292 13524
rect 5348 13468 5516 13524
rect 5572 13468 5582 13524
rect 6290 13468 6300 13524
rect 6356 13468 6972 13524
rect 7028 13468 7644 13524
rect 7700 13468 7710 13524
rect 7970 13468 7980 13524
rect 8036 13468 8540 13524
rect 8596 13468 8606 13524
rect 9090 13468 9100 13524
rect 9156 13468 15484 13524
rect 15540 13468 17948 13524
rect 18004 13468 18844 13524
rect 18900 13468 20860 13524
rect 20916 13468 20926 13524
rect 21410 13468 21420 13524
rect 21476 13468 22540 13524
rect 22596 13468 22606 13524
rect 25442 13468 25452 13524
rect 25508 13468 25676 13524
rect 25732 13468 25742 13524
rect 26310 13468 26348 13524
rect 26404 13468 26414 13524
rect 26898 13468 26908 13524
rect 26964 13468 32060 13524
rect 32116 13468 33180 13524
rect 33236 13468 33246 13524
rect 34514 13468 34524 13524
rect 34580 13468 35196 13524
rect 35252 13468 37772 13524
rect 37828 13468 39676 13524
rect 39732 13468 39742 13524
rect 40898 13468 40908 13524
rect 40964 13468 42868 13524
rect 42812 13412 42868 13468
rect 14018 13356 14028 13412
rect 14084 13356 16716 13412
rect 16772 13356 16782 13412
rect 23762 13356 23772 13412
rect 23828 13356 27356 13412
rect 27412 13356 27422 13412
rect 34374 13356 34412 13412
rect 34468 13356 34478 13412
rect 42802 13356 42812 13412
rect 42868 13356 42878 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 6374 13244 6412 13300
rect 6468 13244 6478 13300
rect 11218 13244 11228 13300
rect 11284 13244 13804 13300
rect 13860 13244 13870 13300
rect 14242 13244 14252 13300
rect 14308 13244 18060 13300
rect 18116 13244 18126 13300
rect 22838 13244 22876 13300
rect 22932 13244 24332 13300
rect 24388 13244 24398 13300
rect 25638 13244 25676 13300
rect 25732 13244 25742 13300
rect 26562 13244 26572 13300
rect 26628 13244 27412 13300
rect 39554 13244 39564 13300
rect 39620 13244 41020 13300
rect 41076 13244 41086 13300
rect 13804 13188 13860 13244
rect 27356 13188 27412 13244
rect 3266 13132 3276 13188
rect 3332 13132 5852 13188
rect 5908 13132 5918 13188
rect 8642 13132 8652 13188
rect 8708 13132 9884 13188
rect 9940 13132 10556 13188
rect 10612 13132 10622 13188
rect 13804 13132 14364 13188
rect 14420 13132 14430 13188
rect 16930 13132 16940 13188
rect 16996 13132 19180 13188
rect 19236 13132 19246 13188
rect 23090 13132 23100 13188
rect 23156 13132 26908 13188
rect 27346 13132 27356 13188
rect 27412 13132 34188 13188
rect 34244 13132 34254 13188
rect 34402 13132 34412 13188
rect 34468 13132 34478 13188
rect 35746 13132 35756 13188
rect 35812 13132 35822 13188
rect 3490 13020 3500 13076
rect 3556 13020 4060 13076
rect 4116 13020 7084 13076
rect 7140 13020 8204 13076
rect 8260 13020 10668 13076
rect 10724 13020 10734 13076
rect 11442 13020 11452 13076
rect 11508 13020 12236 13076
rect 12292 13020 12302 13076
rect 16370 13020 16380 13076
rect 16436 13020 18508 13076
rect 18564 13020 18574 13076
rect 18722 13020 18732 13076
rect 18788 13020 20748 13076
rect 20804 13020 21644 13076
rect 21700 13020 21710 13076
rect 25228 13020 25452 13076
rect 25508 13020 25518 13076
rect 25228 12964 25284 13020
rect 3332 12908 9100 12964
rect 9156 12908 9166 12964
rect 9650 12908 9660 12964
rect 9716 12908 9996 12964
rect 10052 12908 10332 12964
rect 10388 12908 10398 12964
rect 18050 12908 18060 12964
rect 18116 12908 20412 12964
rect 20468 12908 20478 12964
rect 23398 12908 23436 12964
rect 23492 12908 23502 12964
rect 25218 12908 25228 12964
rect 25284 12908 25294 12964
rect 3332 12516 3388 12908
rect 26852 12852 26908 13132
rect 34412 13076 34468 13132
rect 28130 13020 28140 13076
rect 28196 13020 29932 13076
rect 29988 13020 29998 13076
rect 33506 13020 33516 13076
rect 33572 13020 34468 13076
rect 34412 12964 34468 13020
rect 33394 12908 33404 12964
rect 33460 12908 34188 12964
rect 34244 12908 34254 12964
rect 34412 12908 35084 12964
rect 35140 12908 35150 12964
rect 35756 12852 35812 13132
rect 35970 13020 35980 13076
rect 36036 13020 39004 13076
rect 39060 13020 39070 13076
rect 39778 13020 39788 13076
rect 39844 13020 40684 13076
rect 40740 13020 40750 13076
rect 41682 13020 41692 13076
rect 41748 13020 43148 13076
rect 43204 13020 43214 13076
rect 38332 12908 40460 12964
rect 40516 12908 40526 12964
rect 42802 12908 42812 12964
rect 42868 12908 43820 12964
rect 43876 12908 43886 12964
rect 38332 12852 38388 12908
rect 7522 12796 7532 12852
rect 7588 12796 10668 12852
rect 10724 12796 10734 12852
rect 12562 12796 12572 12852
rect 12628 12796 13468 12852
rect 13524 12796 13534 12852
rect 14578 12796 14588 12852
rect 14644 12796 15148 12852
rect 15204 12796 15214 12852
rect 17154 12796 17164 12852
rect 17220 12796 19292 12852
rect 19348 12796 19358 12852
rect 21746 12796 21756 12852
rect 21812 12796 22428 12852
rect 22484 12796 22494 12852
rect 26852 12796 35812 12852
rect 38322 12796 38332 12852
rect 38388 12796 38398 12852
rect 38518 12796 38556 12852
rect 38612 12796 38622 12852
rect 43026 12796 43036 12852
rect 43092 12796 47852 12852
rect 47908 12796 47918 12852
rect 17164 12740 17220 12796
rect 4162 12684 4172 12740
rect 4228 12684 7532 12740
rect 7588 12684 7598 12740
rect 7970 12684 7980 12740
rect 8036 12684 8316 12740
rect 8372 12684 8382 12740
rect 10546 12684 10556 12740
rect 10612 12684 11788 12740
rect 11844 12684 11854 12740
rect 12226 12684 12236 12740
rect 12292 12684 17220 12740
rect 17724 12684 18620 12740
rect 18676 12684 18686 12740
rect 21634 12684 21644 12740
rect 21700 12684 34076 12740
rect 34132 12684 34748 12740
rect 34804 12684 34814 12740
rect 34972 12684 37100 12740
rect 37156 12684 37166 12740
rect 17724 12628 17780 12684
rect 34972 12628 35028 12684
rect 49200 12628 50000 12656
rect 4834 12572 4844 12628
rect 4900 12572 7644 12628
rect 7700 12572 7710 12628
rect 11890 12572 11900 12628
rect 11956 12572 13916 12628
rect 13972 12572 13982 12628
rect 16818 12572 16828 12628
rect 16884 12572 17780 12628
rect 18162 12572 18172 12628
rect 18228 12572 18238 12628
rect 20738 12572 20748 12628
rect 20804 12572 23100 12628
rect 23156 12572 23166 12628
rect 25554 12572 25564 12628
rect 25620 12572 26796 12628
rect 26852 12572 26862 12628
rect 33170 12572 33180 12628
rect 33236 12572 35028 12628
rect 36306 12572 36316 12628
rect 36372 12572 40348 12628
rect 40404 12572 41468 12628
rect 41524 12572 41534 12628
rect 46274 12572 46284 12628
rect 46340 12572 46900 12628
rect 47618 12572 47628 12628
rect 47684 12572 48188 12628
rect 48244 12572 50000 12628
rect 18172 12516 18228 12572
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 46844 12516 46900 12572
rect 49200 12544 50000 12572
rect 1922 12460 1932 12516
rect 1988 12460 3388 12516
rect 5730 12460 5740 12516
rect 5796 12460 6188 12516
rect 6244 12460 6254 12516
rect 7074 12460 7084 12516
rect 7140 12460 9548 12516
rect 9604 12460 13636 12516
rect 13794 12460 13804 12516
rect 13860 12460 13898 12516
rect 14364 12460 16716 12516
rect 16772 12460 16782 12516
rect 18172 12460 19628 12516
rect 19684 12460 19694 12516
rect 28690 12460 28700 12516
rect 28756 12460 32060 12516
rect 32116 12460 33068 12516
rect 33124 12460 33134 12516
rect 34850 12460 34860 12516
rect 34916 12460 36988 12516
rect 37044 12460 37054 12516
rect 46834 12460 46844 12516
rect 46900 12460 46910 12516
rect 13580 12404 13636 12460
rect 14364 12404 14420 12460
rect 6738 12348 6748 12404
rect 6804 12348 7420 12404
rect 7476 12348 7486 12404
rect 8082 12348 8092 12404
rect 8148 12348 10108 12404
rect 10164 12348 10174 12404
rect 11666 12348 11676 12404
rect 11732 12348 13356 12404
rect 13412 12348 13422 12404
rect 13580 12348 14420 12404
rect 14550 12348 14588 12404
rect 14644 12348 14654 12404
rect 15026 12348 15036 12404
rect 15092 12292 15148 12404
rect 15922 12348 15932 12404
rect 15988 12348 16268 12404
rect 16324 12348 18508 12404
rect 18564 12348 19964 12404
rect 20020 12348 20030 12404
rect 25302 12348 25340 12404
rect 25396 12348 25406 12404
rect 26338 12348 26348 12404
rect 26404 12348 28476 12404
rect 28532 12348 29372 12404
rect 29428 12348 29438 12404
rect 31126 12348 31164 12404
rect 31220 12348 31230 12404
rect 34402 12348 34412 12404
rect 34468 12348 36204 12404
rect 36260 12348 36270 12404
rect 36642 12348 36652 12404
rect 36708 12348 39004 12404
rect 39060 12348 39070 12404
rect 44146 12348 44156 12404
rect 44212 12348 44940 12404
rect 44996 12348 45276 12404
rect 45332 12348 45342 12404
rect 36204 12292 36260 12348
rect 3826 12236 3836 12292
rect 3892 12236 6188 12292
rect 6244 12236 6254 12292
rect 7298 12236 7308 12292
rect 7364 12236 8652 12292
rect 8708 12236 8718 12292
rect 10546 12236 10556 12292
rect 10612 12236 14476 12292
rect 14532 12236 14542 12292
rect 15092 12236 15372 12292
rect 15428 12236 15438 12292
rect 15698 12236 15708 12292
rect 15764 12236 16380 12292
rect 16436 12236 16446 12292
rect 19394 12236 19404 12292
rect 19460 12236 24108 12292
rect 24164 12236 24174 12292
rect 26002 12236 26012 12292
rect 26068 12236 27020 12292
rect 27076 12236 27468 12292
rect 27524 12236 29036 12292
rect 29092 12236 29820 12292
rect 29876 12236 29886 12292
rect 31266 12236 31276 12292
rect 31332 12236 31836 12292
rect 31892 12236 31902 12292
rect 34636 12236 35812 12292
rect 36204 12236 37100 12292
rect 37156 12236 37166 12292
rect 34636 12180 34692 12236
rect 35756 12180 35812 12236
rect 3042 12124 3052 12180
rect 3108 12124 3948 12180
rect 4004 12124 4014 12180
rect 6402 12124 6412 12180
rect 6468 12124 7868 12180
rect 7924 12124 7934 12180
rect 9090 12124 9100 12180
rect 9156 12124 10220 12180
rect 10276 12124 10286 12180
rect 10882 12124 10892 12180
rect 10948 12124 12348 12180
rect 12404 12124 13468 12180
rect 13524 12124 14028 12180
rect 14084 12124 14094 12180
rect 14354 12124 14364 12180
rect 14420 12124 14812 12180
rect 14868 12124 14878 12180
rect 17602 12124 17612 12180
rect 17668 12124 18620 12180
rect 18676 12124 18686 12180
rect 19030 12124 19068 12180
rect 19124 12124 19134 12180
rect 20962 12124 20972 12180
rect 21028 12124 25116 12180
rect 25172 12124 25182 12180
rect 26114 12124 26124 12180
rect 26180 12124 27580 12180
rect 27636 12124 27646 12180
rect 28130 12124 28140 12180
rect 28196 12124 29484 12180
rect 29540 12124 29550 12180
rect 30146 12124 30156 12180
rect 30212 12124 34692 12180
rect 34850 12124 34860 12180
rect 34916 12124 35532 12180
rect 35588 12124 35598 12180
rect 35756 12124 36316 12180
rect 36372 12124 36382 12180
rect 46722 12124 46732 12180
rect 46788 12124 47852 12180
rect 47908 12124 47918 12180
rect 20972 12068 21028 12124
rect 2818 12012 2828 12068
rect 2884 12012 8820 12068
rect 8978 12012 8988 12068
rect 9044 12012 9884 12068
rect 9940 12012 17164 12068
rect 17220 12012 17230 12068
rect 18050 12012 18060 12068
rect 18116 12012 21028 12068
rect 24210 12012 24220 12068
rect 24276 12012 26348 12068
rect 26404 12012 26414 12068
rect 31042 12012 31052 12068
rect 31108 12012 31612 12068
rect 31668 12012 31678 12068
rect 34962 12012 34972 12068
rect 35028 12012 35644 12068
rect 35700 12012 36876 12068
rect 36932 12012 36942 12068
rect 41122 12012 41132 12068
rect 41188 12012 42364 12068
rect 42420 12012 42430 12068
rect 45938 12012 45948 12068
rect 46004 12012 47516 12068
rect 47572 12012 48188 12068
rect 48244 12012 48254 12068
rect 8764 11956 8820 12012
rect 5954 11900 5964 11956
rect 6020 11900 7196 11956
rect 7252 11900 7532 11956
rect 7588 11900 7598 11956
rect 8764 11900 11228 11956
rect 11284 11900 11294 11956
rect 11778 11900 11788 11956
rect 11844 11900 13020 11956
rect 13076 11900 13086 11956
rect 15026 11900 15036 11956
rect 15092 11900 17612 11956
rect 17668 11900 18508 11956
rect 18564 11900 18574 11956
rect 18834 11900 18844 11956
rect 18900 11900 18956 11956
rect 19012 11900 19022 11956
rect 19618 11900 19628 11956
rect 19684 11900 26460 11956
rect 26516 11900 26526 11956
rect 34850 11900 34860 11956
rect 34916 11900 35868 11956
rect 35924 11900 35934 11956
rect 2258 11788 2268 11844
rect 2324 11788 3052 11844
rect 3108 11788 3118 11844
rect 8428 11788 9660 11844
rect 9716 11788 9726 11844
rect 10210 11788 10220 11844
rect 10276 11788 10314 11844
rect 11442 11788 11452 11844
rect 11508 11788 13132 11844
rect 13188 11788 13198 11844
rect 16930 11788 16940 11844
rect 16996 11788 18060 11844
rect 18116 11788 18126 11844
rect 18274 11788 18284 11844
rect 18340 11788 18396 11844
rect 18452 11788 18462 11844
rect 20850 11788 20860 11844
rect 20916 11788 21532 11844
rect 21588 11788 21598 11844
rect 21970 11788 21980 11844
rect 22036 11788 23660 11844
rect 23716 11788 24668 11844
rect 24724 11788 24734 11844
rect 27906 11788 27916 11844
rect 27972 11788 29260 11844
rect 29316 11788 29708 11844
rect 29764 11788 29774 11844
rect 30034 11788 30044 11844
rect 30100 11788 30492 11844
rect 30548 11788 30828 11844
rect 30884 11788 30894 11844
rect 33170 11788 33180 11844
rect 33236 11788 33740 11844
rect 33796 11788 33806 11844
rect 36978 11788 36988 11844
rect 37044 11788 38332 11844
rect 38388 11788 38398 11844
rect 43474 11788 43484 11844
rect 43540 11788 44380 11844
rect 44436 11788 44446 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 8428 11732 8484 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 6850 11676 6860 11732
rect 6916 11676 7196 11732
rect 7252 11676 7262 11732
rect 7858 11676 7868 11732
rect 7924 11676 8484 11732
rect 10546 11676 10556 11732
rect 10612 11676 12236 11732
rect 12292 11676 12302 11732
rect 13010 11676 13020 11732
rect 13076 11676 13804 11732
rect 13860 11676 13870 11732
rect 14354 11676 14364 11732
rect 14420 11676 15036 11732
rect 15092 11676 15102 11732
rect 16482 11676 16492 11732
rect 16548 11676 21308 11732
rect 21364 11676 21374 11732
rect 22306 11676 22316 11732
rect 22372 11676 23436 11732
rect 23492 11676 23502 11732
rect 34626 11676 34636 11732
rect 34692 11676 34702 11732
rect 35532 11676 40572 11732
rect 40628 11676 41132 11732
rect 41188 11676 41198 11732
rect 34636 11620 34692 11676
rect 35532 11620 35588 11676
rect 5058 11564 5068 11620
rect 5124 11564 6972 11620
rect 7028 11564 7038 11620
rect 12114 11564 12124 11620
rect 12180 11564 13412 11620
rect 14578 11564 14588 11620
rect 14644 11564 18396 11620
rect 18452 11564 18462 11620
rect 20290 11564 20300 11620
rect 20356 11564 21420 11620
rect 21476 11564 21486 11620
rect 22642 11564 22652 11620
rect 22708 11564 23100 11620
rect 23156 11564 23166 11620
rect 23538 11564 23548 11620
rect 23604 11564 23996 11620
rect 24052 11564 26908 11620
rect 31378 11564 31388 11620
rect 31444 11564 34076 11620
rect 34132 11564 34142 11620
rect 34636 11564 35588 11620
rect 36530 11564 36540 11620
rect 36596 11564 37436 11620
rect 37492 11564 37502 11620
rect 45714 11564 45724 11620
rect 45780 11564 46396 11620
rect 46452 11564 46462 11620
rect 13356 11508 13412 11564
rect 26852 11508 26908 11564
rect 3490 11452 3500 11508
rect 3556 11452 12460 11508
rect 12516 11452 12526 11508
rect 13346 11452 13356 11508
rect 13412 11452 13422 11508
rect 13580 11452 15148 11508
rect 15250 11452 15260 11508
rect 15316 11452 15354 11508
rect 17938 11452 17948 11508
rect 18004 11452 18284 11508
rect 18340 11452 18350 11508
rect 20626 11452 20636 11508
rect 20692 11452 21644 11508
rect 21700 11452 24780 11508
rect 24836 11452 24846 11508
rect 26852 11452 33460 11508
rect 33618 11452 33628 11508
rect 33684 11452 34748 11508
rect 34804 11452 35868 11508
rect 35924 11452 35934 11508
rect 36866 11452 36876 11508
rect 36932 11452 37548 11508
rect 37604 11452 37614 11508
rect 41458 11452 41468 11508
rect 41524 11452 42364 11508
rect 42420 11452 43036 11508
rect 43092 11452 43102 11508
rect 43474 11452 43484 11508
rect 43540 11452 48300 11508
rect 48356 11452 48366 11508
rect 13580 11396 13636 11452
rect 6290 11340 6300 11396
rect 6356 11340 6748 11396
rect 6804 11340 6814 11396
rect 8082 11340 8092 11396
rect 8148 11340 8988 11396
rect 9044 11340 9054 11396
rect 10658 11340 10668 11396
rect 10724 11340 11116 11396
rect 11172 11340 11182 11396
rect 11330 11340 11340 11396
rect 11396 11340 11900 11396
rect 11956 11340 13636 11396
rect 15092 11396 15148 11452
rect 33404 11396 33460 11452
rect 43484 11396 43540 11452
rect 15092 11340 23324 11396
rect 23380 11340 29708 11396
rect 29764 11340 29774 11396
rect 30818 11340 30828 11396
rect 30884 11340 31948 11396
rect 32004 11340 32172 11396
rect 32228 11340 32238 11396
rect 33404 11340 34076 11396
rect 34132 11340 34142 11396
rect 34514 11340 34524 11396
rect 34580 11340 35084 11396
rect 35140 11340 35150 11396
rect 35522 11340 35532 11396
rect 35588 11340 35980 11396
rect 36036 11340 36046 11396
rect 37090 11340 37100 11396
rect 37156 11340 37996 11396
rect 38052 11340 40236 11396
rect 40292 11340 41132 11396
rect 41188 11340 42028 11396
rect 42084 11340 43540 11396
rect 45154 11340 45164 11396
rect 45220 11340 46508 11396
rect 46564 11340 47628 11396
rect 47684 11340 47694 11396
rect 8642 11228 8652 11284
rect 8708 11228 10556 11284
rect 10612 11228 10622 11284
rect 11218 11228 11228 11284
rect 11284 11228 12012 11284
rect 12068 11228 12078 11284
rect 14476 11228 14812 11284
rect 14868 11228 16828 11284
rect 16884 11228 16894 11284
rect 17154 11228 17164 11284
rect 17220 11228 25340 11284
rect 25396 11228 25406 11284
rect 4498 11116 4508 11172
rect 4564 11116 5852 11172
rect 5908 11116 5918 11172
rect 6934 11116 6972 11172
rect 7028 11116 7038 11172
rect 8866 11116 8876 11172
rect 8932 11116 11788 11172
rect 11844 11116 11854 11172
rect 14476 11060 14532 11228
rect 29708 11172 29764 11340
rect 33730 11228 33740 11284
rect 33796 11228 34188 11284
rect 34244 11228 41020 11284
rect 41076 11228 41086 11284
rect 44930 11228 44940 11284
rect 44996 11228 45276 11284
rect 45332 11228 46396 11284
rect 46452 11228 46462 11284
rect 46834 11228 46844 11284
rect 46900 11228 47012 11284
rect 15092 11116 21476 11172
rect 22306 11116 22316 11172
rect 22372 11116 23548 11172
rect 23604 11116 23614 11172
rect 27766 11116 27804 11172
rect 27860 11116 28140 11172
rect 28196 11116 28206 11172
rect 29708 11116 34748 11172
rect 34804 11116 34814 11172
rect 45154 11116 45164 11172
rect 45220 11116 46060 11172
rect 46116 11116 46126 11172
rect 6066 11004 6076 11060
rect 6132 11004 14252 11060
rect 14308 11004 14318 11060
rect 14466 11004 14476 11060
rect 14532 11004 14542 11060
rect 14774 11004 14812 11060
rect 14868 11004 14878 11060
rect 15092 10948 15148 11116
rect 21420 11060 21476 11116
rect 22316 11060 22372 11116
rect 34748 11060 34804 11116
rect 46956 11060 47012 11228
rect 21046 11004 21084 11060
rect 21140 11004 21150 11060
rect 21420 11004 22372 11060
rect 34402 11004 34412 11060
rect 34468 11004 34524 11060
rect 34580 11004 34590 11060
rect 34748 11004 36092 11060
rect 36148 11004 38444 11060
rect 38500 11004 38510 11060
rect 44258 11004 44268 11060
rect 44324 11004 44828 11060
rect 44884 11004 47012 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 3042 10892 3052 10948
rect 3108 10892 11452 10948
rect 11508 10892 11518 10948
rect 12450 10892 12460 10948
rect 12516 10892 13356 10948
rect 13412 10892 15148 10948
rect 18610 10892 18620 10948
rect 18676 10892 19516 10948
rect 19572 10892 19582 10948
rect 20188 10892 20748 10948
rect 20804 10892 20814 10948
rect 21186 10892 21196 10948
rect 21252 10892 21420 10948
rect 21476 10892 21486 10948
rect 34066 10892 34076 10948
rect 34132 10892 34860 10948
rect 34916 10892 34926 10948
rect 20188 10836 20244 10892
rect 2930 10780 2940 10836
rect 2996 10780 7196 10836
rect 7252 10780 7262 10836
rect 14018 10780 14028 10836
rect 14084 10780 14588 10836
rect 14644 10780 14654 10836
rect 16258 10780 16268 10836
rect 16324 10780 17276 10836
rect 17332 10780 17724 10836
rect 17780 10780 17790 10836
rect 18732 10780 20244 10836
rect 20402 10780 20412 10836
rect 20468 10780 23884 10836
rect 23940 10780 23950 10836
rect 27346 10780 27356 10836
rect 27412 10780 28140 10836
rect 28196 10780 29260 10836
rect 29316 10780 30940 10836
rect 30996 10780 31006 10836
rect 18732 10724 18788 10780
rect 5618 10668 5628 10724
rect 5684 10668 6972 10724
rect 7028 10668 7038 10724
rect 12674 10668 12684 10724
rect 12740 10668 13580 10724
rect 13636 10668 13646 10724
rect 14242 10668 14252 10724
rect 14308 10668 18788 10724
rect 18918 10668 18956 10724
rect 19012 10668 19460 10724
rect 20738 10668 20748 10724
rect 20804 10668 21868 10724
rect 21924 10668 21934 10724
rect 23762 10668 23772 10724
rect 23828 10668 26348 10724
rect 26404 10668 30156 10724
rect 30212 10668 30222 10724
rect 33282 10668 33292 10724
rect 33348 10668 35308 10724
rect 35364 10668 36204 10724
rect 36260 10668 36270 10724
rect 43138 10668 43148 10724
rect 43204 10668 45500 10724
rect 45556 10668 45566 10724
rect 15260 10612 15316 10668
rect 6188 10556 11340 10612
rect 11396 10556 11406 10612
rect 12562 10556 12572 10612
rect 12628 10556 14476 10612
rect 14532 10556 14542 10612
rect 15250 10556 15260 10612
rect 15316 10556 15326 10612
rect 15586 10556 15596 10612
rect 15652 10556 16380 10612
rect 16436 10556 16446 10612
rect 17826 10556 17836 10612
rect 17892 10556 19180 10612
rect 19236 10556 19246 10612
rect 6188 10500 6244 10556
rect 19404 10500 19460 10668
rect 46956 10612 47012 11004
rect 21074 10556 21084 10612
rect 21140 10556 22988 10612
rect 23044 10556 23054 10612
rect 30818 10556 30828 10612
rect 30884 10556 32060 10612
rect 32116 10556 40012 10612
rect 40068 10556 40078 10612
rect 46946 10556 46956 10612
rect 47012 10556 47022 10612
rect 2146 10444 2156 10500
rect 2212 10444 6188 10500
rect 6244 10444 6254 10500
rect 9090 10444 9100 10500
rect 9156 10444 9166 10500
rect 12870 10444 12908 10500
rect 12964 10444 12974 10500
rect 13458 10444 13468 10500
rect 13524 10444 13804 10500
rect 13860 10444 15260 10500
rect 15316 10444 15326 10500
rect 19404 10444 24892 10500
rect 24948 10444 25228 10500
rect 25284 10444 25294 10500
rect 30034 10444 30044 10500
rect 30100 10444 30716 10500
rect 30772 10444 30782 10500
rect 30930 10444 30940 10500
rect 30996 10444 31948 10500
rect 32004 10444 32172 10500
rect 32228 10444 32508 10500
rect 32564 10444 33628 10500
rect 33684 10444 35756 10500
rect 35812 10444 36428 10500
rect 36484 10444 36494 10500
rect 39218 10444 39228 10500
rect 39284 10444 39676 10500
rect 39732 10444 40908 10500
rect 40964 10444 40974 10500
rect 9100 10276 9156 10444
rect 21186 10332 21196 10388
rect 21252 10332 21980 10388
rect 22036 10332 22046 10388
rect 23510 10332 23548 10388
rect 23604 10332 27244 10388
rect 27300 10332 27804 10388
rect 27860 10332 27870 10388
rect 29586 10332 29596 10388
rect 29652 10332 30156 10388
rect 30212 10332 35644 10388
rect 35700 10332 35710 10388
rect 35858 10332 35868 10388
rect 35924 10332 37772 10388
rect 37828 10332 37838 10388
rect 5282 10220 5292 10276
rect 5348 10220 6636 10276
rect 6692 10220 6702 10276
rect 9100 10220 15372 10276
rect 15428 10220 15438 10276
rect 20962 10220 20972 10276
rect 21028 10220 22092 10276
rect 22148 10220 23212 10276
rect 23268 10220 23278 10276
rect 29362 10220 29372 10276
rect 29428 10220 33180 10276
rect 33236 10220 33246 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 21644 10164 21700 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 6962 10108 6972 10164
rect 7028 10108 7308 10164
rect 7364 10108 18956 10164
rect 19012 10108 19022 10164
rect 21634 10108 21644 10164
rect 21700 10108 21710 10164
rect 23314 10108 23324 10164
rect 23380 10108 23996 10164
rect 24052 10108 24062 10164
rect 33282 10108 33292 10164
rect 33348 10108 34300 10164
rect 34356 10108 34366 10164
rect 36530 10108 36540 10164
rect 36596 10108 36988 10164
rect 37044 10108 37660 10164
rect 37716 10108 38556 10164
rect 38612 10108 38622 10164
rect 8754 9996 8764 10052
rect 8820 9996 9772 10052
rect 9828 9996 12908 10052
rect 12964 9996 12974 10052
rect 15922 9996 15932 10052
rect 15988 9996 19852 10052
rect 19908 9996 19918 10052
rect 27122 9996 27132 10052
rect 27188 9996 27804 10052
rect 27860 9996 37212 10052
rect 37268 9996 37278 10052
rect 41682 9996 41692 10052
rect 41748 9996 42476 10052
rect 42532 9996 42812 10052
rect 42868 9996 42878 10052
rect 7634 9884 7644 9940
rect 7700 9884 8092 9940
rect 8148 9884 8158 9940
rect 10070 9884 10108 9940
rect 10164 9884 10174 9940
rect 12002 9884 12012 9940
rect 12068 9884 12078 9940
rect 15092 9884 16044 9940
rect 16100 9884 16110 9940
rect 16370 9884 16380 9940
rect 16436 9884 18732 9940
rect 18788 9884 18798 9940
rect 21046 9884 21084 9940
rect 21140 9884 21150 9940
rect 35298 9884 35308 9940
rect 35364 9884 40124 9940
rect 40180 9884 40190 9940
rect 12012 9828 12068 9884
rect 15092 9828 15148 9884
rect 3826 9772 3836 9828
rect 3892 9772 10332 9828
rect 10388 9772 10398 9828
rect 12012 9772 15148 9828
rect 15698 9772 15708 9828
rect 15764 9772 16268 9828
rect 16324 9772 17724 9828
rect 17780 9772 18620 9828
rect 18676 9772 19404 9828
rect 19460 9772 24332 9828
rect 24388 9772 24398 9828
rect 24882 9772 24892 9828
rect 24948 9772 28588 9828
rect 28644 9772 28654 9828
rect 30604 9772 36092 9828
rect 36148 9772 37996 9828
rect 38052 9772 38062 9828
rect 40338 9772 40348 9828
rect 40404 9772 41916 9828
rect 41972 9772 43036 9828
rect 43092 9772 43102 9828
rect 30604 9716 30660 9772
rect 2034 9660 2044 9716
rect 2100 9660 5964 9716
rect 6020 9660 6030 9716
rect 7858 9660 7868 9716
rect 7924 9660 9660 9716
rect 9716 9660 9726 9716
rect 14802 9660 14812 9716
rect 14868 9660 15148 9716
rect 15204 9660 20748 9716
rect 20804 9660 20814 9716
rect 23090 9660 23100 9716
rect 23156 9660 23436 9716
rect 23492 9660 23502 9716
rect 28242 9660 28252 9716
rect 28308 9660 30660 9716
rect 30818 9660 30828 9716
rect 30884 9660 33180 9716
rect 33236 9660 33246 9716
rect 34178 9660 34188 9716
rect 34244 9660 36652 9716
rect 36708 9660 36718 9716
rect 38658 9660 38668 9716
rect 38724 9660 41020 9716
rect 41076 9660 41086 9716
rect 3378 9548 3388 9604
rect 3444 9548 8428 9604
rect 8484 9548 8494 9604
rect 10294 9548 10332 9604
rect 10388 9548 10398 9604
rect 17714 9548 17724 9604
rect 17780 9548 18172 9604
rect 18228 9548 22428 9604
rect 22484 9548 22494 9604
rect 28466 9548 28476 9604
rect 28532 9548 31164 9604
rect 31220 9548 31230 9604
rect 36418 9548 36428 9604
rect 36484 9548 37212 9604
rect 37268 9548 37278 9604
rect 44482 9548 44492 9604
rect 44548 9548 44940 9604
rect 44996 9548 45006 9604
rect 5058 9436 5068 9492
rect 5124 9436 5516 9492
rect 5572 9436 6020 9492
rect 7522 9436 7532 9492
rect 7588 9436 8316 9492
rect 8372 9436 8382 9492
rect 9314 9436 9324 9492
rect 9380 9436 11004 9492
rect 11060 9436 11070 9492
rect 30258 9436 30268 9492
rect 30324 9436 37772 9492
rect 37828 9436 37838 9492
rect 5964 9380 6020 9436
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 3378 9324 3388 9380
rect 3444 9324 4172 9380
rect 4228 9324 5740 9380
rect 5796 9324 5806 9380
rect 5964 9324 19404 9380
rect 19460 9324 19470 9380
rect 25554 9324 25564 9380
rect 25620 9324 29372 9380
rect 29428 9324 29438 9380
rect 2930 9212 2940 9268
rect 2996 9212 4060 9268
rect 4116 9212 4126 9268
rect 5506 9212 5516 9268
rect 5572 9212 6412 9268
rect 6468 9212 6972 9268
rect 7028 9212 14700 9268
rect 14756 9212 14766 9268
rect 16790 9212 16828 9268
rect 16884 9212 18284 9268
rect 18340 9212 18350 9268
rect 20290 9212 20300 9268
rect 20356 9212 25676 9268
rect 25732 9212 26012 9268
rect 26068 9212 26078 9268
rect 26450 9212 26460 9268
rect 26516 9212 26526 9268
rect 29474 9212 29484 9268
rect 29540 9212 30604 9268
rect 30660 9212 30670 9268
rect 35634 9212 35644 9268
rect 35700 9212 37100 9268
rect 37156 9212 37166 9268
rect 39330 9212 39340 9268
rect 39396 9212 39900 9268
rect 39956 9212 43484 9268
rect 43540 9212 43550 9268
rect 4274 9100 4284 9156
rect 4340 9100 13356 9156
rect 13412 9100 13422 9156
rect 20626 9100 20636 9156
rect 20692 9100 22092 9156
rect 22148 9100 22158 9156
rect 2034 8988 2044 9044
rect 2100 8988 5404 9044
rect 5460 8988 5470 9044
rect 6514 8988 6524 9044
rect 6580 8988 7196 9044
rect 7252 8988 7980 9044
rect 8036 8988 8046 9044
rect 11218 8988 11228 9044
rect 11284 8988 11788 9044
rect 14690 8988 14700 9044
rect 14756 8988 15260 9044
rect 15316 8988 15326 9044
rect 21410 8988 21420 9044
rect 21476 8988 22204 9044
rect 22260 8988 22270 9044
rect 4946 8876 4956 8932
rect 5012 8876 7868 8932
rect 7924 8876 7934 8932
rect 11732 8820 11788 8988
rect 26012 8932 26068 9212
rect 26460 9156 26516 9212
rect 26460 9100 26796 9156
rect 26852 9100 29148 9156
rect 29204 9100 29820 9156
rect 29876 9100 29886 9156
rect 31154 9100 31164 9156
rect 31220 9100 31948 9156
rect 32004 9100 32014 9156
rect 40450 9100 40460 9156
rect 40516 9100 43260 9156
rect 43316 9100 43326 9156
rect 29586 8988 29596 9044
rect 29652 8988 30828 9044
rect 30884 8988 30894 9044
rect 31826 8988 31836 9044
rect 31892 8988 35308 9044
rect 35364 8988 35374 9044
rect 36082 8988 36092 9044
rect 36148 8988 37212 9044
rect 37268 8988 37278 9044
rect 38612 8988 47852 9044
rect 47908 8988 47918 9044
rect 12898 8876 12908 8932
rect 12964 8876 14476 8932
rect 14532 8876 14542 8932
rect 19254 8876 19292 8932
rect 19348 8876 19358 8932
rect 19506 8876 19516 8932
rect 19572 8876 21868 8932
rect 21924 8876 21934 8932
rect 22092 8876 23436 8932
rect 23492 8876 23502 8932
rect 26012 8876 32788 8932
rect 34402 8876 34412 8932
rect 34468 8876 35420 8932
rect 35476 8876 35486 8932
rect 22092 8820 22148 8876
rect 32732 8820 32788 8876
rect 38612 8820 38668 8988
rect 42466 8876 42476 8932
rect 42532 8876 43820 8932
rect 43876 8876 43886 8932
rect 3266 8764 3276 8820
rect 3332 8764 5012 8820
rect 7410 8764 7420 8820
rect 7476 8764 8764 8820
rect 8820 8764 8830 8820
rect 11732 8764 13468 8820
rect 13524 8764 14028 8820
rect 14084 8764 22148 8820
rect 23314 8764 23324 8820
rect 23380 8764 28140 8820
rect 28196 8764 28206 8820
rect 32732 8764 38668 8820
rect 4956 8708 5012 8764
rect 4956 8652 7644 8708
rect 7700 8652 7710 8708
rect 7970 8652 7980 8708
rect 8036 8652 8876 8708
rect 8932 8652 8942 8708
rect 12674 8652 12684 8708
rect 12740 8652 13804 8708
rect 13860 8652 20860 8708
rect 20916 8652 22764 8708
rect 22820 8652 22830 8708
rect 22988 8652 26908 8708
rect 27010 8652 27020 8708
rect 27076 8652 27804 8708
rect 27860 8652 27870 8708
rect 35858 8652 35868 8708
rect 35924 8652 36316 8708
rect 36372 8652 36382 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 5516 8540 10220 8596
rect 10276 8540 10286 8596
rect 12786 8540 12796 8596
rect 12852 8540 13244 8596
rect 13300 8540 14924 8596
rect 14980 8540 14990 8596
rect 0 8372 800 8400
rect 0 8316 4060 8372
rect 4116 8316 4126 8372
rect 0 8288 800 8316
rect 5516 8260 5572 8540
rect 22988 8484 23044 8652
rect 26852 8596 26908 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 26852 8540 27636 8596
rect 37090 8540 37100 8596
rect 37156 8540 38332 8596
rect 38388 8540 42812 8596
rect 42868 8540 42878 8596
rect 6822 8428 6860 8484
rect 6916 8428 6926 8484
rect 12124 8428 13916 8484
rect 13972 8428 13982 8484
rect 14802 8428 14812 8484
rect 14868 8428 15148 8484
rect 15204 8428 15214 8484
rect 18610 8428 18620 8484
rect 18676 8428 21084 8484
rect 21140 8428 22988 8484
rect 23044 8428 23054 8484
rect 24658 8428 24668 8484
rect 24724 8428 26908 8484
rect 26964 8428 26974 8484
rect 12124 8372 12180 8428
rect 27580 8372 27636 8540
rect 35970 8428 35980 8484
rect 36036 8428 36074 8484
rect 37202 8428 37212 8484
rect 37268 8428 41356 8484
rect 41412 8428 41422 8484
rect 10770 8316 10780 8372
rect 10836 8316 11676 8372
rect 11732 8316 12012 8372
rect 12068 8316 12180 8372
rect 19170 8316 19180 8372
rect 19236 8316 19292 8372
rect 19348 8316 19358 8372
rect 19842 8316 19852 8372
rect 19908 8316 21532 8372
rect 21588 8316 21598 8372
rect 27570 8316 27580 8372
rect 27636 8316 28588 8372
rect 28644 8316 32620 8372
rect 32676 8316 32686 8372
rect 34738 8316 34748 8372
rect 34804 8316 37100 8372
rect 37156 8316 37166 8372
rect 37324 8316 38444 8372
rect 38500 8316 38510 8372
rect 40114 8316 40124 8372
rect 40180 8316 40796 8372
rect 40852 8316 42252 8372
rect 42308 8316 42318 8372
rect 47394 8316 47404 8372
rect 47460 8316 48188 8372
rect 48244 8316 48254 8372
rect 3714 8204 3724 8260
rect 3780 8204 5572 8260
rect 6290 8204 6300 8260
rect 6356 8204 8204 8260
rect 8260 8204 9100 8260
rect 9156 8204 9166 8260
rect 10098 8204 10108 8260
rect 10164 8204 13804 8260
rect 13860 8204 13870 8260
rect 15026 8204 15036 8260
rect 15092 8204 21196 8260
rect 21252 8204 21262 8260
rect 21410 8204 21420 8260
rect 21476 8204 23884 8260
rect 23940 8204 23950 8260
rect 25890 8204 25900 8260
rect 25956 8204 29708 8260
rect 29764 8204 29774 8260
rect 32274 8204 32284 8260
rect 32340 8204 33292 8260
rect 33348 8204 33358 8260
rect 34962 8204 34972 8260
rect 35028 8204 35532 8260
rect 35588 8204 36204 8260
rect 36260 8204 36270 8260
rect 37324 8148 37380 8316
rect 37762 8204 37772 8260
rect 37828 8204 37838 8260
rect 37986 8204 37996 8260
rect 38052 8204 41020 8260
rect 41076 8204 41086 8260
rect 41234 8204 41244 8260
rect 41300 8204 42140 8260
rect 42196 8204 42206 8260
rect 42802 8204 42812 8260
rect 42868 8204 44156 8260
rect 44212 8204 44222 8260
rect 44482 8204 44492 8260
rect 44548 8204 45388 8260
rect 45444 8204 45454 8260
rect 5730 8092 5740 8148
rect 5796 8092 8092 8148
rect 8148 8092 8158 8148
rect 8428 8092 10444 8148
rect 10500 8092 10510 8148
rect 12786 8092 12796 8148
rect 12852 8092 13468 8148
rect 13524 8092 13534 8148
rect 15586 8092 15596 8148
rect 15652 8092 16828 8148
rect 16884 8092 16894 8148
rect 17042 8092 17052 8148
rect 17108 8092 18844 8148
rect 18900 8092 18910 8148
rect 20402 8092 20412 8148
rect 20468 8092 21756 8148
rect 21812 8092 21822 8148
rect 23090 8092 23100 8148
rect 23156 8092 26348 8148
rect 26404 8092 26414 8148
rect 29586 8092 29596 8148
rect 29652 8092 30492 8148
rect 30548 8092 31276 8148
rect 31332 8092 31342 8148
rect 34178 8092 34188 8148
rect 34244 8092 35420 8148
rect 35476 8092 35486 8148
rect 35746 8092 35756 8148
rect 35812 8092 37100 8148
rect 37156 8092 37380 8148
rect 37772 8148 37828 8204
rect 37772 8092 40012 8148
rect 40068 8092 43148 8148
rect 43204 8092 43214 8148
rect 8428 8036 8484 8092
rect 2818 7980 2828 8036
rect 2884 7980 3388 8036
rect 6962 7980 6972 8036
rect 7028 7980 7532 8036
rect 7588 7980 7598 8036
rect 7858 7980 7868 8036
rect 7924 7980 8428 8036
rect 8484 7980 8494 8036
rect 10210 7980 10220 8036
rect 10276 7980 15148 8036
rect 15922 7980 15932 8036
rect 15988 7980 16940 8036
rect 16996 7980 17006 8036
rect 17826 7980 17836 8036
rect 17892 7980 18508 8036
rect 18564 7980 18574 8036
rect 18732 7980 21980 8036
rect 22036 7980 22046 8036
rect 26562 7980 26572 8036
rect 26628 7980 27132 8036
rect 27188 7980 28140 8036
rect 28196 7980 29148 8036
rect 29204 7980 29214 8036
rect 29362 7980 29372 8036
rect 29428 7980 30268 8036
rect 30324 7980 30334 8036
rect 34850 7980 34860 8036
rect 34916 7980 35196 8036
rect 35252 7980 35262 8036
rect 35522 7980 35532 8036
rect 35588 7980 35644 8036
rect 35700 7980 35710 8036
rect 37426 7980 37436 8036
rect 37492 7980 38668 8036
rect 38724 7980 39788 8036
rect 39844 7980 39854 8036
rect 40124 7980 40236 8036
rect 40292 7980 40852 8036
rect 41906 7980 41916 8036
rect 41972 7980 43260 8036
rect 43316 7980 43326 8036
rect 43810 7980 43820 8036
rect 43876 7980 44940 8036
rect 44996 7980 45006 8036
rect 3332 7924 3388 7980
rect 3332 7868 4620 7924
rect 4676 7868 7644 7924
rect 7700 7868 9436 7924
rect 9492 7868 9502 7924
rect 15092 7812 15148 7980
rect 18732 7924 18788 7980
rect 40124 7924 40180 7980
rect 16930 7868 16940 7924
rect 16996 7868 18788 7924
rect 21522 7868 21532 7924
rect 21588 7868 23212 7924
rect 23268 7868 33852 7924
rect 33908 7868 33918 7924
rect 34290 7868 34300 7924
rect 34356 7868 38556 7924
rect 38612 7868 39676 7924
rect 39732 7868 40180 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 40796 7812 40852 7980
rect 41010 7868 41020 7924
rect 41076 7868 42812 7924
rect 42868 7868 43372 7924
rect 43428 7868 43438 7924
rect 43820 7812 43876 7980
rect 6514 7756 6524 7812
rect 6580 7756 12908 7812
rect 12964 7756 12974 7812
rect 15092 7756 18620 7812
rect 18676 7756 18686 7812
rect 20290 7756 20300 7812
rect 20356 7756 20860 7812
rect 20916 7756 20926 7812
rect 21410 7756 21420 7812
rect 21476 7756 24220 7812
rect 24276 7756 24286 7812
rect 32274 7756 32284 7812
rect 32340 7756 33292 7812
rect 33348 7756 35084 7812
rect 35140 7756 35150 7812
rect 40796 7756 43876 7812
rect 49200 7700 50000 7728
rect 6850 7644 6860 7700
rect 6916 7644 7588 7700
rect 10322 7644 10332 7700
rect 10388 7644 10892 7700
rect 10948 7644 12348 7700
rect 12404 7644 12414 7700
rect 16902 7644 16940 7700
rect 16996 7644 17006 7700
rect 18834 7644 18844 7700
rect 18900 7644 19292 7700
rect 19348 7644 21644 7700
rect 21700 7644 21710 7700
rect 27794 7644 27804 7700
rect 27860 7644 29484 7700
rect 29540 7644 29550 7700
rect 30370 7644 30380 7700
rect 30436 7644 30940 7700
rect 30996 7644 31006 7700
rect 33730 7644 33740 7700
rect 33796 7644 34636 7700
rect 34692 7644 34702 7700
rect 35830 7644 35868 7700
rect 35924 7644 35934 7700
rect 38882 7644 38892 7700
rect 38948 7644 39228 7700
rect 39284 7644 39294 7700
rect 40226 7644 40236 7700
rect 40292 7644 40908 7700
rect 40964 7644 40974 7700
rect 41234 7644 41244 7700
rect 41300 7644 41580 7700
rect 41636 7644 41646 7700
rect 44146 7644 44156 7700
rect 44212 7644 45052 7700
rect 45108 7644 45118 7700
rect 48178 7644 48188 7700
rect 48244 7644 50000 7700
rect 4162 7532 4172 7588
rect 4228 7532 5628 7588
rect 5684 7532 5694 7588
rect 7532 7476 7588 7644
rect 49200 7616 50000 7644
rect 9762 7532 9772 7588
rect 9828 7532 10780 7588
rect 10836 7532 10846 7588
rect 13458 7532 13468 7588
rect 13524 7532 15820 7588
rect 15876 7532 15886 7588
rect 17490 7532 17500 7588
rect 17556 7532 18452 7588
rect 18582 7532 18620 7588
rect 18676 7532 18686 7588
rect 19058 7532 19068 7588
rect 19124 7532 21084 7588
rect 21140 7532 21150 7588
rect 21746 7532 21756 7588
rect 21812 7532 24220 7588
rect 24276 7532 25116 7588
rect 25172 7532 25182 7588
rect 25778 7532 25788 7588
rect 25844 7532 26348 7588
rect 26404 7532 33068 7588
rect 33124 7532 33134 7588
rect 36194 7532 36204 7588
rect 36260 7532 36764 7588
rect 36820 7532 36830 7588
rect 37202 7532 37212 7588
rect 37268 7532 39116 7588
rect 39172 7532 39182 7588
rect 40338 7532 40348 7588
rect 40404 7532 42476 7588
rect 42532 7532 42542 7588
rect 44454 7532 44492 7588
rect 44548 7532 44558 7588
rect 18396 7476 18452 7532
rect 6934 7420 6972 7476
rect 7028 7420 7038 7476
rect 7522 7420 7532 7476
rect 7588 7420 7598 7476
rect 9202 7420 9212 7476
rect 9268 7420 9996 7476
rect 10052 7420 10062 7476
rect 16706 7420 16716 7476
rect 16772 7420 17276 7476
rect 17332 7420 18172 7476
rect 18228 7420 18238 7476
rect 18396 7420 23604 7476
rect 24546 7420 24556 7476
rect 24612 7420 26460 7476
rect 26516 7420 30268 7476
rect 30324 7420 31276 7476
rect 31332 7420 31342 7476
rect 33842 7420 33852 7476
rect 33908 7420 37100 7476
rect 37156 7420 37166 7476
rect 38098 7420 38108 7476
rect 38164 7420 38668 7476
rect 38724 7420 38734 7476
rect 39778 7420 39788 7476
rect 39844 7420 41804 7476
rect 41860 7420 41870 7476
rect 43698 7420 43708 7476
rect 43764 7420 45276 7476
rect 45332 7420 46956 7476
rect 47012 7420 47516 7476
rect 47572 7420 47582 7476
rect 3154 7308 3164 7364
rect 3220 7308 8988 7364
rect 9044 7308 9054 7364
rect 10658 7308 10668 7364
rect 10724 7308 14252 7364
rect 14308 7308 15148 7364
rect 16258 7308 16268 7364
rect 16324 7308 17500 7364
rect 17556 7308 17566 7364
rect 18386 7308 18396 7364
rect 18452 7308 18508 7364
rect 18564 7308 18574 7364
rect 19740 7308 22764 7364
rect 22820 7308 23324 7364
rect 23380 7308 23390 7364
rect 15092 7252 15148 7308
rect 19740 7252 19796 7308
rect 23548 7252 23604 7420
rect 24994 7308 25004 7364
rect 25060 7308 26124 7364
rect 26180 7308 26348 7364
rect 26404 7308 26414 7364
rect 27430 7308 27468 7364
rect 27524 7308 27534 7364
rect 30370 7308 30380 7364
rect 30436 7308 32172 7364
rect 32228 7308 32238 7364
rect 32610 7308 32620 7364
rect 32676 7308 37884 7364
rect 37940 7308 37950 7364
rect 38322 7308 38332 7364
rect 38388 7308 38892 7364
rect 38948 7308 38958 7364
rect 15092 7196 19796 7252
rect 19954 7196 19964 7252
rect 20020 7196 20412 7252
rect 20468 7196 20478 7252
rect 21186 7196 21196 7252
rect 21252 7196 22204 7252
rect 22260 7196 22270 7252
rect 23548 7196 29596 7252
rect 29652 7196 29662 7252
rect 36418 7196 36428 7252
rect 36484 7196 36988 7252
rect 37044 7196 37772 7252
rect 37828 7196 38220 7252
rect 38276 7196 38286 7252
rect 11218 7084 11228 7140
rect 11284 7084 11294 7140
rect 18834 7084 18844 7140
rect 18900 7084 19852 7140
rect 19908 7084 19918 7140
rect 20962 7084 20972 7140
rect 21028 7084 21420 7140
rect 21476 7084 21486 7140
rect 40114 7084 40124 7140
rect 40180 7084 41244 7140
rect 41300 7084 41310 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 5954 6972 5964 7028
rect 6020 6972 7980 7028
rect 8036 6972 8046 7028
rect 5964 6916 6020 6972
rect 2706 6860 2716 6916
rect 2772 6860 6020 6916
rect 9090 6860 9100 6916
rect 9156 6860 9604 6916
rect 9548 6804 9604 6860
rect 11228 6804 11284 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 17714 6972 17724 7028
rect 17780 6972 18284 7028
rect 18340 6972 22372 7028
rect 24546 6972 24556 7028
rect 24612 6972 32732 7028
rect 32788 6972 32798 7028
rect 35606 6972 35644 7028
rect 35700 6972 35710 7028
rect 39330 6972 39340 7028
rect 39396 6972 41468 7028
rect 41524 6972 43260 7028
rect 43316 6972 43326 7028
rect 22316 6916 22372 6972
rect 16706 6860 16716 6916
rect 16772 6860 22092 6916
rect 22148 6860 22158 6916
rect 22316 6860 26908 6916
rect 26964 6860 27804 6916
rect 27860 6860 28364 6916
rect 28420 6860 28430 6916
rect 32274 6860 32284 6916
rect 32340 6860 33516 6916
rect 33572 6860 37212 6916
rect 37268 6860 37278 6916
rect 38098 6860 38108 6916
rect 38164 6860 38780 6916
rect 38836 6860 38846 6916
rect 6738 6748 6748 6804
rect 6804 6748 7868 6804
rect 7924 6748 9324 6804
rect 9380 6748 9390 6804
rect 9538 6748 9548 6804
rect 9604 6748 9614 6804
rect 9762 6748 9772 6804
rect 9828 6748 11452 6804
rect 11508 6748 11518 6804
rect 20178 6748 20188 6804
rect 20244 6748 21756 6804
rect 21812 6748 21822 6804
rect 27122 6748 27132 6804
rect 27188 6748 28812 6804
rect 28868 6748 28878 6804
rect 31714 6748 31724 6804
rect 31780 6748 32396 6804
rect 32452 6748 32462 6804
rect 32610 6748 32620 6804
rect 32676 6748 34860 6804
rect 34916 6748 34926 6804
rect 35970 6748 35980 6804
rect 36036 6748 36876 6804
rect 36932 6748 36942 6804
rect 37762 6748 37772 6804
rect 37828 6748 38892 6804
rect 38948 6748 40124 6804
rect 40180 6748 40190 6804
rect 3826 6636 3836 6692
rect 3892 6636 6860 6692
rect 6916 6636 6926 6692
rect 7410 6636 7420 6692
rect 7476 6636 9212 6692
rect 9268 6636 9278 6692
rect 9538 6636 9548 6692
rect 9604 6636 14140 6692
rect 14196 6636 15148 6692
rect 16370 6636 16380 6692
rect 16436 6636 17500 6692
rect 17556 6636 18060 6692
rect 18116 6636 19348 6692
rect 19506 6636 19516 6692
rect 19572 6636 20636 6692
rect 20692 6636 22316 6692
rect 22372 6636 22382 6692
rect 24882 6636 24892 6692
rect 24948 6636 26684 6692
rect 26740 6636 26750 6692
rect 27346 6636 27356 6692
rect 27412 6636 27468 6692
rect 27524 6636 27534 6692
rect 28018 6636 28028 6692
rect 28084 6636 29932 6692
rect 29988 6636 29998 6692
rect 30482 6636 30492 6692
rect 30548 6636 31500 6692
rect 31556 6636 33068 6692
rect 33124 6636 33134 6692
rect 36278 6636 36316 6692
rect 36372 6636 36382 6692
rect 46946 6636 46956 6692
rect 47012 6636 47852 6692
rect 47908 6636 47918 6692
rect 3378 6524 3388 6580
rect 3444 6524 3454 6580
rect 4274 6524 4284 6580
rect 4340 6524 5516 6580
rect 5572 6524 5582 6580
rect 5842 6524 5852 6580
rect 5908 6524 8988 6580
rect 9044 6524 9054 6580
rect 9650 6524 9660 6580
rect 9716 6524 11004 6580
rect 11060 6524 11070 6580
rect 12534 6524 12572 6580
rect 12628 6524 12638 6580
rect 3388 6468 3444 6524
rect 15092 6468 15148 6636
rect 19292 6580 19348 6636
rect 16706 6524 16716 6580
rect 16772 6524 18844 6580
rect 18900 6524 18910 6580
rect 19292 6524 23100 6580
rect 23156 6524 27916 6580
rect 27972 6524 27982 6580
rect 31266 6524 31276 6580
rect 31332 6524 33292 6580
rect 33348 6524 33358 6580
rect 35746 6524 35756 6580
rect 35812 6524 38556 6580
rect 38612 6524 39788 6580
rect 39844 6524 39854 6580
rect 42130 6524 42140 6580
rect 42196 6524 44940 6580
rect 44996 6524 45006 6580
rect 45154 6524 45164 6580
rect 45220 6524 46060 6580
rect 46116 6524 47180 6580
rect 47236 6524 47246 6580
rect 45164 6468 45220 6524
rect 3388 6412 6076 6468
rect 6132 6412 6142 6468
rect 6402 6412 6412 6468
rect 6468 6412 7084 6468
rect 7140 6412 7150 6468
rect 7410 6412 7420 6468
rect 7476 6412 8316 6468
rect 8372 6412 9324 6468
rect 9380 6412 9390 6468
rect 11218 6412 11228 6468
rect 11284 6412 13468 6468
rect 13524 6412 13916 6468
rect 13972 6412 13982 6468
rect 15092 6412 17724 6468
rect 17780 6412 17790 6468
rect 18610 6412 18620 6468
rect 18676 6412 26908 6468
rect 27794 6412 27804 6468
rect 27860 6412 29596 6468
rect 29652 6412 29662 6468
rect 33618 6412 33628 6468
rect 33684 6412 34300 6468
rect 34356 6412 35196 6468
rect 35252 6412 37436 6468
rect 37492 6412 37502 6468
rect 39554 6412 39564 6468
rect 39620 6412 40236 6468
rect 40292 6412 40302 6468
rect 41682 6412 41692 6468
rect 41748 6412 42476 6468
rect 42532 6412 42542 6468
rect 44370 6412 44380 6468
rect 44436 6412 45220 6468
rect 46162 6412 46172 6468
rect 46228 6412 47628 6468
rect 47684 6412 48188 6468
rect 48244 6412 48254 6468
rect 18620 6356 18676 6412
rect 8530 6300 8540 6356
rect 8596 6300 10108 6356
rect 10164 6300 10668 6356
rect 10724 6300 10734 6356
rect 14578 6300 14588 6356
rect 14644 6300 18676 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 26852 6244 26908 6412
rect 27010 6300 27020 6356
rect 27076 6300 27356 6356
rect 27412 6300 27422 6356
rect 29484 6300 30940 6356
rect 30996 6300 31006 6356
rect 34850 6300 34860 6356
rect 34916 6300 40908 6356
rect 40964 6300 40974 6356
rect 43698 6300 43708 6356
rect 43764 6300 45388 6356
rect 45444 6300 46620 6356
rect 46676 6300 47068 6356
rect 47124 6300 47134 6356
rect 29484 6244 29540 6300
rect 5170 6188 5180 6244
rect 5236 6188 13692 6244
rect 13748 6188 14364 6244
rect 14420 6188 14924 6244
rect 14980 6188 14990 6244
rect 26852 6188 29484 6244
rect 29540 6188 29550 6244
rect 30258 6188 30268 6244
rect 30324 6188 31948 6244
rect 32004 6188 32014 6244
rect 34738 6188 34748 6244
rect 34804 6188 35756 6244
rect 35812 6188 36204 6244
rect 36260 6188 36270 6244
rect 40338 6188 40348 6244
rect 40404 6188 42140 6244
rect 42196 6188 42206 6244
rect 6178 6076 6188 6132
rect 6244 6076 7084 6132
rect 7140 6076 8092 6132
rect 8148 6076 8158 6132
rect 8978 6076 8988 6132
rect 9044 6076 9772 6132
rect 9828 6076 10892 6132
rect 10948 6076 10958 6132
rect 12898 6076 12908 6132
rect 12964 6076 13468 6132
rect 13524 6076 14476 6132
rect 14532 6076 14542 6132
rect 16818 6076 16828 6132
rect 16884 6076 17500 6132
rect 17556 6076 17948 6132
rect 18004 6076 18014 6132
rect 19282 6076 19292 6132
rect 19348 6076 19964 6132
rect 20020 6076 20030 6132
rect 20738 6076 20748 6132
rect 20804 6076 22988 6132
rect 23044 6076 23054 6132
rect 24556 6076 26124 6132
rect 26180 6076 26190 6132
rect 26786 6076 26796 6132
rect 26852 6076 27356 6132
rect 27412 6076 27422 6132
rect 28354 6076 28364 6132
rect 28420 6076 30604 6132
rect 30660 6076 30670 6132
rect 34066 6076 34076 6132
rect 34132 6076 35980 6132
rect 36036 6076 36428 6132
rect 36484 6076 36494 6132
rect 37174 6076 37212 6132
rect 37268 6076 37278 6132
rect 24556 6020 24612 6076
rect 7746 5964 7756 6020
rect 7812 5964 8428 6020
rect 8484 5964 8494 6020
rect 11442 5964 11452 6020
rect 11508 5964 11676 6020
rect 11732 5964 11742 6020
rect 13122 5964 13132 6020
rect 13188 5964 13692 6020
rect 13748 5964 13758 6020
rect 14140 5964 18620 6020
rect 18676 5964 22540 6020
rect 22596 5964 24556 6020
rect 24612 5964 24622 6020
rect 25554 5964 25564 6020
rect 25620 5964 27020 6020
rect 27076 5964 27086 6020
rect 27458 5964 27468 6020
rect 27524 5964 28588 6020
rect 28644 5964 29148 6020
rect 29204 5964 29214 6020
rect 30604 5964 30828 6020
rect 30884 5964 32956 6020
rect 33012 5964 33964 6020
rect 34020 5964 34030 6020
rect 41010 5964 41020 6020
rect 41076 5964 41356 6020
rect 41412 5964 41422 6020
rect 46050 5964 46060 6020
rect 46116 5964 46956 6020
rect 47012 5964 47022 6020
rect 14140 5908 14196 5964
rect 30604 5908 30660 5964
rect 7634 5852 7644 5908
rect 7700 5852 8540 5908
rect 8596 5852 8606 5908
rect 8978 5852 8988 5908
rect 9044 5852 9660 5908
rect 9716 5852 9726 5908
rect 10210 5852 10220 5908
rect 10276 5852 10892 5908
rect 10948 5852 10958 5908
rect 14130 5852 14140 5908
rect 14196 5852 14206 5908
rect 14690 5852 14700 5908
rect 14756 5852 15148 5908
rect 15474 5852 15484 5908
rect 15540 5852 17612 5908
rect 17668 5852 17678 5908
rect 23762 5852 23772 5908
rect 23828 5852 24108 5908
rect 24164 5852 25340 5908
rect 25396 5852 25406 5908
rect 25778 5852 25788 5908
rect 25844 5852 26908 5908
rect 27794 5852 27804 5908
rect 27860 5852 28476 5908
rect 28532 5852 28542 5908
rect 30594 5852 30604 5908
rect 30660 5852 30670 5908
rect 32498 5852 32508 5908
rect 32564 5852 32844 5908
rect 32900 5852 34412 5908
rect 34468 5852 34478 5908
rect 15092 5796 15148 5852
rect 26852 5796 26908 5852
rect 4610 5740 4620 5796
rect 4676 5740 5628 5796
rect 5684 5740 5694 5796
rect 6290 5740 6300 5796
rect 6356 5740 7308 5796
rect 7364 5740 7374 5796
rect 8642 5740 8652 5796
rect 8708 5740 11228 5796
rect 11284 5740 11294 5796
rect 11442 5740 11452 5796
rect 11508 5740 11546 5796
rect 15092 5740 17724 5796
rect 17780 5740 18284 5796
rect 18340 5740 18350 5796
rect 18946 5740 18956 5796
rect 19012 5740 20076 5796
rect 20132 5740 21196 5796
rect 21252 5740 21262 5796
rect 21746 5740 21756 5796
rect 21812 5740 22316 5796
rect 22372 5740 23436 5796
rect 23492 5740 23502 5796
rect 26852 5740 27468 5796
rect 27524 5740 27860 5796
rect 28130 5740 28140 5796
rect 28196 5740 29036 5796
rect 29092 5740 29102 5796
rect 30818 5740 30828 5796
rect 30884 5740 31500 5796
rect 31556 5740 31566 5796
rect 32722 5740 32732 5796
rect 32788 5740 33740 5796
rect 33796 5740 33806 5796
rect 40898 5740 40908 5796
rect 40964 5740 43932 5796
rect 43988 5740 43998 5796
rect 27804 5684 27860 5740
rect 9986 5628 9996 5684
rect 10052 5628 10668 5684
rect 10724 5628 12572 5684
rect 12628 5628 12638 5684
rect 22978 5628 22988 5684
rect 23044 5628 24556 5684
rect 24612 5628 26908 5684
rect 27804 5628 31052 5684
rect 31108 5628 31118 5684
rect 32162 5628 32172 5684
rect 32228 5628 33180 5684
rect 33236 5628 33246 5684
rect 34066 5628 34076 5684
rect 34132 5628 34972 5684
rect 35028 5628 35038 5684
rect 35830 5628 35868 5684
rect 35924 5628 35934 5684
rect 26852 5572 26908 5628
rect 10882 5516 10892 5572
rect 10948 5516 12460 5572
rect 12516 5516 12526 5572
rect 14354 5516 14364 5572
rect 14420 5516 18508 5572
rect 18564 5516 18574 5572
rect 23874 5516 23884 5572
rect 23940 5516 24332 5572
rect 24388 5516 24398 5572
rect 26852 5516 32508 5572
rect 32564 5516 32574 5572
rect 33842 5516 33852 5572
rect 33908 5516 34188 5572
rect 34244 5516 34254 5572
rect 36754 5516 36764 5572
rect 36820 5516 37324 5572
rect 37380 5516 38780 5572
rect 38836 5516 38846 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 7634 5404 7644 5460
rect 7700 5404 8764 5460
rect 8820 5404 8830 5460
rect 12226 5404 12236 5460
rect 12292 5404 12572 5460
rect 12628 5404 14252 5460
rect 14308 5404 14318 5460
rect 22530 5404 22540 5460
rect 22596 5404 23324 5460
rect 23380 5404 24780 5460
rect 24836 5404 33516 5460
rect 33572 5404 34076 5460
rect 34132 5404 34142 5460
rect 38994 5404 39004 5460
rect 39060 5404 39788 5460
rect 39844 5404 39854 5460
rect 5730 5292 5740 5348
rect 5796 5292 8092 5348
rect 8148 5292 8158 5348
rect 11106 5292 11116 5348
rect 11172 5292 14364 5348
rect 14420 5292 14924 5348
rect 14980 5292 14990 5348
rect 19170 5292 19180 5348
rect 19236 5292 19628 5348
rect 19684 5292 19694 5348
rect 23426 5292 23436 5348
rect 23492 5292 24444 5348
rect 24500 5292 24510 5348
rect 31490 5292 31500 5348
rect 31556 5292 33404 5348
rect 33460 5292 34916 5348
rect 3826 5180 3836 5236
rect 3892 5180 4620 5236
rect 4676 5180 5068 5236
rect 5124 5180 6188 5236
rect 6244 5180 6692 5236
rect 10994 5180 11004 5236
rect 11060 5180 11070 5236
rect 12338 5180 12348 5236
rect 12404 5180 14028 5236
rect 14084 5180 16604 5236
rect 16660 5180 16670 5236
rect 18162 5180 18172 5236
rect 18228 5180 20748 5236
rect 20804 5180 20814 5236
rect 26450 5180 26460 5236
rect 26516 5180 27244 5236
rect 27300 5180 27310 5236
rect 31378 5180 31388 5236
rect 31444 5180 34636 5236
rect 34692 5180 34702 5236
rect 6636 5012 6692 5180
rect 7970 5068 7980 5124
rect 8036 5068 8652 5124
rect 8708 5068 8718 5124
rect 9538 5068 9548 5124
rect 9604 5068 10220 5124
rect 10276 5068 10286 5124
rect 11004 5012 11060 5180
rect 34860 5124 34916 5292
rect 12674 5068 12684 5124
rect 12740 5068 13580 5124
rect 13636 5068 13646 5124
rect 15250 5068 15260 5124
rect 15316 5068 15484 5124
rect 15540 5068 17052 5124
rect 17108 5068 17118 5124
rect 19618 5068 19628 5124
rect 19684 5068 20412 5124
rect 20468 5068 20478 5124
rect 21186 5068 21196 5124
rect 21252 5068 22204 5124
rect 22260 5068 22270 5124
rect 25778 5068 25788 5124
rect 25844 5068 27468 5124
rect 27524 5068 28028 5124
rect 28084 5068 28094 5124
rect 32050 5068 32060 5124
rect 32116 5068 33740 5124
rect 33796 5068 33806 5124
rect 34738 5068 34748 5124
rect 34804 5068 34916 5124
rect 46946 5068 46956 5124
rect 47012 5068 47852 5124
rect 47908 5068 47918 5124
rect 6636 4956 8764 5012
rect 8820 4956 9884 5012
rect 9940 4956 9950 5012
rect 11004 4956 13804 5012
rect 13860 4956 15148 5012
rect 16034 4956 16044 5012
rect 16100 4956 18396 5012
rect 18452 4956 18462 5012
rect 20290 4956 20300 5012
rect 20356 4956 21084 5012
rect 21140 4956 22764 5012
rect 22820 4956 23660 5012
rect 23716 4956 25004 5012
rect 25060 4956 25070 5012
rect 29362 4956 29372 5012
rect 29428 4956 30268 5012
rect 30324 4956 31612 5012
rect 31668 4956 31678 5012
rect 35970 4956 35980 5012
rect 36036 4956 37212 5012
rect 37268 4956 38892 5012
rect 38948 4956 38958 5012
rect 44482 4956 44492 5012
rect 44548 4956 47628 5012
rect 47684 4956 48188 5012
rect 48244 4956 48254 5012
rect 15092 4900 15148 4956
rect 8306 4844 8316 4900
rect 8372 4844 12796 4900
rect 12852 4844 12862 4900
rect 13234 4844 13244 4900
rect 13300 4844 14252 4900
rect 14308 4844 14318 4900
rect 15092 4844 19964 4900
rect 20020 4844 20030 4900
rect 22418 4844 22428 4900
rect 22484 4844 23100 4900
rect 23156 4844 23166 4900
rect 36082 4844 36092 4900
rect 36148 4844 38444 4900
rect 38500 4844 38510 4900
rect 42578 4844 42588 4900
rect 42644 4844 43708 4900
rect 43764 4844 43774 4900
rect 44146 4844 44156 4900
rect 44212 4844 44492 4900
rect 44548 4844 44940 4900
rect 44996 4844 45006 4900
rect 8418 4732 8428 4788
rect 8484 4732 9772 4788
rect 9828 4732 9838 4788
rect 10434 4732 10444 4788
rect 10500 4732 15596 4788
rect 15652 4732 15662 4788
rect 16482 4732 16492 4788
rect 16548 4732 17276 4788
rect 17332 4732 17342 4788
rect 18946 4732 18956 4788
rect 19012 4732 19292 4788
rect 19348 4732 19358 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 10770 4620 10780 4676
rect 10836 4620 11564 4676
rect 11620 4620 11630 4676
rect 12226 4620 12236 4676
rect 12292 4620 14924 4676
rect 14980 4620 14990 4676
rect 9874 4508 9884 4564
rect 9940 4508 13580 4564
rect 13636 4508 13646 4564
rect 14998 4508 15036 4564
rect 15092 4508 15102 4564
rect 19506 4508 19516 4564
rect 19572 4508 20076 4564
rect 20132 4508 20142 4564
rect 24098 4508 24108 4564
rect 24164 4508 26236 4564
rect 26292 4508 26302 4564
rect 39106 4508 39116 4564
rect 39172 4508 40124 4564
rect 40180 4508 41020 4564
rect 41076 4508 42588 4564
rect 42644 4508 42654 4564
rect 13010 4396 13020 4452
rect 13076 4396 34860 4452
rect 34916 4396 34926 4452
rect 20738 4284 20748 4340
rect 20804 4284 21420 4340
rect 21476 4284 21486 4340
rect 14130 4172 14140 4228
rect 14196 4172 18060 4228
rect 18116 4172 18126 4228
rect 18274 4172 18284 4228
rect 18340 4172 19516 4228
rect 19572 4172 19582 4228
rect 23090 4172 23100 4228
rect 23156 4172 23660 4228
rect 23716 4172 23726 4228
rect 36278 4172 36316 4228
rect 36372 4172 36382 4228
rect 18386 4060 18396 4116
rect 18452 4060 31164 4116
rect 31220 4060 31230 4116
rect 39666 4060 39676 4116
rect 39732 4060 41916 4116
rect 41972 4060 41982 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 15138 3836 15148 3892
rect 15204 3836 15214 3892
rect 15148 3780 15204 3836
rect 9986 3724 9996 3780
rect 10052 3724 15204 3780
rect 8866 3612 8876 3668
rect 8932 3612 10780 3668
rect 10836 3612 10846 3668
rect 13570 3612 13580 3668
rect 13636 3612 17724 3668
rect 17780 3612 17790 3668
rect 18834 3612 18844 3668
rect 18900 3612 21420 3668
rect 21476 3612 21868 3668
rect 21924 3612 24108 3668
rect 24164 3612 24174 3668
rect 26226 3612 26236 3668
rect 26292 3612 28588 3668
rect 28644 3612 28654 3668
rect 42578 3612 42588 3668
rect 42644 3612 43820 3668
rect 43876 3612 43886 3668
rect 37874 3500 37884 3556
rect 37940 3500 47628 3556
rect 47684 3500 47694 3556
rect 9538 3388 9548 3444
rect 9604 3388 10892 3444
rect 10948 3388 11788 3444
rect 11844 3388 12684 3444
rect 12740 3388 15260 3444
rect 15316 3388 15326 3444
rect 46946 3388 46956 3444
rect 47012 3388 48076 3444
rect 48132 3388 48142 3444
rect 4050 3276 4060 3332
rect 4116 3276 25228 3332
rect 25284 3276 25294 3332
rect 23650 3164 23660 3220
rect 23716 3164 33628 3220
rect 33684 3164 33694 3220
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 9314 2940 9324 2996
rect 9380 2940 28924 2996
rect 28980 2940 28990 2996
rect 3378 2828 3388 2884
rect 3444 2828 21084 2884
rect 21140 2828 21150 2884
rect 49200 2772 50000 2800
rect 9538 2716 9548 2772
rect 9604 2716 27580 2772
rect 27636 2716 27646 2772
rect 48178 2716 48188 2772
rect 48244 2716 50000 2772
rect 49200 2688 50000 2716
rect 9538 2604 9548 2660
rect 9604 2604 34412 2660
rect 34468 2604 34478 2660
rect 18498 2492 18508 2548
rect 18564 2492 23660 2548
rect 23716 2492 23726 2548
rect 13346 2380 13356 2436
rect 13412 2380 23548 2436
rect 23604 2380 23614 2436
rect 6738 2268 6748 2324
rect 6804 2268 32284 2324
rect 32340 2268 32350 2324
rect 12786 1596 12796 1652
rect 12852 1596 24892 1652
rect 24948 1596 24958 1652
rect 12898 1484 12908 1540
rect 12964 1484 30380 1540
rect 30436 1484 30446 1540
rect 10770 1372 10780 1428
rect 10836 1372 24556 1428
rect 24612 1372 24622 1428
rect 15026 1260 15036 1316
rect 15092 1260 25788 1316
rect 25844 1260 25854 1316
rect 7634 1148 7644 1204
rect 7700 1148 25788 1204
rect 25844 1148 25854 1204
<< via3 >>
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 48076 44156 48132 44212
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 37548 43484 37604 43540
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 38892 42812 38948 42868
rect 43708 42812 43764 42868
rect 45164 42812 45220 42868
rect 25340 42588 25396 42644
rect 16716 42476 16772 42532
rect 40012 42476 40068 42532
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 44940 42028 44996 42084
rect 43708 41804 43764 41860
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 26124 40908 26180 40964
rect 38892 41132 38948 41188
rect 41244 41020 41300 41076
rect 44940 41020 44996 41076
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 43484 40460 43540 40516
rect 13132 40348 13188 40404
rect 14476 40236 14532 40292
rect 40012 40124 40068 40180
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 11004 38892 11060 38948
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 17724 38220 17780 38276
rect 37548 38108 37604 38164
rect 45164 37884 45220 37940
rect 48076 37884 48132 37940
rect 5516 37772 5572 37828
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 37548 37548 37604 37604
rect 44492 37436 44548 37492
rect 26124 37212 26180 37268
rect 18844 37100 18900 37156
rect 18732 36988 18788 37044
rect 43484 36988 43540 37044
rect 44492 36876 44548 36932
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 5516 36764 5572 36820
rect 8540 36764 8596 36820
rect 19628 36316 19684 36372
rect 7532 36204 7588 36260
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 14476 35980 14532 36036
rect 19628 35980 19684 36036
rect 23212 35756 23268 35812
rect 25340 35756 25396 35812
rect 41244 35532 41300 35588
rect 8540 35420 8596 35476
rect 16716 35420 16772 35476
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 16604 35196 16660 35252
rect 19516 35084 19572 35140
rect 34636 35084 34692 35140
rect 35644 35084 35700 35140
rect 19628 34860 19684 34916
rect 18508 34748 18564 34804
rect 5180 34636 5236 34692
rect 13132 34636 13188 34692
rect 35644 34636 35700 34692
rect 6076 34412 6132 34468
rect 23884 34524 23940 34580
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 23996 34412 24052 34468
rect 22652 34188 22708 34244
rect 29596 34300 29652 34356
rect 18732 34076 18788 34132
rect 19516 34076 19572 34132
rect 23884 33740 23940 33796
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 5628 33628 5684 33684
rect 1708 33180 1764 33236
rect 4172 33180 4228 33236
rect 7532 33180 7588 33236
rect 14924 33180 14980 33236
rect 2044 33068 2100 33124
rect 13692 33068 13748 33124
rect 20412 33068 20468 33124
rect 2268 32956 2324 33012
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 16492 32844 16548 32900
rect 23436 32844 23492 32900
rect 4956 32732 5012 32788
rect 26684 32732 26740 32788
rect 3388 32620 3444 32676
rect 14924 32396 14980 32452
rect 2604 32172 2660 32228
rect 8428 32172 8484 32228
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 8540 32060 8596 32116
rect 11004 31948 11060 32004
rect 22652 31724 22708 31780
rect 8876 31612 8932 31668
rect 2604 31500 2660 31556
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 13580 31276 13636 31332
rect 5292 30940 5348 30996
rect 22428 30828 22484 30884
rect 21532 30716 21588 30772
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 17948 30492 18004 30548
rect 25900 30380 25956 30436
rect 5068 30268 5124 30324
rect 16604 30268 16660 30324
rect 19068 30268 19124 30324
rect 19628 30268 19684 30324
rect 23996 30268 24052 30324
rect 3388 30156 3444 30212
rect 8876 30156 8932 30212
rect 16492 30156 16548 30212
rect 21308 30156 21364 30212
rect 2268 30044 2324 30100
rect 4172 30044 4228 30100
rect 18844 30044 18900 30100
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 23436 29708 23492 29764
rect 2044 29484 2100 29540
rect 8428 29484 8484 29540
rect 8540 29260 8596 29316
rect 5068 29148 5124 29204
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 13580 29484 13636 29540
rect 17948 29484 18004 29540
rect 20412 29484 20468 29540
rect 5628 29148 5684 29204
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 13692 28924 13748 28980
rect 26236 28924 26292 28980
rect 6076 28812 6132 28868
rect 18508 28812 18564 28868
rect 4956 28700 5012 28756
rect 1708 28588 1764 28644
rect 18844 28588 18900 28644
rect 26236 28476 26292 28532
rect 22428 28364 22484 28420
rect 5180 28252 5236 28308
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 19068 28140 19124 28196
rect 21532 28140 21588 28196
rect 18508 27692 18564 27748
rect 19628 27580 19684 27636
rect 34636 27468 34692 27524
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 6860 27132 6916 27188
rect 20188 27132 20244 27188
rect 6076 26684 6132 26740
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 25900 26460 25956 26516
rect 26684 26460 26740 26516
rect 17948 25900 18004 25956
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 18284 25676 18340 25732
rect 21308 25676 21364 25732
rect 19068 25340 19124 25396
rect 18508 25228 18564 25284
rect 19628 25228 19684 25284
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 5292 24892 5348 24948
rect 17948 24780 18004 24836
rect 18284 24780 18340 24836
rect 18844 24780 18900 24836
rect 25228 24668 25284 24724
rect 19628 24332 19684 24388
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 6860 23884 6916 23940
rect 17500 23884 17556 23940
rect 29596 23884 29652 23940
rect 17612 23548 17668 23604
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 23212 23324 23268 23380
rect 27916 23212 27972 23268
rect 19068 22876 19124 22932
rect 27916 22764 27972 22820
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19180 22540 19236 22596
rect 25340 22428 25396 22484
rect 25116 22204 25172 22260
rect 37436 22204 37492 22260
rect 20188 22092 20244 22148
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 25340 21756 25396 21812
rect 20300 21644 20356 21700
rect 5068 21532 5124 21588
rect 17500 21420 17556 21476
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 4060 20972 4116 21028
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19292 20860 19348 20916
rect 19404 20636 19460 20692
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 17500 20300 17556 20356
rect 18396 20300 18452 20356
rect 25116 20188 25172 20244
rect 19180 20076 19236 20132
rect 17612 19964 17668 20020
rect 19292 19852 19348 19908
rect 23884 19740 23940 19796
rect 19292 19628 19348 19684
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 17388 19516 17444 19572
rect 23660 19516 23716 19572
rect 23884 19516 23940 19572
rect 17164 19292 17220 19348
rect 19628 19292 19684 19348
rect 20300 19180 20356 19236
rect 25116 19180 25172 19236
rect 6076 19068 6132 19124
rect 18396 18844 18452 18900
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 16828 18732 16884 18788
rect 17388 18732 17444 18788
rect 17612 18732 17668 18788
rect 20748 18732 20804 18788
rect 23660 18732 23716 18788
rect 14588 18620 14644 18676
rect 37436 18508 37492 18564
rect 10220 18396 10276 18452
rect 16940 18284 16996 18340
rect 17724 18284 17780 18340
rect 23660 18284 23716 18340
rect 23884 18172 23940 18228
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 20748 17948 20804 18004
rect 10220 17836 10276 17892
rect 20412 17836 20468 17892
rect 18284 17724 18340 17780
rect 23436 17612 23492 17668
rect 28364 17500 28420 17556
rect 25788 17388 25844 17444
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4956 17164 5012 17220
rect 19628 17164 19684 17220
rect 20188 17164 20244 17220
rect 10108 17052 10164 17108
rect 20412 17052 20468 17108
rect 4060 16828 4116 16884
rect 5068 16828 5124 16884
rect 18396 16828 18452 16884
rect 25788 16828 25844 16884
rect 6076 16604 6132 16660
rect 4956 16492 5012 16548
rect 18284 16492 18340 16548
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 17500 16380 17556 16436
rect 5068 16044 5124 16100
rect 19404 16044 19460 16100
rect 20412 16044 20468 16100
rect 4844 15932 4900 15988
rect 20748 15932 20804 15988
rect 22876 15932 22932 15988
rect 25340 15932 25396 15988
rect 6188 15820 6244 15876
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 18284 15596 18340 15652
rect 6412 15260 6468 15316
rect 25340 15260 25396 15316
rect 17164 15148 17220 15204
rect 21756 15036 21812 15092
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19628 14700 19684 14756
rect 18396 14588 18452 14644
rect 28364 14588 28420 14644
rect 4844 14364 4900 14420
rect 21756 14364 21812 14420
rect 23100 14364 23156 14420
rect 26348 14252 26404 14308
rect 18620 14140 18676 14196
rect 27580 14140 27636 14196
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 7532 14028 7588 14084
rect 13804 14028 13860 14084
rect 25676 14028 25732 14084
rect 10220 13804 10276 13860
rect 26908 13804 26964 13860
rect 27580 13804 27636 13860
rect 15372 13692 15428 13748
rect 19404 13692 19460 13748
rect 38612 13692 38668 13748
rect 15036 13580 15092 13636
rect 25564 13580 25620 13636
rect 25788 13580 25844 13636
rect 31164 13580 31220 13636
rect 18844 13468 18900 13524
rect 25452 13468 25508 13524
rect 26348 13468 26404 13524
rect 26908 13468 26964 13524
rect 34412 13356 34468 13412
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 6412 13244 6468 13300
rect 22876 13244 22932 13300
rect 25676 13244 25732 13300
rect 25452 13020 25508 13076
rect 23436 12908 23492 12964
rect 13468 12796 13524 12852
rect 19292 12796 19348 12852
rect 38556 12796 38612 12852
rect 7532 12684 7588 12740
rect 23100 12572 23156 12628
rect 25564 12572 25620 12628
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 6188 12460 6244 12516
rect 13804 12460 13860 12516
rect 14588 12348 14644 12404
rect 25340 12348 25396 12404
rect 31164 12348 31220 12404
rect 19404 12236 19460 12292
rect 14812 12124 14868 12180
rect 17612 12124 17668 12180
rect 19068 12124 19124 12180
rect 18060 12012 18116 12068
rect 18844 11900 18900 11956
rect 10220 11788 10276 11844
rect 18060 11788 18116 11844
rect 18284 11788 18340 11844
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 13356 11452 13412 11508
rect 15260 11452 15316 11508
rect 35980 11340 36036 11396
rect 6972 11116 7028 11172
rect 27804 11116 27860 11172
rect 14252 11004 14308 11060
rect 14812 11004 14868 11060
rect 21084 11004 21140 11060
rect 34412 11004 34468 11060
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 21420 10892 21476 10948
rect 14252 10668 14308 10724
rect 18956 10668 19012 10724
rect 12572 10556 12628 10612
rect 12908 10444 12964 10500
rect 15260 10444 15316 10500
rect 23548 10332 23604 10388
rect 15372 10220 15428 10276
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 18956 10108 19012 10164
rect 10108 9884 10164 9940
rect 21084 9884 21140 9940
rect 10332 9548 10388 9604
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 16828 9212 16884 9268
rect 13356 9100 13412 9156
rect 37212 8988 37268 9044
rect 19292 8876 19348 8932
rect 13468 8764 13524 8820
rect 7644 8652 7700 8708
rect 36316 8652 36372 8708
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 6860 8428 6916 8484
rect 26908 8428 26964 8484
rect 35980 8428 36036 8484
rect 19292 8316 19348 8372
rect 21420 8204 21476 8260
rect 35644 7980 35700 8036
rect 16940 7868 16996 7924
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 16940 7644 16996 7700
rect 35868 7644 35924 7700
rect 18620 7532 18676 7588
rect 44492 7532 44548 7588
rect 6972 7420 7028 7476
rect 18396 7308 18452 7364
rect 27468 7308 27524 7364
rect 21420 7084 21476 7140
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 35644 6972 35700 7028
rect 27804 6860 27860 6916
rect 9548 6748 9604 6804
rect 11452 6748 11508 6804
rect 6860 6636 6916 6692
rect 27468 6636 27524 6692
rect 36316 6636 36372 6692
rect 12572 6524 12628 6580
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 37212 6076 37268 6132
rect 27468 5964 27524 6020
rect 11452 5740 11508 5796
rect 35868 5628 35924 5684
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 44492 4844 44548 4900
rect 18956 4732 19012 4788
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 15036 4508 15092 4564
rect 36316 4172 36372 4228
rect 18396 4060 18452 4116
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 25228 3276 25284 3332
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 9548 2604 9604 2660
rect 13356 2380 13412 2436
rect 23548 2380 23604 2436
rect 12908 1484 12964 1540
rect 7644 1148 7700 1204
rect 25788 1148 25844 1204
<< metal4 >>
rect 4448 46284 4768 46316
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 19808 45500 20128 46316
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 16716 42532 16772 42542
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 13132 40404 13188 40414
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 11004 38948 11060 38958
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 5516 37828 5572 37838
rect 5516 36820 5572 37772
rect 5516 36754 5572 36764
rect 8540 36820 8596 36830
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 7532 36260 7588 36270
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 1708 33236 1764 33246
rect 1708 28644 1764 33180
rect 4172 33236 4228 33246
rect 2044 33124 2100 33134
rect 2044 29540 2100 33068
rect 2268 33012 2324 33022
rect 2268 30100 2324 32956
rect 3388 32676 3444 32686
rect 2604 32228 2660 32238
rect 2604 31556 2660 32172
rect 2604 31490 2660 31500
rect 3388 30212 3444 32620
rect 3388 30146 3444 30156
rect 2268 30034 2324 30044
rect 4172 30100 4228 33180
rect 4172 30034 4228 30044
rect 4448 32172 4768 33684
rect 5180 34692 5236 34702
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 2044 29474 2100 29484
rect 1708 28578 1764 28588
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4956 32788 5012 32798
rect 4956 28756 5012 32732
rect 5068 30324 5124 30334
rect 5068 29204 5124 30268
rect 5068 29138 5124 29148
rect 4956 28690 5012 28700
rect 5180 28308 5236 34636
rect 6076 34468 6132 34478
rect 5628 33684 5684 33694
rect 5180 28242 5236 28252
rect 5292 30996 5348 31006
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 5292 24948 5348 30940
rect 5628 29204 5684 33628
rect 5628 29138 5684 29148
rect 6076 28868 6132 34412
rect 7532 33236 7588 36204
rect 8540 35476 8596 36764
rect 8540 35410 8596 35420
rect 7532 33170 7588 33180
rect 8428 32228 8484 32238
rect 8428 29540 8484 32172
rect 8428 29474 8484 29484
rect 8540 32116 8596 32126
rect 8540 29316 8596 32060
rect 11004 32004 11060 38892
rect 13132 34692 13188 40348
rect 14476 40292 14532 40302
rect 14476 36036 14532 40236
rect 14476 35970 14532 35980
rect 16716 35476 16772 42476
rect 19808 42364 20128 43876
rect 35168 46284 35488 46316
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 48076 44212 48132 44222
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 16716 35410 16772 35420
rect 17724 38276 17780 38286
rect 13132 34626 13188 34636
rect 16604 35252 16660 35262
rect 14924 33236 14980 33246
rect 11004 31938 11060 31948
rect 13692 33124 13748 33134
rect 8876 31668 8932 31678
rect 8876 30212 8932 31612
rect 8876 30146 8932 30156
rect 13580 31332 13636 31342
rect 13580 29540 13636 31276
rect 13580 29474 13636 29484
rect 8540 29250 8596 29260
rect 13692 28980 13748 33068
rect 14924 32452 14980 33180
rect 14924 32386 14980 32396
rect 16492 32900 16548 32910
rect 16492 30212 16548 32844
rect 16604 30324 16660 35196
rect 16604 30258 16660 30268
rect 16492 30146 16548 30156
rect 13692 28914 13748 28924
rect 6076 26740 6132 28812
rect 6076 26674 6132 26684
rect 6860 27188 6916 27198
rect 5292 24882 5348 24892
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 6860 23940 6916 27132
rect 6860 23874 6916 23884
rect 17500 23940 17556 23950
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4060 21028 4116 21038
rect 4060 16884 4116 20972
rect 4060 16818 4116 16828
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 5068 21588 5124 21598
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4956 17220 5012 17230
rect 4956 16548 5012 17164
rect 4956 16482 5012 16492
rect 5068 16884 5124 21532
rect 17500 21476 17556 23884
rect 17500 21410 17556 21420
rect 17612 23604 17668 23614
rect 17500 20356 17556 20366
rect 17388 19572 17444 19582
rect 17164 19348 17220 19358
rect 4448 14924 4768 16436
rect 5068 16100 5124 16828
rect 6076 19124 6132 19134
rect 6076 16660 6132 19068
rect 16828 18788 16884 18798
rect 14588 18676 14644 18686
rect 10220 18452 10276 18462
rect 10220 17892 10276 18396
rect 6076 16594 6132 16604
rect 10108 17108 10164 17118
rect 5068 16034 5124 16044
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4844 15988 4900 15998
rect 4844 14420 4900 15932
rect 4844 14354 4900 14364
rect 6188 15876 6244 15886
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 6188 12516 6244 15820
rect 6412 15316 6468 15326
rect 6412 13300 6468 15260
rect 6412 13234 6468 13244
rect 7532 14084 7588 14094
rect 7532 12740 7588 14028
rect 7532 12674 7588 12684
rect 6188 12450 6244 12460
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 6972 11172 7028 11182
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 6860 8484 6916 8494
rect 6860 6692 6916 8428
rect 6972 7476 7028 11116
rect 10108 9940 10164 17052
rect 10220 15148 10276 17836
rect 10220 15092 10388 15148
rect 10220 13860 10276 13870
rect 10220 11844 10276 13804
rect 10220 11778 10276 11788
rect 10108 9874 10164 9884
rect 10332 9604 10388 15092
rect 13804 14084 13860 14094
rect 13468 12852 13524 12862
rect 13356 11508 13412 11518
rect 10332 9538 10388 9548
rect 12572 10612 12628 10622
rect 6972 7410 7028 7420
rect 7644 8708 7700 8718
rect 6860 6626 6916 6636
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 7644 1204 7700 8652
rect 9548 6804 9604 6814
rect 9548 2660 9604 6748
rect 11452 6804 11508 6814
rect 11452 5796 11508 6748
rect 12572 6580 12628 10556
rect 12572 6514 12628 6524
rect 12908 10500 12964 10510
rect 11452 5730 11508 5740
rect 9548 2594 9604 2604
rect 12908 1540 12964 10444
rect 13356 9156 13412 11452
rect 13356 2436 13412 9100
rect 13468 8820 13524 12796
rect 13804 12516 13860 14028
rect 13804 12450 13860 12460
rect 14588 12404 14644 18620
rect 15372 13748 15428 13758
rect 14588 12338 14644 12348
rect 15036 13636 15092 13646
rect 14812 12180 14868 12190
rect 14252 11060 14308 11070
rect 14252 10724 14308 11004
rect 14812 11060 14868 12124
rect 14812 10994 14868 11004
rect 14252 10658 14308 10668
rect 13468 8754 13524 8764
rect 15036 4564 15092 13580
rect 15260 11508 15316 11518
rect 15260 10500 15316 11452
rect 15260 10434 15316 10444
rect 15372 10276 15428 13692
rect 15372 10210 15428 10220
rect 16828 9268 16884 18732
rect 16828 9202 16884 9212
rect 16940 18340 16996 18350
rect 16940 7924 16996 18284
rect 17164 15204 17220 19292
rect 17388 18788 17444 19516
rect 17388 18722 17444 18732
rect 17500 16436 17556 20300
rect 17612 20020 17668 23548
rect 17612 19954 17668 19964
rect 17500 16370 17556 16380
rect 17612 18788 17668 18798
rect 17164 15138 17220 15148
rect 17612 12180 17668 18732
rect 17724 18340 17780 38220
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 18844 37156 18900 37166
rect 18732 37044 18788 37054
rect 18508 34804 18564 34814
rect 17948 30548 18004 30558
rect 17948 29540 18004 30492
rect 17948 29474 18004 29484
rect 18508 28868 18564 34748
rect 18732 34132 18788 36988
rect 18732 34066 18788 34076
rect 18844 30100 18900 37100
rect 19628 36372 19684 36382
rect 19628 36036 19684 36316
rect 19628 35970 19684 35980
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19516 35140 19572 35150
rect 19516 34132 19572 35084
rect 19516 34066 19572 34076
rect 19628 34916 19684 34926
rect 18844 30034 18900 30044
rect 19068 30324 19124 30334
rect 18508 28802 18564 28812
rect 18844 28644 18900 28654
rect 18508 27748 18564 27758
rect 17948 25956 18004 25966
rect 17948 24836 18004 25900
rect 17948 24770 18004 24780
rect 18284 25732 18340 25742
rect 18284 24836 18340 25676
rect 18508 25284 18564 27692
rect 18508 25218 18564 25228
rect 18284 24770 18340 24780
rect 18844 24836 18900 28588
rect 19068 28196 19124 30268
rect 19628 30324 19684 34860
rect 19628 30258 19684 30268
rect 19808 34524 20128 36036
rect 25340 42644 25396 42654
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 23212 35812 23268 35822
rect 22652 34244 22708 34254
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19068 25396 19124 28140
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 20412 33124 20468 33134
rect 20412 29540 20468 33068
rect 22652 31780 22708 34188
rect 22652 31714 22708 31724
rect 22428 30884 22484 30894
rect 21532 30772 21588 30782
rect 20412 29474 20468 29484
rect 21308 30212 21364 30222
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19068 25330 19124 25340
rect 19628 27636 19684 27646
rect 18844 24770 18900 24780
rect 19628 25284 19684 27580
rect 19628 24388 19684 25228
rect 19068 22932 19124 22942
rect 18396 20356 18452 20366
rect 18396 18900 18452 20300
rect 18396 18834 18452 18844
rect 17724 18274 17780 18284
rect 18284 17780 18340 17790
rect 18284 16548 18340 17724
rect 18284 16482 18340 16492
rect 18396 16884 18452 16894
rect 17612 12114 17668 12124
rect 18284 15652 18340 15662
rect 18060 12068 18116 12078
rect 18060 11844 18116 12012
rect 18060 11778 18116 11788
rect 18284 11844 18340 15596
rect 18284 11778 18340 11788
rect 18396 14644 18452 16828
rect 16940 7700 16996 7868
rect 16940 7634 16996 7644
rect 15036 4498 15092 4508
rect 18396 7364 18452 14588
rect 18620 14196 18676 14206
rect 18620 7588 18676 14140
rect 18844 13524 18900 13534
rect 18844 11956 18900 13468
rect 19068 12180 19124 22876
rect 19180 22596 19236 22606
rect 19180 20132 19236 22540
rect 19180 20066 19236 20076
rect 19292 20916 19348 20926
rect 19292 19908 19348 20860
rect 19292 19842 19348 19852
rect 19404 20692 19460 20702
rect 19292 19684 19348 19694
rect 19292 12852 19348 19628
rect 19292 12786 19348 12796
rect 19404 16100 19460 20636
rect 19628 19348 19684 24332
rect 19628 19282 19684 19292
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19404 13748 19460 16044
rect 19628 17220 19684 17230
rect 19628 14756 19684 17164
rect 19628 14690 19684 14700
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 20188 27188 20244 27198
rect 20188 22148 20244 27132
rect 21308 25732 21364 30156
rect 21532 28196 21588 30716
rect 22428 28420 22484 30828
rect 22428 28354 22484 28364
rect 21532 28130 21588 28140
rect 21308 25666 21364 25676
rect 23212 23380 23268 35756
rect 25340 35812 25396 42588
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 26124 40964 26180 40974
rect 26124 37268 26180 40908
rect 26124 37202 26180 37212
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 25340 35746 25396 35756
rect 35168 36876 35488 38388
rect 37548 43540 37604 43550
rect 37548 38164 37604 43484
rect 38892 42868 38948 42878
rect 38892 41188 38948 42812
rect 43708 42868 43764 42878
rect 38892 41122 38948 41132
rect 40012 42532 40068 42542
rect 40012 40180 40068 42476
rect 43708 41860 43764 42812
rect 45164 42868 45220 42878
rect 43708 41794 43764 41804
rect 44940 42084 44996 42094
rect 40012 40114 40068 40124
rect 41244 41076 41300 41086
rect 37548 37604 37604 38108
rect 37548 37538 37604 37548
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 41244 35588 41300 41020
rect 44940 41076 44996 42028
rect 44940 41010 44996 41020
rect 43484 40516 43540 40526
rect 43484 37044 43540 40460
rect 45164 37940 45220 42812
rect 45164 37874 45220 37884
rect 48076 37940 48132 44156
rect 48076 37874 48132 37884
rect 43484 36978 43540 36988
rect 44492 37492 44548 37502
rect 44492 36932 44548 37436
rect 44492 36866 44548 36876
rect 41244 35522 41300 35532
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 34636 35140 34692 35150
rect 23884 34580 23940 34590
rect 23884 33796 23940 34524
rect 23884 33730 23940 33740
rect 23996 34468 24052 34478
rect 23436 32900 23492 32910
rect 23436 29764 23492 32844
rect 23996 30324 24052 34412
rect 29596 34356 29652 34366
rect 26684 32788 26740 32798
rect 23996 30258 24052 30268
rect 25900 30436 25956 30446
rect 23436 29698 23492 29708
rect 25900 26516 25956 30380
rect 26236 28980 26292 28990
rect 26236 28532 26292 28924
rect 26236 28466 26292 28476
rect 25900 26450 25956 26460
rect 26684 26516 26740 32732
rect 26684 26450 26740 26460
rect 23212 23314 23268 23324
rect 25228 24724 25284 24734
rect 20188 17220 20244 22092
rect 25116 22260 25172 22270
rect 20300 21700 20356 21710
rect 20300 19236 20356 21644
rect 25116 20244 25172 22204
rect 23884 19796 23940 19806
rect 20300 19170 20356 19180
rect 23660 19572 23716 19582
rect 20748 18788 20804 18798
rect 20748 18004 20804 18732
rect 23660 18788 23716 19516
rect 23660 18340 23716 18732
rect 23660 18274 23716 18284
rect 23884 19572 23940 19740
rect 23884 18228 23940 19516
rect 25116 19236 25172 20188
rect 25116 19170 25172 19180
rect 23884 18162 23940 18172
rect 20188 17154 20244 17164
rect 20412 17892 20468 17902
rect 20412 17108 20468 17836
rect 20412 16100 20468 17052
rect 20412 16034 20468 16044
rect 20748 15988 20804 17948
rect 23436 17668 23492 17678
rect 20748 15922 20804 15932
rect 22876 15988 22932 15998
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19404 12292 19460 13692
rect 19404 12226 19460 12236
rect 19808 14140 20128 15652
rect 21756 15092 21812 15102
rect 21756 14420 21812 15036
rect 21756 14354 21812 14364
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 22876 13300 22932 15932
rect 22876 13234 22932 13244
rect 23100 14420 23156 14430
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 23100 12628 23156 14364
rect 23436 12964 23492 17612
rect 23436 12898 23492 12908
rect 23100 12562 23156 12572
rect 19068 12114 19124 12124
rect 18844 11890 18900 11900
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 18620 7522 18676 7532
rect 18956 10724 19012 10734
rect 18956 10164 19012 10668
rect 18396 4116 18452 7308
rect 18956 4788 19012 10108
rect 19808 9436 20128 10948
rect 21084 11060 21140 11070
rect 21084 9940 21140 11004
rect 21084 9874 21140 9884
rect 21420 10948 21476 10958
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19292 8932 19348 8942
rect 19292 8372 19348 8876
rect 19292 8306 19348 8316
rect 18956 4722 19012 4732
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 21420 8260 21476 10892
rect 21420 7140 21476 8204
rect 21420 7074 21476 7084
rect 23548 10388 23604 10398
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 18396 4050 18452 4060
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 13356 2370 13412 2380
rect 23548 2436 23604 10332
rect 25228 3332 25284 24668
rect 29596 23940 29652 34300
rect 34636 27524 34692 35084
rect 34636 27458 34692 27468
rect 35168 33740 35488 35252
rect 35644 35140 35700 35150
rect 35644 34692 35700 35084
rect 35644 34626 35700 34636
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 29596 23874 29652 23884
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 27916 23268 27972 23278
rect 27916 22820 27972 23212
rect 27916 22754 27972 22764
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 25340 22484 25396 22494
rect 25340 21812 25396 22428
rect 25340 21746 25396 21756
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 37436 22260 37492 22270
rect 37436 18564 37492 22204
rect 37436 18498 37492 18508
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 28364 17556 28420 17566
rect 25788 17444 25844 17454
rect 25788 16884 25844 17388
rect 25340 15988 25396 15998
rect 25340 15316 25396 15932
rect 25340 12404 25396 15260
rect 25676 14084 25732 14094
rect 25564 13636 25620 13646
rect 25452 13524 25508 13534
rect 25452 13076 25508 13468
rect 25452 13010 25508 13020
rect 25564 12628 25620 13580
rect 25676 13300 25732 14028
rect 25676 13234 25732 13244
rect 25788 13636 25844 16828
rect 28364 14644 28420 17500
rect 28364 14578 28420 14588
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 25564 12562 25620 12572
rect 25340 12338 25396 12348
rect 25228 3266 25284 3276
rect 23548 2370 23604 2380
rect 12908 1474 12964 1484
rect 7644 1138 7700 1148
rect 25788 1204 25844 13580
rect 26348 14308 26404 14318
rect 26348 13524 26404 14252
rect 27580 14196 27636 14206
rect 26348 13458 26404 13468
rect 26908 13860 26964 13870
rect 26908 13524 26964 13804
rect 27580 13860 27636 14140
rect 27580 13794 27636 13804
rect 26908 8484 26964 13468
rect 31164 13636 31220 13646
rect 31164 12404 31220 13580
rect 31164 12338 31220 12348
rect 34412 13412 34468 13422
rect 26908 8418 26964 8428
rect 27804 11172 27860 11182
rect 27468 7364 27524 7374
rect 27468 6692 27524 7308
rect 27804 6916 27860 11116
rect 34412 11060 34468 13356
rect 34412 10994 34468 11004
rect 35168 13356 35488 14868
rect 38612 13748 38668 13758
rect 38612 13618 38668 13692
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 38556 13562 38668 13618
rect 38556 12852 38612 13562
rect 38556 12786 38612 12796
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 27804 6850 27860 6860
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35980 11396 36036 11406
rect 35980 8484 36036 11340
rect 37212 9044 37268 9054
rect 35980 8418 36036 8428
rect 36316 8708 36372 8718
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 27468 6020 27524 6636
rect 27468 5954 27524 5964
rect 35168 5516 35488 7028
rect 35644 8036 35700 8046
rect 35644 7028 35700 7980
rect 35644 6962 35700 6972
rect 35868 7700 35924 7710
rect 35868 5684 35924 7644
rect 35868 5618 35924 5628
rect 36316 6692 36372 8652
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 36316 4228 36372 6636
rect 37212 6132 37268 8988
rect 37212 6066 37268 6076
rect 44492 7588 44548 7598
rect 44492 4900 44548 7532
rect 44492 4834 44548 4844
rect 36316 4162 36372 4172
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 25788 1138 25844 1148
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1259_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1260_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19376 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1261_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 21728 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1262_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18704 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1263_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20496 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1264_
timestamp 1698431365
transform -1 0 23408 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1265_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21392 0 1 25088
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1266_
timestamp 1698431365
transform -1 0 17024 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1267_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19936 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1268_
timestamp 1698431365
transform 1 0 12208 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1269_
timestamp 1698431365
transform -1 0 19712 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1270_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22624 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1271_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23632 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1272_
timestamp 1698431365
transform 1 0 21392 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1273_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22288 0 1 26656
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1274_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19040 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1275_
timestamp 1698431365
transform 1 0 20048 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1276_
timestamp 1698431365
transform 1 0 19264 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1277_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15008 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1278_
timestamp 1698431365
transform 1 0 19264 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1279_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22624 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1280_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32704 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1281_
timestamp 1698431365
transform -1 0 31920 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1282_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1283_
timestamp 1698431365
transform -1 0 23968 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1284_
timestamp 1698431365
transform 1 0 24864 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1285_
timestamp 1698431365
transform -1 0 30800 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1286_
timestamp 1698431365
transform -1 0 28336 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1287_
timestamp 1698431365
transform 1 0 32032 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1288_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22064 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1289_
timestamp 1698431365
transform -1 0 31136 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1290_
timestamp 1698431365
transform 1 0 30352 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1291_
timestamp 1698431365
transform -1 0 30688 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1292_
timestamp 1698431365
transform -1 0 29904 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1293_
timestamp 1698431365
transform -1 0 29904 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1294_
timestamp 1698431365
transform -1 0 31248 0 -1 26656
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1295_
timestamp 1698431365
transform -1 0 27552 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1296_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 27328 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1297_
timestamp 1698431365
transform 1 0 34272 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1298_
timestamp 1698431365
transform -1 0 34720 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1299_
timestamp 1698431365
transform -1 0 30688 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1300_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28000 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1301_
timestamp 1698431365
transform -1 0 11872 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _1302_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19824 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1303_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11760 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1304_
timestamp 1698431365
transform -1 0 17024 0 -1 23520
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1305_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _1306_
timestamp 1698431365
transform -1 0 9184 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _1307_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9520 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1308_
timestamp 1698431365
transform 1 0 10192 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1309_
timestamp 1698431365
transform 1 0 15344 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1310_
timestamp 1698431365
transform -1 0 14000 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__or2_4  _1311_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1312_
timestamp 1698431365
transform 1 0 11424 0 -1 26656
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1313_
timestamp 1698431365
transform -1 0 10192 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1314_
timestamp 1698431365
transform -1 0 6160 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1315_
timestamp 1698431365
transform 1 0 6272 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1316_
timestamp 1698431365
transform 1 0 12432 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1317_
timestamp 1698431365
transform -1 0 12768 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1318_
timestamp 1698431365
transform 1 0 2352 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _1319_
timestamp 1698431365
transform -1 0 3808 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1320_
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1321_
timestamp 1698431365
transform 1 0 6160 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1322_
timestamp 1698431365
transform -1 0 4592 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1323_
timestamp 1698431365
transform 1 0 3136 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1324_
timestamp 1698431365
transform 1 0 4816 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1325_
timestamp 1698431365
transform 1 0 6272 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1326_
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1327_
timestamp 1698431365
transform 1 0 7392 0 1 23520
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1328_
timestamp 1698431365
transform 1 0 4368 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _1329_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1330_
timestamp 1698431365
transform -1 0 9184 0 -1 26656
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1331_
timestamp 1698431365
transform -1 0 2576 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _1332_
timestamp 1698431365
transform -1 0 4480 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1333_
timestamp 1698431365
transform 1 0 6272 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1334_
timestamp 1698431365
transform 1 0 2576 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1335_
timestamp 1698431365
transform 1 0 7504 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _1336_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10080 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1337_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9968 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1338_
timestamp 1698431365
transform 1 0 28000 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1339_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1340_
timestamp 1698431365
transform 1 0 27888 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1341_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32592 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1342_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30128 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1343_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 21056 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1344_
timestamp 1698431365
transform 1 0 13552 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1345_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23632 0 -1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1346_
timestamp 1698431365
transform -1 0 28224 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1347_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32704 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1348_
timestamp 1698431365
transform -1 0 32704 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1349_
timestamp 1698431365
transform -1 0 31136 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1350_
timestamp 1698431365
transform 1 0 30688 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1351_
timestamp 1698431365
transform -1 0 25648 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1352_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32256 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1353_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31472 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1354_
timestamp 1698431365
transform 1 0 19936 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1355_
timestamp 1698431365
transform -1 0 11872 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1356_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16800 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1357_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13104 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1358_
timestamp 1698431365
transform -1 0 13104 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1359_
timestamp 1698431365
transform -1 0 18032 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1360_
timestamp 1698431365
transform 1 0 18704 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1361_
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1362_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18256 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1363_
timestamp 1698431365
transform 1 0 7168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1364_
timestamp 1698431365
transform 1 0 4368 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1365_
timestamp 1698431365
transform 1 0 6160 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1366_
timestamp 1698431365
transform -1 0 5264 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1367_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4480 0 -1 26656
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1368_
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1369_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7168 0 1 26656
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1370_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9856 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1371_
timestamp 1698431365
transform 1 0 31136 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1372_
timestamp 1698431365
transform -1 0 33152 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1373_
timestamp 1698431365
transform 1 0 31584 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1374_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31136 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1375_
timestamp 1698431365
transform 1 0 30240 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1376_
timestamp 1698431365
transform -1 0 10192 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1377_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6608 0 1 20384
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1378_
timestamp 1698431365
transform -1 0 18032 0 -1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1379_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13104 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1380_
timestamp 1698431365
transform 1 0 15344 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1381_
timestamp 1698431365
transform 1 0 17248 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1382_
timestamp 1698431365
transform 1 0 2240 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1383_
timestamp 1698431365
transform -1 0 2688 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1384_
timestamp 1698431365
transform -1 0 2576 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1385_
timestamp 1698431365
transform 1 0 6272 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1386_
timestamp 1698431365
transform -1 0 7168 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1387_
timestamp 1698431365
transform 1 0 5600 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1388_
timestamp 1698431365
transform -1 0 6832 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1389_
timestamp 1698431365
transform -1 0 5264 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1390_
timestamp 1698431365
transform 1 0 5936 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1391_
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1392_
timestamp 1698431365
transform -1 0 16352 0 -1 25088
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1393_
timestamp 1698431365
transform -1 0 10640 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1394_
timestamp 1698431365
transform -1 0 16240 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1395_
timestamp 1698431365
transform -1 0 12544 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1396_
timestamp 1698431365
transform -1 0 13328 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1397_
timestamp 1698431365
transform 1 0 13552 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1398_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12544 0 -1 29792
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1399_
timestamp 1698431365
transform 1 0 16128 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1400_
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1401_
timestamp 1698431365
transform 1 0 27328 0 -1 20384
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1402_
timestamp 1698431365
transform -1 0 26432 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1403_
timestamp 1698431365
transform 1 0 30800 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1404_
timestamp 1698431365
transform 1 0 26880 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1405_
timestamp 1698431365
transform -1 0 28784 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1406_
timestamp 1698431365
transform -1 0 30800 0 -1 23520
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1407_
timestamp 1698431365
transform 1 0 17472 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1408_
timestamp 1698431365
transform -1 0 22848 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1409_
timestamp 1698431365
transform -1 0 20944 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1410_
timestamp 1698431365
transform -1 0 20944 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1411_
timestamp 1698431365
transform -1 0 21728 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1412_
timestamp 1698431365
transform 1 0 21616 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1413_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20944 0 -1 29792
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1414_
timestamp 1698431365
transform 1 0 26880 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1415_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26096 0 1 31360
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1416_
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1417_
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1418_
timestamp 1698431365
transform -1 0 31024 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1419_
timestamp 1698431365
transform 1 0 26320 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1420_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28672 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1421_
timestamp 1698431365
transform -1 0 27328 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1422_
timestamp 1698431365
transform 1 0 27776 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1423_
timestamp 1698431365
transform 1 0 27888 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1424_
timestamp 1698431365
transform -1 0 28672 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1425_
timestamp 1698431365
transform -1 0 23632 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1426_
timestamp 1698431365
transform -1 0 27328 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1427_
timestamp 1698431365
transform -1 0 30128 0 -1 21952
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1428_
timestamp 1698431365
transform 1 0 19712 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1429_
timestamp 1698431365
transform 1 0 20160 0 1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1430_
timestamp 1698431365
transform -1 0 18816 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1431_
timestamp 1698431365
transform 1 0 19824 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1432_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19376 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1433_
timestamp 1698431365
transform 1 0 23408 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1434_
timestamp 1698431365
transform 1 0 4480 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1435_
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _1436_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4704 0 -1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1437_
timestamp 1698431365
transform -1 0 18704 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1438_
timestamp 1698431365
transform -1 0 13104 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1439_
timestamp 1698431365
transform 1 0 18032 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1440_
timestamp 1698431365
transform -1 0 17808 0 1 28224
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1441_
timestamp 1698431365
transform 1 0 13776 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1442_
timestamp 1698431365
transform -1 0 16912 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1443_
timestamp 1698431365
transform -1 0 13440 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1444_
timestamp 1698431365
transform 1 0 15120 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1445_
timestamp 1698431365
transform 1 0 23296 0 1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1446_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23968 0 1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1447_
timestamp 1698431365
transform 1 0 28336 0 -1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1448_
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1449_
timestamp 1698431365
transform 1 0 30128 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1450_
timestamp 1698431365
transform -1 0 26544 0 -1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1451_
timestamp 1698431365
transform -1 0 26208 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1452_
timestamp 1698431365
transform 1 0 23632 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1453_
timestamp 1698431365
transform 1 0 25312 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1454_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1455_
timestamp 1698431365
transform 1 0 20272 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1456_
timestamp 1698431365
transform 1 0 23072 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1457_
timestamp 1698431365
transform -1 0 28784 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1458_
timestamp 1698431365
transform 1 0 26432 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1459_
timestamp 1698431365
transform 1 0 26208 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1460_
timestamp 1698431365
transform -1 0 13440 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1461_
timestamp 1698431365
transform -1 0 9744 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1462_
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1463_
timestamp 1698431365
transform -1 0 16128 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1464_
timestamp 1698431365
transform 1 0 12096 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1465_
timestamp 1698431365
transform -1 0 9072 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1466_
timestamp 1698431365
transform 1 0 13440 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1467_
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1468_
timestamp 1698431365
transform 1 0 15680 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1469_
timestamp 1698431365
transform 1 0 27664 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1470_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 -1 34496
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1471_
timestamp 1698431365
transform 1 0 33152 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1472_
timestamp 1698431365
transform 1 0 34496 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1473_
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1474_
timestamp 1698431365
transform 1 0 30240 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1475_
timestamp 1698431365
transform -1 0 24864 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1476_
timestamp 1698431365
transform 1 0 26656 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1477_
timestamp 1698431365
transform 1 0 27552 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1478_
timestamp 1698431365
transform -1 0 28784 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1479_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20048 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1480_
timestamp 1698431365
transform 1 0 20944 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1481_
timestamp 1698431365
transform 1 0 23968 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1482_
timestamp 1698431365
transform -1 0 25760 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1483_
timestamp 1698431365
transform 1 0 22176 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1484_
timestamp 1698431365
transform 1 0 11424 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1485_
timestamp 1698431365
transform -1 0 17248 0 1 31360
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1486_
timestamp 1698431365
transform 1 0 19376 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1487_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11424 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1488_
timestamp 1698431365
transform -1 0 10304 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1489_
timestamp 1698431365
transform -1 0 5600 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1490_
timestamp 1698431365
transform -1 0 5264 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1491_
timestamp 1698431365
transform 1 0 7392 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1492_
timestamp 1698431365
transform 1 0 9184 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1493_
timestamp 1698431365
transform -1 0 12992 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1494_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14448 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1495_
timestamp 1698431365
transform 1 0 12992 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1496_
timestamp 1698431365
transform 1 0 22624 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1497_
timestamp 1698431365
transform 1 0 29792 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1498_
timestamp 1698431365
transform 1 0 30464 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1499_
timestamp 1698431365
transform -1 0 36288 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1500_
timestamp 1698431365
transform -1 0 24864 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1501_
timestamp 1698431365
transform -1 0 24864 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1502_
timestamp 1698431365
transform -1 0 23072 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1503_
timestamp 1698431365
transform 1 0 23632 0 1 23520
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1504_
timestamp 1698431365
transform -1 0 24864 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1505_
timestamp 1698431365
transform 1 0 22064 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1506_
timestamp 1698431365
transform 1 0 23184 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1507_
timestamp 1698431365
transform 1 0 24304 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1508_
timestamp 1698431365
transform 1 0 23968 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1509_
timestamp 1698431365
transform 1 0 24304 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1510_
timestamp 1698431365
transform -1 0 24304 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1511_
timestamp 1698431365
transform 1 0 22848 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1512_
timestamp 1698431365
transform -1 0 19152 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1513_
timestamp 1698431365
transform -1 0 19264 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1514_
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1515_
timestamp 1698431365
transform 1 0 16800 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1516_
timestamp 1698431365
transform 1 0 5824 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1517_
timestamp 1698431365
transform 1 0 4480 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1518_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11088 0 1 31360
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1519_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8960 0 -1 29792
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1520_
timestamp 1698431365
transform 1 0 7840 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1521_
timestamp 1698431365
transform 1 0 10752 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1522_
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1523_
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1524_
timestamp 1698431365
transform 1 0 23296 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1525_
timestamp 1698431365
transform -1 0 23184 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1526_
timestamp 1698431365
transform -1 0 24192 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1527_
timestamp 1698431365
transform 1 0 22064 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1528_
timestamp 1698431365
transform -1 0 24416 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1529_
timestamp 1698431365
transform 1 0 29456 0 -1 39200
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1530_
timestamp 1698431365
transform 1 0 29120 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1531_
timestamp 1698431365
transform -1 0 31696 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1532_
timestamp 1698431365
transform -1 0 32256 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1533_
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1534_
timestamp 1698431365
transform 1 0 37184 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1535_
timestamp 1698431365
transform 1 0 28784 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1536_
timestamp 1698431365
transform 1 0 33152 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1537_
timestamp 1698431365
transform 1 0 24192 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1538_
timestamp 1698431365
transform -1 0 22848 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1539_
timestamp 1698431365
transform 1 0 22736 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1540_
timestamp 1698431365
transform 1 0 22176 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1541_
timestamp 1698431365
transform 1 0 24752 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1542_
timestamp 1698431365
transform -1 0 6832 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1543_
timestamp 1698431365
transform -1 0 9072 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1544_
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1545_
timestamp 1698431365
transform 1 0 11536 0 1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1546_
timestamp 1698431365
transform 1 0 10864 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1547_
timestamp 1698431365
transform -1 0 9408 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1548_
timestamp 1698431365
transform -1 0 10528 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1549_
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1550_
timestamp 1698431365
transform 1 0 10976 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1551_
timestamp 1698431365
transform -1 0 9184 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1552_
timestamp 1698431365
transform 1 0 9184 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1553_
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1554_
timestamp 1698431365
transform -1 0 13776 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1555_
timestamp 1698431365
transform -1 0 13104 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1556_
timestamp 1698431365
transform 1 0 12656 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1557_
timestamp 1698431365
transform 1 0 23408 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1558_
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1559_
timestamp 1698431365
transform 1 0 19264 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1560_
timestamp 1698431365
transform 1 0 25984 0 1 25088
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1561_
timestamp 1698431365
transform 1 0 25648 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1562_
timestamp 1698431365
transform 1 0 28000 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1563_
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1564_
timestamp 1698431365
transform 1 0 29456 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1565_
timestamp 1698431365
transform -1 0 45136 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1566_
timestamp 1698431365
transform 1 0 31024 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1567_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30576 0 1 39200
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1568_
timestamp 1698431365
transform 1 0 30240 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1569_
timestamp 1698431365
transform 1 0 22736 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1570_
timestamp 1698431365
transform -1 0 26768 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1571_
timestamp 1698431365
transform -1 0 26096 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1572_
timestamp 1698431365
transform 1 0 27776 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1573_
timestamp 1698431365
transform -1 0 23968 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1574_
timestamp 1698431365
transform -1 0 25536 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1575_
timestamp 1698431365
transform -1 0 22848 0 1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1576_
timestamp 1698431365
transform 1 0 21616 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1577_
timestamp 1698431365
transform -1 0 22064 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1578_
timestamp 1698431365
transform 1 0 22064 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1579_
timestamp 1698431365
transform 1 0 22512 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1580_
timestamp 1698431365
transform 1 0 7168 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1581_
timestamp 1698431365
transform -1 0 10528 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1582_
timestamp 1698431365
transform -1 0 7392 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1583_
timestamp 1698431365
transform -1 0 9072 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1584_
timestamp 1698431365
transform -1 0 8400 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1585_
timestamp 1698431365
transform 1 0 8064 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1586_
timestamp 1698431365
transform -1 0 14560 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1587_
timestamp 1698431365
transform -1 0 11424 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1588_
timestamp 1698431365
transform 1 0 9632 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1589_
timestamp 1698431365
transform 1 0 9072 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1590_
timestamp 1698431365
transform 1 0 11536 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1591_
timestamp 1698431365
transform 1 0 11424 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1592_
timestamp 1698431365
transform 1 0 9296 0 1 42336
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1593_
timestamp 1698431365
transform 1 0 22512 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1594_
timestamp 1698431365
transform 1 0 29792 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1595_
timestamp 1698431365
transform 1 0 35056 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1596_
timestamp 1698431365
transform 1 0 35728 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1597_
timestamp 1698431365
transform 1 0 29120 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1598_
timestamp 1698431365
transform 1 0 31696 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1599_
timestamp 1698431365
transform 1 0 31136 0 1 42336
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1600_
timestamp 1698431365
transform -1 0 23520 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1601_
timestamp 1698431365
transform 1 0 27104 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1602_
timestamp 1698431365
transform -1 0 24976 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1603_
timestamp 1698431365
transform 1 0 23408 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1604_
timestamp 1698431365
transform -1 0 5264 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1605_
timestamp 1698431365
transform 1 0 12432 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1606_
timestamp 1698431365
transform 1 0 11424 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1607_
timestamp 1698431365
transform 1 0 12320 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1608_
timestamp 1698431365
transform 1 0 12432 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1609_
timestamp 1698431365
transform 1 0 13776 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1610_
timestamp 1698431365
transform -1 0 13888 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1611_
timestamp 1698431365
transform 1 0 9632 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1612_
timestamp 1698431365
transform -1 0 11872 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1613_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11424 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1614_
timestamp 1698431365
transform 1 0 10416 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1615_
timestamp 1698431365
transform 1 0 12320 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1616_
timestamp 1698431365
transform 1 0 23520 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1617_
timestamp 1698431365
transform 1 0 28560 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1618_
timestamp 1698431365
transform 1 0 31360 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1619_
timestamp 1698431365
transform 1 0 39088 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1620_
timestamp 1698431365
transform -1 0 24640 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1621_
timestamp 1698431365
transform -1 0 24640 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1622_
timestamp 1698431365
transform 1 0 24640 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1623_
timestamp 1698431365
transform 1 0 24192 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1624_
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1625_
timestamp 1698431365
transform 1 0 11872 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1626_
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1627_
timestamp 1698431365
transform -1 0 34384 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1628_
timestamp 1698431365
transform 1 0 29792 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1629_
timestamp 1698431365
transform 1 0 29904 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1630_
timestamp 1698431365
transform 1 0 31360 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1631_
timestamp 1698431365
transform 1 0 43680 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1632_
timestamp 1698431365
transform 1 0 32704 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1633_
timestamp 1698431365
transform -1 0 34384 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1634_
timestamp 1698431365
transform 1 0 39872 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1635_
timestamp 1698431365
transform -1 0 45136 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1636_
timestamp 1698431365
transform -1 0 47376 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1637_
timestamp 1698431365
transform -1 0 46704 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1638_
timestamp 1698431365
transform 1 0 43120 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1639_
timestamp 1698431365
transform -1 0 45024 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1640_
timestamp 1698431365
transform 1 0 15680 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1641_
timestamp 1698431365
transform -1 0 28896 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1642_
timestamp 1698431365
transform -1 0 26880 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1643_
timestamp 1698431365
transform -1 0 24192 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1644_
timestamp 1698431365
transform 1 0 11424 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1645_
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1646_
timestamp 1698431365
transform -1 0 23072 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1647_
timestamp 1698431365
transform 1 0 22736 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1648_
timestamp 1698431365
transform -1 0 17920 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1649_
timestamp 1698431365
transform -1 0 18368 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1650_
timestamp 1698431365
transform 1 0 18368 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1651_
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1652_
timestamp 1698431365
transform -1 0 29680 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1653_
timestamp 1698431365
transform 1 0 29344 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1654_
timestamp 1698431365
transform 1 0 16576 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1655_
timestamp 1698431365
transform -1 0 48160 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1656_
timestamp 1698431365
transform -1 0 20384 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1657_
timestamp 1698431365
transform 1 0 19376 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1658_
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1659_
timestamp 1698431365
transform -1 0 14784 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1660_
timestamp 1698431365
transform -1 0 23520 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1661_
timestamp 1698431365
transform 1 0 17360 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1662_
timestamp 1698431365
transform -1 0 16128 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1663_
timestamp 1698431365
transform -1 0 34720 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1664_
timestamp 1698431365
transform -1 0 30576 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1665_
timestamp 1698431365
transform -1 0 17024 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1666_
timestamp 1698431365
transform 1 0 18144 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1667_
timestamp 1698431365
transform -1 0 48048 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1668_
timestamp 1698431365
transform -1 0 25984 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1669_
timestamp 1698431365
transform -1 0 18144 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1670_
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1671_
timestamp 1698431365
transform -1 0 30576 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1672_
timestamp 1698431365
transform -1 0 28784 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1673_
timestamp 1698431365
transform 1 0 26768 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1674_
timestamp 1698431365
transform -1 0 27216 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1675_
timestamp 1698431365
transform 1 0 27664 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1676_
timestamp 1698431365
transform 1 0 26768 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1677_
timestamp 1698431365
transform 1 0 27328 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1678_
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1679_
timestamp 1698431365
transform -1 0 28784 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1680_
timestamp 1698431365
transform 1 0 26992 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1681_
timestamp 1698431365
transform 1 0 28000 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1682_
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1683_
timestamp 1698431365
transform 1 0 28784 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1684_
timestamp 1698431365
transform 1 0 27216 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1685_
timestamp 1698431365
transform 1 0 26432 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1686_
timestamp 1698431365
transform -1 0 34384 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1687_
timestamp 1698431365
transform 1 0 23296 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1688_
timestamp 1698431365
transform 1 0 27328 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1689_
timestamp 1698431365
transform 1 0 27440 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1690_
timestamp 1698431365
transform 1 0 28112 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1691_
timestamp 1698431365
transform -1 0 32368 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1692_
timestamp 1698431365
transform -1 0 31808 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1693_
timestamp 1698431365
transform 1 0 30464 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1694_
timestamp 1698431365
transform 1 0 29344 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1695_
timestamp 1698431365
transform -1 0 32256 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1696_
timestamp 1698431365
transform 1 0 30464 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1697_
timestamp 1698431365
transform 1 0 22512 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1698_
timestamp 1698431365
transform 1 0 18144 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1699_
timestamp 1698431365
transform -1 0 32368 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1700_
timestamp 1698431365
transform 1 0 31584 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1701_
timestamp 1698431365
transform -1 0 33824 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1702_
timestamp 1698431365
transform -1 0 33824 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1703_
timestamp 1698431365
transform -1 0 44240 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1704_
timestamp 1698431365
transform -1 0 43008 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1705_
timestamp 1698431365
transform -1 0 35952 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1706_
timestamp 1698431365
transform -1 0 34384 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1707_
timestamp 1698431365
transform 1 0 31472 0 1 25088
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1708_
timestamp 1698431365
transform 1 0 34832 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1709_
timestamp 1698431365
transform -1 0 35280 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1710_
timestamp 1698431365
transform -1 0 35728 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1711_
timestamp 1698431365
transform -1 0 34608 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1712_
timestamp 1698431365
transform 1 0 25200 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1713_
timestamp 1698431365
transform 1 0 26208 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1714_
timestamp 1698431365
transform 1 0 26432 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1715_
timestamp 1698431365
transform -1 0 42112 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1716_
timestamp 1698431365
transform -1 0 39984 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1717_
timestamp 1698431365
transform -1 0 22512 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1718_
timestamp 1698431365
transform -1 0 26544 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1719_
timestamp 1698431365
transform 1 0 25536 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1720_
timestamp 1698431365
transform -1 0 25984 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1721_
timestamp 1698431365
transform -1 0 23968 0 1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1722_
timestamp 1698431365
transform -1 0 21840 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1723_
timestamp 1698431365
transform -1 0 23632 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1724_
timestamp 1698431365
transform 1 0 20384 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1725_
timestamp 1698431365
transform 1 0 21280 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1726_
timestamp 1698431365
transform -1 0 20944 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1727_
timestamp 1698431365
transform 1 0 18592 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1728_
timestamp 1698431365
transform -1 0 18256 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1729_
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1730_
timestamp 1698431365
transform -1 0 19936 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1731_
timestamp 1698431365
transform 1 0 19264 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1732_
timestamp 1698431365
transform 1 0 19040 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1733_
timestamp 1698431365
transform -1 0 21840 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1734_
timestamp 1698431365
transform -1 0 22960 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1735_
timestamp 1698431365
transform -1 0 19040 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1736_
timestamp 1698431365
transform -1 0 19376 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1737_
timestamp 1698431365
transform 1 0 18928 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1738_
timestamp 1698431365
transform -1 0 20832 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1739_
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1740_
timestamp 1698431365
transform 1 0 19488 0 -1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1741_
timestamp 1698431365
transform -1 0 21840 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1742_
timestamp 1698431365
transform 1 0 19936 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1743_
timestamp 1698431365
transform 1 0 21504 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1744_
timestamp 1698431365
transform 1 0 20608 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1745_
timestamp 1698431365
transform -1 0 23968 0 -1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1746_
timestamp 1698431365
transform -1 0 21952 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1747_
timestamp 1698431365
transform -1 0 20944 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1748_
timestamp 1698431365
transform -1 0 22512 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1749_
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1750_
timestamp 1698431365
transform 1 0 18816 0 -1 42336
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1751_
timestamp 1698431365
transform -1 0 21392 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1752_
timestamp 1698431365
transform 1 0 11424 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1753_
timestamp 1698431365
transform -1 0 21616 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1754_
timestamp 1698431365
transform 1 0 17248 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1755_
timestamp 1698431365
transform -1 0 19600 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1756_
timestamp 1698431365
transform 1 0 17920 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1757_
timestamp 1698431365
transform -1 0 19712 0 1 39200
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1758_
timestamp 1698431365
transform -1 0 15792 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1759_
timestamp 1698431365
transform 1 0 16464 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1760_
timestamp 1698431365
transform -1 0 18144 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1761_
timestamp 1698431365
transform -1 0 18144 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1762_
timestamp 1698431365
transform 1 0 8176 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1763_
timestamp 1698431365
transform 1 0 11312 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1764_
timestamp 1698431365
transform 1 0 9184 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1765_
timestamp 1698431365
transform 1 0 8624 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1766_
timestamp 1698431365
transform 1 0 9632 0 -1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1767_
timestamp 1698431365
transform -1 0 11424 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1768_
timestamp 1698431365
transform 1 0 9632 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1769_
timestamp 1698431365
transform 1 0 7616 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1770_
timestamp 1698431365
transform 1 0 10304 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1771_
timestamp 1698431365
transform -1 0 15568 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1772_
timestamp 1698431365
transform 1 0 13440 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1773_
timestamp 1698431365
transform 1 0 14000 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1774_
timestamp 1698431365
transform 1 0 14560 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1775_
timestamp 1698431365
transform -1 0 15568 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1776_
timestamp 1698431365
transform -1 0 17696 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1777_
timestamp 1698431365
transform -1 0 17024 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1778_
timestamp 1698431365
transform 1 0 14112 0 -1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1779_
timestamp 1698431365
transform -1 0 16912 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1780_
timestamp 1698431365
transform 1 0 14560 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1781_
timestamp 1698431365
transform 1 0 14112 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1782_
timestamp 1698431365
transform 1 0 15344 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1783_
timestamp 1698431365
transform -1 0 16240 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1784_
timestamp 1698431365
transform 1 0 9520 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1785_
timestamp 1698431365
transform 1 0 11760 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1786_
timestamp 1698431365
transform 1 0 11872 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1787_
timestamp 1698431365
transform -1 0 10864 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1788_
timestamp 1698431365
transform 1 0 10192 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1789_
timestamp 1698431365
transform 1 0 10192 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1790_
timestamp 1698431365
transform 1 0 3360 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1791_
timestamp 1698431365
transform -1 0 5264 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1792_
timestamp 1698431365
transform -1 0 5712 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1793_
timestamp 1698431365
transform 1 0 5712 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1794_
timestamp 1698431365
transform -1 0 5264 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1795_
timestamp 1698431365
transform 1 0 3920 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1796_
timestamp 1698431365
transform -1 0 3920 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1797_
timestamp 1698431365
transform -1 0 3696 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1798_
timestamp 1698431365
transform 1 0 3024 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1799_
timestamp 1698431365
transform 1 0 2128 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1800_
timestamp 1698431365
transform 1 0 39984 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1801_
timestamp 1698431365
transform -1 0 14336 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1802_
timestamp 1698431365
transform -1 0 5152 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1803_
timestamp 1698431365
transform -1 0 4592 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1804_
timestamp 1698431365
transform -1 0 4816 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1805_
timestamp 1698431365
transform 1 0 1680 0 1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1806_
timestamp 1698431365
transform 1 0 4256 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1807_
timestamp 1698431365
transform 1 0 2688 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1808_
timestamp 1698431365
transform -1 0 6608 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1809_
timestamp 1698431365
transform -1 0 5040 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1810_
timestamp 1698431365
transform 1 0 6048 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1811_
timestamp 1698431365
transform -1 0 6048 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1812_
timestamp 1698431365
transform 1 0 3136 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1813_
timestamp 1698431365
transform 1 0 2800 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1814_
timestamp 1698431365
transform -1 0 6048 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1815_
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1816_
timestamp 1698431365
transform -1 0 6944 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1817_
timestamp 1698431365
transform 1 0 13888 0 1 42336
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1818_
timestamp 1698431365
transform -1 0 16240 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1819_
timestamp 1698431365
transform 1 0 15120 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1820_
timestamp 1698431365
transform -1 0 29904 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1821_
timestamp 1698431365
transform 1 0 32480 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1822_
timestamp 1698431365
transform 1 0 16016 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1823_
timestamp 1698431365
transform -1 0 15120 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1824_
timestamp 1698431365
transform -1 0 5264 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1825_
timestamp 1698431365
transform 1 0 1792 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1826_
timestamp 1698431365
transform -1 0 2688 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1827_
timestamp 1698431365
transform -1 0 4256 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1828_
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1829_
timestamp 1698431365
transform 1 0 3696 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1830_
timestamp 1698431365
transform -1 0 2240 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1831_
timestamp 1698431365
transform 1 0 2128 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1832_
timestamp 1698431365
transform 1 0 2800 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1833_
timestamp 1698431365
transform 1 0 2240 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1834_
timestamp 1698431365
transform -1 0 7392 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1835_
timestamp 1698431365
transform 1 0 3584 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1836_
timestamp 1698431365
transform -1 0 2688 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1837_
timestamp 1698431365
transform -1 0 4144 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1838_
timestamp 1698431365
transform 1 0 2688 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1839_
timestamp 1698431365
transform 1 0 2688 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1840_
timestamp 1698431365
transform -1 0 8064 0 1 31360
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1841_
timestamp 1698431365
transform 1 0 6944 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1842_
timestamp 1698431365
transform -1 0 6272 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1843_
timestamp 1698431365
transform -1 0 6832 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1844_
timestamp 1698431365
transform -1 0 5936 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1845_
timestamp 1698431365
transform 1 0 4256 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1846_
timestamp 1698431365
transform -1 0 6160 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1847_
timestamp 1698431365
transform 1 0 2800 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1848_
timestamp 1698431365
transform 1 0 2464 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1849_
timestamp 1698431365
transform -1 0 7392 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1850_
timestamp 1698431365
transform -1 0 6944 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1851_
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1852_
timestamp 1698431365
transform 1 0 5936 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1853_
timestamp 1698431365
transform 1 0 7280 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1854_
timestamp 1698431365
transform 1 0 6160 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1855_
timestamp 1698431365
transform -1 0 6160 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1856_
timestamp 1698431365
transform 1 0 7056 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1857_
timestamp 1698431365
transform -1 0 7168 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1858_
timestamp 1698431365
transform -1 0 7616 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1859_
timestamp 1698431365
transform 1 0 6272 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1860_
timestamp 1698431365
transform -1 0 6272 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1861_
timestamp 1698431365
transform -1 0 41104 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1862_
timestamp 1698431365
transform 1 0 6720 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1863_
timestamp 1698431365
transform -1 0 8512 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1864_
timestamp 1698431365
transform 1 0 7280 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1865_
timestamp 1698431365
transform 1 0 6496 0 1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1866_
timestamp 1698431365
transform -1 0 9072 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1867_
timestamp 1698431365
transform 1 0 7392 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1868_
timestamp 1698431365
transform 1 0 6832 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1869_
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1870_
timestamp 1698431365
transform 1 0 6720 0 1 43904
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1871_
timestamp 1698431365
transform 1 0 9184 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1872_
timestamp 1698431365
transform 1 0 7056 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1873_
timestamp 1698431365
transform -1 0 9856 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1874_
timestamp 1698431365
transform -1 0 8624 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1875_
timestamp 1698431365
transform 1 0 7504 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1876_
timestamp 1698431365
transform -1 0 13104 0 1 43904
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1877_
timestamp 1698431365
transform -1 0 10528 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1878_
timestamp 1698431365
transform 1 0 12320 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1879_
timestamp 1698431365
transform 1 0 10416 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1880_
timestamp 1698431365
transform -1 0 32144 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1881_
timestamp 1698431365
transform 1 0 12880 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1882_
timestamp 1698431365
transform 1 0 12656 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1883_
timestamp 1698431365
transform 1 0 45360 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1884_
timestamp 1698431365
transform 1 0 39984 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1885_
timestamp 1698431365
transform 1 0 42000 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1886_
timestamp 1698431365
transform -1 0 44128 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1887_
timestamp 1698431365
transform -1 0 43120 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1888_
timestamp 1698431365
transform 1 0 41440 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1889_
timestamp 1698431365
transform 1 0 46144 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1890_
timestamp 1698431365
transform 1 0 46144 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1891_
timestamp 1698431365
transform 1 0 45248 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1892_
timestamp 1698431365
transform -1 0 45360 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1893_
timestamp 1698431365
transform -1 0 47712 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1894_
timestamp 1698431365
transform 1 0 47040 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1895_
timestamp 1698431365
transform 1 0 39872 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1896_
timestamp 1698431365
transform -1 0 46816 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1897_
timestamp 1698431365
transform -1 0 43680 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1898_
timestamp 1698431365
transform 1 0 44800 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1899_
timestamp 1698431365
transform -1 0 29232 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1900_
timestamp 1698431365
transform 1 0 43120 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1901_
timestamp 1698431365
transform -1 0 46480 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1902_
timestamp 1698431365
transform 1 0 43792 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1903_
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1904_
timestamp 1698431365
transform 1 0 42448 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1905_
timestamp 1698431365
transform 1 0 44016 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1906_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33040 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1907_
timestamp 1698431365
transform 1 0 41552 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1908_
timestamp 1698431365
transform 1 0 43568 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1909_
timestamp 1698431365
transform -1 0 45024 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1910_
timestamp 1698431365
transform -1 0 43008 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1911_
timestamp 1698431365
transform -1 0 44352 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1912_
timestamp 1698431365
transform 1 0 41440 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1913_
timestamp 1698431365
transform 1 0 43008 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1914_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42672 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1915_
timestamp 1698431365
transform -1 0 41440 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1916_
timestamp 1698431365
transform -1 0 45920 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1917_
timestamp 1698431365
transform 1 0 44128 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1918_
timestamp 1698431365
transform -1 0 45360 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1919_
timestamp 1698431365
transform 1 0 43792 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1920_
timestamp 1698431365
transform 1 0 43344 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1921_
timestamp 1698431365
transform 1 0 44800 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1922_
timestamp 1698431365
transform 1 0 43568 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1923_
timestamp 1698431365
transform 1 0 44240 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1924_
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1925_
timestamp 1698431365
transform 1 0 47376 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1926_
timestamp 1698431365
transform 1 0 45920 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1927_
timestamp 1698431365
transform 1 0 46480 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1928_
timestamp 1698431365
transform 1 0 47376 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1929_
timestamp 1698431365
transform 1 0 47152 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1930_
timestamp 1698431365
transform -1 0 47376 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1931_
timestamp 1698431365
transform -1 0 47152 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1932_
timestamp 1698431365
transform 1 0 43792 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1933_
timestamp 1698431365
transform 1 0 47152 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1934_
timestamp 1698431365
transform 1 0 45360 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1935_
timestamp 1698431365
transform -1 0 47152 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1936_
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1937_
timestamp 1698431365
transform -1 0 47488 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1938_
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1939_
timestamp 1698431365
transform 1 0 46032 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1940_
timestamp 1698431365
transform -1 0 46704 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1941_
timestamp 1698431365
transform -1 0 46256 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1942_
timestamp 1698431365
transform 1 0 45248 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1943_
timestamp 1698431365
transform -1 0 47824 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1944_
timestamp 1698431365
transform 1 0 46704 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1945_
timestamp 1698431365
transform -1 0 47264 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1946_
timestamp 1698431365
transform 1 0 47376 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1947_
timestamp 1698431365
transform 1 0 44912 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1948_
timestamp 1698431365
transform 1 0 47824 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1949_
timestamp 1698431365
transform 1 0 45696 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1950_
timestamp 1698431365
transform -1 0 47376 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1951_
timestamp 1698431365
transform 1 0 45024 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1952_
timestamp 1698431365
transform 1 0 47264 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1953_
timestamp 1698431365
transform 1 0 46704 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1954_
timestamp 1698431365
transform 1 0 47264 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1955_
timestamp 1698431365
transform 1 0 47600 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1956_
timestamp 1698431365
transform -1 0 47264 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1957_
timestamp 1698431365
transform 1 0 46592 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1958_
timestamp 1698431365
transform -1 0 47040 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1959_
timestamp 1698431365
transform 1 0 46144 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1960_
timestamp 1698431365
transform -1 0 46592 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1961_
timestamp 1698431365
transform -1 0 46144 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1962_
timestamp 1698431365
transform -1 0 44016 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1963_
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1964_
timestamp 1698431365
transform -1 0 39200 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1965_
timestamp 1698431365
transform 1 0 39200 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1966_
timestamp 1698431365
transform 1 0 42448 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1967_
timestamp 1698431365
transform 1 0 41552 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1968_
timestamp 1698431365
transform -1 0 48160 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1969_
timestamp 1698431365
transform 1 0 45360 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1970_
timestamp 1698431365
transform 1 0 46480 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1971_
timestamp 1698431365
transform 1 0 47040 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1972_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 48384 0 -1 26656
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1973_
timestamp 1698431365
transform -1 0 48384 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1974_
timestamp 1698431365
transform -1 0 41328 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1975_
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1976_
timestamp 1698431365
transform -1 0 42000 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1977_
timestamp 1698431365
transform 1 0 40656 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1978_
timestamp 1698431365
transform 1 0 47152 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1979_
timestamp 1698431365
transform 1 0 46816 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1980_
timestamp 1698431365
transform -1 0 37520 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1981_
timestamp 1698431365
transform -1 0 14560 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1982_
timestamp 1698431365
transform 1 0 25312 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1983_
timestamp 1698431365
transform 1 0 33152 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1984_
timestamp 1698431365
transform 1 0 39088 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1985_
timestamp 1698431365
transform 1 0 38752 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1986_
timestamp 1698431365
transform 1 0 39536 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1987_
timestamp 1698431365
transform -1 0 39088 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1988_
timestamp 1698431365
transform 1 0 39536 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1989_
timestamp 1698431365
transform -1 0 38304 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1990_
timestamp 1698431365
transform 1 0 39536 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1991_
timestamp 1698431365
transform 1 0 37744 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1992_
timestamp 1698431365
transform -1 0 39312 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1993_
timestamp 1698431365
transform 1 0 35952 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1994_
timestamp 1698431365
transform -1 0 38528 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1995_
timestamp 1698431365
transform -1 0 37744 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1996_
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1997_
timestamp 1698431365
transform -1 0 36624 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1998_
timestamp 1698431365
transform -1 0 38080 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1999_
timestamp 1698431365
transform -1 0 38640 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2000_
timestamp 1698431365
transform -1 0 38752 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2001_
timestamp 1698431365
transform 1 0 40320 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2002_
timestamp 1698431365
transform -1 0 39424 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2003_
timestamp 1698431365
transform 1 0 38640 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2004_
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2005_
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2006_
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2007_
timestamp 1698431365
transform 1 0 37744 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2008_
timestamp 1698431365
transform -1 0 39760 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2009_
timestamp 1698431365
transform 1 0 34272 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2010_
timestamp 1698431365
transform -1 0 38640 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2011_
timestamp 1698431365
transform -1 0 39200 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2012_
timestamp 1698431365
transform -1 0 38304 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2013_
timestamp 1698431365
transform -1 0 37968 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2014_
timestamp 1698431365
transform -1 0 37296 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2015_
timestamp 1698431365
transform 1 0 34272 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2016_
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2017_
timestamp 1698431365
transform 1 0 35168 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2018_
timestamp 1698431365
transform 1 0 34272 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2019_
timestamp 1698431365
transform 1 0 34048 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2020_
timestamp 1698431365
transform 1 0 34608 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2021_
timestamp 1698431365
transform 1 0 35616 0 -1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2022_
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2023_
timestamp 1698431365
transform -1 0 34944 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2024_
timestamp 1698431365
transform 1 0 33600 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2025_
timestamp 1698431365
transform -1 0 33376 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2026_
timestamp 1698431365
transform -1 0 32704 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2027_
timestamp 1698431365
transform -1 0 34608 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2028_
timestamp 1698431365
transform 1 0 31024 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2029_
timestamp 1698431365
transform -1 0 33152 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2030_
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2031_
timestamp 1698431365
transform 1 0 31696 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2032_
timestamp 1698431365
transform 1 0 29904 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2033_
timestamp 1698431365
transform 1 0 30240 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2034_
timestamp 1698431365
transform 1 0 25872 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2035_
timestamp 1698431365
transform -1 0 34272 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2036_
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2037_
timestamp 1698431365
transform 1 0 26992 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2038_
timestamp 1698431365
transform 1 0 26096 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2039_
timestamp 1698431365
transform 1 0 27216 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2040_
timestamp 1698431365
transform 1 0 27888 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2041_
timestamp 1698431365
transform 1 0 25424 0 1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2042_
timestamp 1698431365
transform 1 0 28000 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2043_
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2044_
timestamp 1698431365
transform -1 0 28000 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2045_
timestamp 1698431365
transform -1 0 27440 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2046_
timestamp 1698431365
transform 1 0 25984 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2047_
timestamp 1698431365
transform 1 0 26880 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2048_
timestamp 1698431365
transform -1 0 28224 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2049_
timestamp 1698431365
transform 1 0 25984 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2050_
timestamp 1698431365
transform 1 0 26544 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2051_
timestamp 1698431365
transform 1 0 25984 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2052_
timestamp 1698431365
transform 1 0 26656 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2053_
timestamp 1698431365
transform 1 0 27664 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2054_
timestamp 1698431365
transform 1 0 27552 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2055_
timestamp 1698431365
transform -1 0 28560 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2056_
timestamp 1698431365
transform 1 0 26320 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2057_
timestamp 1698431365
transform -1 0 25760 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2058_
timestamp 1698431365
transform 1 0 23520 0 1 43904
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2059_
timestamp 1698431365
transform 1 0 25872 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2060_
timestamp 1698431365
transform 1 0 24192 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2061_
timestamp 1698431365
transform -1 0 25872 0 -1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2062_
timestamp 1698431365
transform -1 0 24752 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2063_
timestamp 1698431365
transform -1 0 21616 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2064_
timestamp 1698431365
transform -1 0 42224 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2065_
timestamp 1698431365
transform 1 0 42224 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2066_
timestamp 1698431365
transform -1 0 33152 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2067_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 43680 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2068_
timestamp 1698431365
transform 1 0 37408 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2069_
timestamp 1698431365
transform -1 0 42336 0 1 9408
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2070_
timestamp 1698431365
transform -1 0 42224 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2071_
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2072_
timestamp 1698431365
transform 1 0 42112 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2073_
timestamp 1698431365
transform -1 0 15344 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2074_
timestamp 1698431365
transform 1 0 37296 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2075_
timestamp 1698431365
transform 1 0 39648 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2076_
timestamp 1698431365
transform 1 0 42112 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2077_
timestamp 1698431365
transform 1 0 31472 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2078_
timestamp 1698431365
transform 1 0 33600 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2079_
timestamp 1698431365
transform -1 0 40544 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2080_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40768 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2081_
timestamp 1698431365
transform 1 0 42336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2082_
timestamp 1698431365
transform 1 0 39648 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2083_
timestamp 1698431365
transform -1 0 38192 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2084_
timestamp 1698431365
transform 1 0 43008 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2085_
timestamp 1698431365
transform -1 0 42112 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2086_
timestamp 1698431365
transform 1 0 40992 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2087_
timestamp 1698431365
transform -1 0 39424 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2088_
timestamp 1698431365
transform 1 0 38416 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2089_
timestamp 1698431365
transform -1 0 39984 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2090_
timestamp 1698431365
transform -1 0 39088 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2091_
timestamp 1698431365
transform 1 0 34272 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2092_
timestamp 1698431365
transform 1 0 39312 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2093_
timestamp 1698431365
transform 1 0 39424 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2094_
timestamp 1698431365
transform 1 0 37520 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2095_
timestamp 1698431365
transform -1 0 38528 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2096_
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2097_
timestamp 1698431365
transform 1 0 38528 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2098_
timestamp 1698431365
transform 1 0 37968 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2099_
timestamp 1698431365
transform 1 0 39424 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2100_
timestamp 1698431365
transform -1 0 34608 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2101_
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2102_
timestamp 1698431365
transform -1 0 36624 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2103_
timestamp 1698431365
transform 1 0 36624 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2104_
timestamp 1698431365
transform 1 0 35616 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2105_
timestamp 1698431365
transform -1 0 37296 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2106_
timestamp 1698431365
transform -1 0 36736 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2107_
timestamp 1698431365
transform 1 0 35168 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2108_
timestamp 1698431365
transform 1 0 35056 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2109_
timestamp 1698431365
transform 1 0 36064 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2110_
timestamp 1698431365
transform -1 0 36064 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2111_
timestamp 1698431365
transform 1 0 35168 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2112_
timestamp 1698431365
transform 1 0 35840 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2113_
timestamp 1698431365
transform -1 0 37744 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2114_
timestamp 1698431365
transform -1 0 36512 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2115_
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2116_
timestamp 1698431365
transform 1 0 35056 0 1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2117_
timestamp 1698431365
transform 1 0 34384 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2118_
timestamp 1698431365
transform 1 0 34608 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2119_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35504 0 -1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2120_
timestamp 1698431365
transform 1 0 33824 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2121_
timestamp 1698431365
transform -1 0 33824 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2122_
timestamp 1698431365
transform -1 0 34608 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2123_
timestamp 1698431365
transform 1 0 33824 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2124_
timestamp 1698431365
transform -1 0 35616 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2125_
timestamp 1698431365
transform -1 0 35616 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2126_
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2127_
timestamp 1698431365
transform 1 0 33824 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2128_
timestamp 1698431365
transform 1 0 33600 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2129_
timestamp 1698431365
transform 1 0 35056 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2130_
timestamp 1698431365
transform -1 0 33824 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2131_
timestamp 1698431365
transform -1 0 33824 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2132_
timestamp 1698431365
transform 1 0 34048 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2133_
timestamp 1698431365
transform -1 0 31248 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2134_
timestamp 1698431365
transform 1 0 21840 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2135_
timestamp 1698431365
transform -1 0 27664 0 1 7840
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2136_
timestamp 1698431365
transform -1 0 32592 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2137_
timestamp 1698431365
transform 1 0 34944 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2138_
timestamp 1698431365
transform 1 0 34048 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2139_
timestamp 1698431365
transform 1 0 30128 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2140_
timestamp 1698431365
transform 1 0 31136 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2141_
timestamp 1698431365
transform 1 0 32928 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2142_
timestamp 1698431365
transform 1 0 22848 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2143_
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2144_
timestamp 1698431365
transform 1 0 34944 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2145_
timestamp 1698431365
transform -1 0 32144 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2146_
timestamp 1698431365
transform 1 0 32032 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2147_
timestamp 1698431365
transform 1 0 31584 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2148_
timestamp 1698431365
transform 1 0 33600 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2149_
timestamp 1698431365
transform -1 0 31584 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2150_
timestamp 1698431365
transform 1 0 23296 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2151_
timestamp 1698431365
transform -1 0 24752 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2152_
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2153_
timestamp 1698431365
transform -1 0 24192 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2154_
timestamp 1698431365
transform -1 0 26656 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2155_
timestamp 1698431365
transform 1 0 23968 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2156_
timestamp 1698431365
transform 1 0 24192 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2157_
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2158_
timestamp 1698431365
transform 1 0 21728 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2159_
timestamp 1698431365
transform -1 0 21952 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2160_
timestamp 1698431365
transform 1 0 21952 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2161_
timestamp 1698431365
transform 1 0 21952 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2162_
timestamp 1698431365
transform -1 0 22400 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2163_
timestamp 1698431365
transform -1 0 20272 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2164_
timestamp 1698431365
transform -1 0 20384 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2165_
timestamp 1698431365
transform -1 0 19488 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2166_
timestamp 1698431365
transform -1 0 20944 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2167_
timestamp 1698431365
transform 1 0 19488 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2168_
timestamp 1698431365
transform -1 0 19824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2169_
timestamp 1698431365
transform 1 0 19936 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2170_
timestamp 1698431365
transform 1 0 21616 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2171_
timestamp 1698431365
transform 1 0 19488 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2172_
timestamp 1698431365
transform 1 0 19376 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2173_
timestamp 1698431365
transform -1 0 21728 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2174_
timestamp 1698431365
transform 1 0 20160 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2175_
timestamp 1698431365
transform 1 0 18928 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2176_
timestamp 1698431365
transform 1 0 23072 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2177_
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2178_
timestamp 1698431365
transform -1 0 22960 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2179_
timestamp 1698431365
transform 1 0 22960 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2180_
timestamp 1698431365
transform -1 0 21392 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2181_
timestamp 1698431365
transform 1 0 22960 0 -1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2182_
timestamp 1698431365
transform 1 0 21280 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2183_
timestamp 1698431365
transform 1 0 23072 0 -1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2184_
timestamp 1698431365
transform -1 0 22960 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2185_
timestamp 1698431365
transform 1 0 21504 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2186_
timestamp 1698431365
transform 1 0 22400 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2187_
timestamp 1698431365
transform -1 0 39872 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2188_
timestamp 1698431365
transform 1 0 22176 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2189_
timestamp 1698431365
transform 1 0 21616 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2190_
timestamp 1698431365
transform 1 0 21728 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2191_
timestamp 1698431365
transform 1 0 23184 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2192_
timestamp 1698431365
transform 1 0 30688 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2193_
timestamp 1698431365
transform 1 0 3360 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2194_
timestamp 1698431365
transform 1 0 2464 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2195_
timestamp 1698431365
transform 1 0 13664 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2196_
timestamp 1698431365
transform 1 0 10864 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2197_
timestamp 1698431365
transform 1 0 8512 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2198_
timestamp 1698431365
transform 1 0 10528 0 -1 7840
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2199_
timestamp 1698431365
transform 1 0 11648 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2200_
timestamp 1698431365
transform 1 0 14784 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2201_
timestamp 1698431365
transform -1 0 14784 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2202_
timestamp 1698431365
transform -1 0 14000 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2203_
timestamp 1698431365
transform 1 0 14224 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2204_
timestamp 1698431365
transform -1 0 13328 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2205_
timestamp 1698431365
transform 1 0 13328 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2206_
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2207_
timestamp 1698431365
transform -1 0 13440 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2208_
timestamp 1698431365
transform -1 0 12768 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2209_
timestamp 1698431365
transform -1 0 10864 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2210_
timestamp 1698431365
transform -1 0 11648 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2211_
timestamp 1698431365
transform -1 0 10416 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2212_
timestamp 1698431365
transform 1 0 10416 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2213_
timestamp 1698431365
transform -1 0 10528 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2214_
timestamp 1698431365
transform -1 0 10528 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2215_
timestamp 1698431365
transform 1 0 9072 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2216_
timestamp 1698431365
transform -1 0 7840 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2217_
timestamp 1698431365
transform 1 0 8176 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2218_
timestamp 1698431365
transform -1 0 10976 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2219_
timestamp 1698431365
transform 1 0 7840 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2220_
timestamp 1698431365
transform -1 0 7840 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2221_
timestamp 1698431365
transform -1 0 7504 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2222_
timestamp 1698431365
transform 1 0 6272 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2223_
timestamp 1698431365
transform -1 0 6608 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2224_
timestamp 1698431365
transform 1 0 7168 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2225_
timestamp 1698431365
transform -1 0 5936 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2226_
timestamp 1698431365
transform -1 0 7392 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2227_
timestamp 1698431365
transform 1 0 7392 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2228_
timestamp 1698431365
transform -1 0 7168 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2229_
timestamp 1698431365
transform 1 0 7168 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2230_
timestamp 1698431365
transform -1 0 5936 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2231_
timestamp 1698431365
transform -1 0 10192 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2232_
timestamp 1698431365
transform -1 0 8064 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2233_
timestamp 1698431365
transform -1 0 7728 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2234_
timestamp 1698431365
transform 1 0 8064 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2235_
timestamp 1698431365
transform -1 0 9520 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2236_
timestamp 1698431365
transform -1 0 9072 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2237_
timestamp 1698431365
transform -1 0 5152 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2238_
timestamp 1698431365
transform -1 0 13104 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2239_
timestamp 1698431365
transform 1 0 7392 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2240_
timestamp 1698431365
transform -1 0 10752 0 1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2241_
timestamp 1698431365
transform 1 0 10976 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2242_
timestamp 1698431365
transform -1 0 9184 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2243_
timestamp 1698431365
transform 1 0 11648 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2244_
timestamp 1698431365
transform 1 0 10192 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2245_
timestamp 1698431365
transform -1 0 11872 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2246_
timestamp 1698431365
transform 1 0 12768 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2247_
timestamp 1698431365
transform 1 0 11872 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2248_
timestamp 1698431365
transform 1 0 11872 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2249_
timestamp 1698431365
transform -1 0 10416 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2250_
timestamp 1698431365
transform -1 0 9744 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2251_
timestamp 1698431365
transform 1 0 10640 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2252_
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2253_
timestamp 1698431365
transform 1 0 9520 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2254_
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2255_
timestamp 1698431365
transform 1 0 32592 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2256_
timestamp 1698431365
transform 1 0 38192 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2257_
timestamp 1698431365
transform 1 0 37072 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2258_
timestamp 1698431365
transform -1 0 40096 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2259_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28000 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2260_
timestamp 1698431365
transform -1 0 31136 0 1 28224
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2261_
timestamp 1698431365
transform 1 0 29456 0 -1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2262_
timestamp 1698431365
transform -1 0 40544 0 -1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2263_
timestamp 1698431365
transform 1 0 38864 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2264_
timestamp 1698431365
transform 1 0 42448 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2265_
timestamp 1698431365
transform -1 0 42224 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2266_
timestamp 1698431365
transform -1 0 42448 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2267_
timestamp 1698431365
transform 1 0 29568 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2268_
timestamp 1698431365
transform 1 0 39088 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2269_
timestamp 1698431365
transform -1 0 40432 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2270_
timestamp 1698431365
transform -1 0 41664 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2271_
timestamp 1698431365
transform -1 0 38976 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2272_
timestamp 1698431365
transform 1 0 37856 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2273_
timestamp 1698431365
transform 1 0 37856 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _2274_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29904 0 -1 32928
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2275_
timestamp 1698431365
transform -1 0 39536 0 -1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2276_
timestamp 1698431365
transform 1 0 37184 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2277_
timestamp 1698431365
transform -1 0 36624 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2278_
timestamp 1698431365
transform 1 0 35616 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2279_
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2280_
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2281_
timestamp 1698431365
transform 1 0 35616 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2282_
timestamp 1698431365
transform -1 0 35616 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2283_
timestamp 1698431365
transform -1 0 37296 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2284_
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2285_
timestamp 1698431365
transform 1 0 36064 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2286_
timestamp 1698431365
transform -1 0 39872 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2287_
timestamp 1698431365
transform -1 0 36400 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2288_
timestamp 1698431365
transform 1 0 31584 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2289_
timestamp 1698431365
transform 1 0 34608 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2290_
timestamp 1698431365
transform 1 0 34160 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2291_
timestamp 1698431365
transform -1 0 41664 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2292_
timestamp 1698431365
transform -1 0 37968 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2293_
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2294_
timestamp 1698431365
transform 1 0 35616 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2295_
timestamp 1698431365
transform 1 0 36400 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2296_
timestamp 1698431365
transform 1 0 37072 0 -1 39200
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2297_
timestamp 1698431365
transform 1 0 39648 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2298_
timestamp 1698431365
transform 1 0 36624 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2299_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2300_
timestamp 1698431365
transform -1 0 40544 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2301_
timestamp 1698431365
transform -1 0 36624 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2302_
timestamp 1698431365
transform 1 0 34384 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2303_
timestamp 1698431365
transform 1 0 36624 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2304_
timestamp 1698431365
transform 1 0 35728 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2305_
timestamp 1698431365
transform -1 0 39648 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2306_
timestamp 1698431365
transform -1 0 38192 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2307_
timestamp 1698431365
transform 1 0 38192 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2308_
timestamp 1698431365
transform 1 0 34048 0 -1 42336
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2309_
timestamp 1698431365
transform 1 0 37408 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2310_
timestamp 1698431365
transform 1 0 38864 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2311_
timestamp 1698431365
transform -1 0 41104 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2312_
timestamp 1698431365
transform -1 0 35056 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2313_
timestamp 1698431365
transform 1 0 38192 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2314_
timestamp 1698431365
transform -1 0 37408 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2315_
timestamp 1698431365
transform 1 0 39536 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2316_
timestamp 1698431365
transform 1 0 37520 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2317_
timestamp 1698431365
transform -1 0 38976 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2318_
timestamp 1698431365
transform -1 0 39424 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2319_
timestamp 1698431365
transform -1 0 40096 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2320_
timestamp 1698431365
transform 1 0 41776 0 1 40768
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2321_
timestamp 1698431365
transform 1 0 46368 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _2322_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 43680 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2323_
timestamp 1698431365
transform 1 0 43568 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2324_
timestamp 1698431365
transform 1 0 46592 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2325_
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2326_
timestamp 1698431365
transform -1 0 43568 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2327_
timestamp 1698431365
transform -1 0 45136 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2328_
timestamp 1698431365
transform 1 0 42560 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2329_
timestamp 1698431365
transform -1 0 45136 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2330_
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2331_
timestamp 1698431365
transform -1 0 44464 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2332_
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2333_
timestamp 1698431365
transform 1 0 45472 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2334_
timestamp 1698431365
transform -1 0 45808 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2335_
timestamp 1698431365
transform 1 0 44576 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2336_
timestamp 1698431365
transform 1 0 46592 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2337_
timestamp 1698431365
transform 1 0 46704 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2338_
timestamp 1698431365
transform -1 0 46704 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2339_
timestamp 1698431365
transform -1 0 47600 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2340_
timestamp 1698431365
transform -1 0 46144 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2341_
timestamp 1698431365
transform 1 0 47264 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2342_
timestamp 1698431365
transform -1 0 46368 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2343_
timestamp 1698431365
transform -1 0 44128 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2344_
timestamp 1698431365
transform 1 0 43344 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2345_
timestamp 1698431365
transform -1 0 44128 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2346_
timestamp 1698431365
transform -1 0 47264 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2347_
timestamp 1698431365
transform -1 0 46368 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2348_
timestamp 1698431365
transform -1 0 44576 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2349_
timestamp 1698431365
transform -1 0 43456 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2350_
timestamp 1698431365
transform -1 0 42000 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2351_
timestamp 1698431365
transform -1 0 41216 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2352_
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2353_
timestamp 1698431365
transform -1 0 41888 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2354_
timestamp 1698431365
transform 1 0 38752 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2355_
timestamp 1698431365
transform 1 0 43792 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2356_
timestamp 1698431365
transform -1 0 44352 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2357_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41328 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2358_
timestamp 1698431365
transform 1 0 42336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2359_
timestamp 1698431365
transform -1 0 42896 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2360_
timestamp 1698431365
transform 1 0 38416 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2361_
timestamp 1698431365
transform -1 0 44688 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _2362_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40992 0 -1 37632
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2363_
timestamp 1698431365
transform 1 0 40544 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2364_
timestamp 1698431365
transform 1 0 42784 0 -1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2365_
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2366_
timestamp 1698431365
transform 1 0 47264 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2367_
timestamp 1698431365
transform -1 0 42224 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2368_
timestamp 1698431365
transform 1 0 41328 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2369_
timestamp 1698431365
transform 1 0 40096 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _2370_
timestamp 1698431365
transform -1 0 43680 0 -1 42336
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2371_
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _2372_
timestamp 1698431365
transform 1 0 38976 0 1 40768
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2373_
timestamp 1698431365
transform -1 0 42672 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _2374_
timestamp 1698431365
transform 1 0 44016 0 -1 40768
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2375_
timestamp 1698431365
transform -1 0 47264 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2376_
timestamp 1698431365
transform 1 0 42896 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2377_
timestamp 1698431365
transform 1 0 44576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2378_
timestamp 1698431365
transform -1 0 46368 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2379_
timestamp 1698431365
transform 1 0 47264 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2380_
timestamp 1698431365
transform -1 0 43008 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2381_
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2382_
timestamp 1698431365
transform 1 0 22848 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2383_
timestamp 1698431365
transform 1 0 16128 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2384_
timestamp 1698431365
transform -1 0 12208 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2385_
timestamp 1698431365
transform 1 0 20160 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2386_
timestamp 1698431365
transform 1 0 18816 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2387_
timestamp 1698431365
transform -1 0 20944 0 1 15680
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2388_
timestamp 1698431365
transform 1 0 25312 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2389_
timestamp 1698431365
transform 1 0 24752 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2390_
timestamp 1698431365
transform 1 0 30128 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2391_
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2392_
timestamp 1698431365
transform 1 0 16688 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2393_
timestamp 1698431365
transform 1 0 25536 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2394_
timestamp 1698431365
transform 1 0 26656 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2395_
timestamp 1698431365
transform 1 0 25984 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2396_
timestamp 1698431365
transform 1 0 24640 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2397_
timestamp 1698431365
transform 1 0 29232 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2398_
timestamp 1698431365
transform 1 0 27440 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2399_
timestamp 1698431365
transform 1 0 28336 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2400_
timestamp 1698431365
transform 1 0 27888 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2401_
timestamp 1698431365
transform -1 0 26768 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2402_
timestamp 1698431365
transform 1 0 26208 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2403_
timestamp 1698431365
transform 1 0 25424 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2404_
timestamp 1698431365
transform -1 0 26208 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2405_
timestamp 1698431365
transform -1 0 24864 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2406_
timestamp 1698431365
transform -1 0 25648 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2407_
timestamp 1698431365
transform -1 0 26880 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2408_
timestamp 1698431365
transform 1 0 25424 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2409_
timestamp 1698431365
transform 1 0 13104 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _2410_
timestamp 1698431365
transform 1 0 16800 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2411_
timestamp 1698431365
transform -1 0 19264 0 1 17248
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2412_
timestamp 1698431365
transform -1 0 15456 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2413_
timestamp 1698431365
transform 1 0 16800 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2414_
timestamp 1698431365
transform 1 0 16128 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2415_
timestamp 1698431365
transform 1 0 14784 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2416_
timestamp 1698431365
transform -1 0 25984 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2417_
timestamp 1698431365
transform 1 0 17584 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2418_
timestamp 1698431365
transform 1 0 18480 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2419_
timestamp 1698431365
transform 1 0 6608 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2420_
timestamp 1698431365
transform 1 0 15456 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2421_
timestamp 1698431365
transform 1 0 20160 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2422_
timestamp 1698431365
transform 1 0 17472 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2423_
timestamp 1698431365
transform 1 0 5712 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2424_
timestamp 1698431365
transform -1 0 10080 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2425_
timestamp 1698431365
transform 1 0 16128 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2426_
timestamp 1698431365
transform 1 0 14896 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2427_
timestamp 1698431365
transform 1 0 18368 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2428_
timestamp 1698431365
transform 1 0 16128 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2429_
timestamp 1698431365
transform -1 0 20160 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2430_
timestamp 1698431365
transform 1 0 17472 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2431_
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2432_
timestamp 1698431365
transform 1 0 3696 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2433_
timestamp 1698431365
transform 1 0 5040 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2434_
timestamp 1698431365
transform 1 0 6496 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2435_
timestamp 1698431365
transform 1 0 5600 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2436_
timestamp 1698431365
transform -1 0 9184 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2437_
timestamp 1698431365
transform 1 0 6608 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2438_
timestamp 1698431365
transform 1 0 6832 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2439_
timestamp 1698431365
transform 1 0 4368 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2440_
timestamp 1698431365
transform 1 0 6384 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2441_
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2442_
timestamp 1698431365
transform 1 0 6496 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2443_
timestamp 1698431365
transform 1 0 5936 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2444_
timestamp 1698431365
transform 1 0 8288 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2445_
timestamp 1698431365
transform 1 0 7392 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2446_
timestamp 1698431365
transform 1 0 29680 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2447_
timestamp 1698431365
transform -1 0 8176 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2448_
timestamp 1698431365
transform 1 0 8176 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2449_
timestamp 1698431365
transform 1 0 22848 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2450_
timestamp 1698431365
transform 1 0 23968 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2451_
timestamp 1698431365
transform -1 0 24416 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2452_
timestamp 1698431365
transform -1 0 24416 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2453_
timestamp 1698431365
transform 1 0 13776 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2454_
timestamp 1698431365
transform 1 0 19264 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2455_
timestamp 1698431365
transform 1 0 21056 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2456_
timestamp 1698431365
transform 1 0 21392 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2457_
timestamp 1698431365
transform 1 0 22288 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2458_
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2459_
timestamp 1698431365
transform 1 0 23744 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2460_
timestamp 1698431365
transform -1 0 25424 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2461_
timestamp 1698431365
transform -1 0 23632 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2462_
timestamp 1698431365
transform 1 0 23744 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2463_
timestamp 1698431365
transform 1 0 20384 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2464_
timestamp 1698431365
transform 1 0 21728 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2465_
timestamp 1698431365
transform -1 0 24080 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2466_
timestamp 1698431365
transform -1 0 22288 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2467_
timestamp 1698431365
transform -1 0 24752 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2468_
timestamp 1698431365
transform 1 0 13552 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2469_
timestamp 1698431365
transform 1 0 19040 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2470_
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2471_
timestamp 1698431365
transform -1 0 22736 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2472_
timestamp 1698431365
transform -1 0 19600 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2473_
timestamp 1698431365
transform 1 0 16240 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2474_
timestamp 1698431365
transform 1 0 19152 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2475_
timestamp 1698431365
transform 1 0 16912 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2476_
timestamp 1698431365
transform 1 0 23072 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2477_
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2478_
timestamp 1698431365
transform 1 0 15232 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2479_
timestamp 1698431365
transform 1 0 18928 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2480_
timestamp 1698431365
transform -1 0 18928 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2481_
timestamp 1698431365
transform -1 0 18368 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2482_
timestamp 1698431365
transform 1 0 16240 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2483_
timestamp 1698431365
transform -1 0 19040 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2484_
timestamp 1698431365
transform -1 0 28784 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2485_
timestamp 1698431365
transform -1 0 8848 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2486_
timestamp 1698431365
transform -1 0 8176 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2487_
timestamp 1698431365
transform -1 0 4368 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2488_
timestamp 1698431365
transform -1 0 6608 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2489_
timestamp 1698431365
transform 1 0 4704 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2490_
timestamp 1698431365
transform -1 0 8176 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2491_
timestamp 1698431365
transform 1 0 5824 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2492_
timestamp 1698431365
transform 1 0 4704 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2493_
timestamp 1698431365
transform 1 0 5824 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2494_
timestamp 1698431365
transform 1 0 4144 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2495_
timestamp 1698431365
transform 1 0 6944 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2496_
timestamp 1698431365
transform -1 0 19264 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2497_
timestamp 1698431365
transform -1 0 16800 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2498_
timestamp 1698431365
transform -1 0 12768 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2499_
timestamp 1698431365
transform -1 0 11312 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2500_
timestamp 1698431365
transform -1 0 10640 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2501_
timestamp 1698431365
transform -1 0 8064 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2502_
timestamp 1698431365
transform 1 0 10304 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2503_
timestamp 1698431365
transform 1 0 9744 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2504_
timestamp 1698431365
transform 1 0 11984 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2505_
timestamp 1698431365
transform 1 0 14336 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2506_
timestamp 1698431365
transform 1 0 11984 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2507_
timestamp 1698431365
transform -1 0 11200 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2508_
timestamp 1698431365
transform -1 0 8064 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2509_
timestamp 1698431365
transform 1 0 11312 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2510_
timestamp 1698431365
transform -1 0 13104 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2511_
timestamp 1698431365
transform -1 0 15008 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2512_
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2513_
timestamp 1698431365
transform 1 0 15008 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2514_
timestamp 1698431365
transform -1 0 15120 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2515_
timestamp 1698431365
transform 1 0 11536 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2516_
timestamp 1698431365
transform 1 0 35392 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2517_
timestamp 1698431365
transform -1 0 33600 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2518_
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2519_
timestamp 1698431365
transform -1 0 32368 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2520_
timestamp 1698431365
transform 1 0 30576 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2521_
timestamp 1698431365
transform -1 0 32256 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2522_
timestamp 1698431365
transform 1 0 31136 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2523_
timestamp 1698431365
transform -1 0 35168 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2524_
timestamp 1698431365
transform 1 0 33152 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2525_
timestamp 1698431365
transform 1 0 33712 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2526_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32032 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2527_
timestamp 1698431365
transform -1 0 16576 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2528_
timestamp 1698431365
transform 1 0 15232 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2529_
timestamp 1698431365
transform -1 0 17024 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2530_
timestamp 1698431365
transform -1 0 17248 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2531_
timestamp 1698431365
transform 1 0 27888 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2532_
timestamp 1698431365
transform 1 0 25536 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2533_
timestamp 1698431365
transform 1 0 27216 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2534_
timestamp 1698431365
transform 1 0 23968 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2535_
timestamp 1698431365
transform 1 0 30688 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2536_
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2537_
timestamp 1698431365
transform 1 0 32256 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2538_
timestamp 1698431365
transform 1 0 30576 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2539_
timestamp 1698431365
transform -1 0 35280 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2540_
timestamp 1698431365
transform -1 0 36176 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2541_
timestamp 1698431365
transform 1 0 23184 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2542_
timestamp 1698431365
transform 1 0 20048 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2543_
timestamp 1698431365
transform 1 0 17248 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2544_
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2545_
timestamp 1698431365
transform 1 0 17248 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2546_
timestamp 1698431365
transform 1 0 18144 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2547_
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2548_
timestamp 1698431365
transform 1 0 13888 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2549_
timestamp 1698431365
transform 1 0 16576 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2550_
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2551_
timestamp 1698431365
transform -1 0 11088 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2552_
timestamp 1698431365
transform -1 0 18592 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2553_
timestamp 1698431365
transform -1 0 18480 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2554_
timestamp 1698431365
transform 1 0 10864 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2555_
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2556_
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2557_
timestamp 1698431365
transform -1 0 4816 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2558_
timestamp 1698431365
transform 1 0 1680 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2559_
timestamp 1698431365
transform -1 0 17024 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2560_
timestamp 1698431365
transform 1 0 13776 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2561_
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2562_
timestamp 1698431365
transform -1 0 4816 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2563_
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2564_
timestamp 1698431365
transform -1 0 9184 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2565_
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2566_
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2567_
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2568_
timestamp 1698431365
transform 1 0 4816 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2569_
timestamp 1698431365
transform 1 0 4704 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2570_
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2571_
timestamp 1698431365
transform 1 0 12992 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2572_
timestamp 1698431365
transform 1 0 41664 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2573_
timestamp 1698431365
transform 1 0 41216 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2574_
timestamp 1698431365
transform 1 0 45136 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2575_
timestamp 1698431365
transform 1 0 45136 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2576_
timestamp 1698431365
transform 1 0 42112 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2577_
timestamp 1698431365
transform 1 0 43120 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2578_
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2579_
timestamp 1698431365
transform -1 0 43344 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2580_
timestamp 1698431365
transform -1 0 44464 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2581_
timestamp 1698431365
transform 1 0 41216 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2582_
timestamp 1698431365
transform 1 0 45136 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2583_
timestamp 1698431365
transform 1 0 45136 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2584_
timestamp 1698431365
transform 1 0 45136 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2585_
timestamp 1698431365
transform 1 0 45136 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2586_
timestamp 1698431365
transform 1 0 42224 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2587_
timestamp 1698431365
transform 1 0 45136 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2588_
timestamp 1698431365
transform 1 0 45136 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2589_
timestamp 1698431365
transform 1 0 45136 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2590_
timestamp 1698431365
transform 1 0 45136 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2591_
timestamp 1698431365
transform 1 0 45136 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2592_
timestamp 1698431365
transform 1 0 44016 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2593_
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2594_
timestamp 1698431365
transform -1 0 44128 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2595_
timestamp 1698431365
transform 1 0 37632 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2596_
timestamp 1698431365
transform 1 0 36288 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2597_
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2598_
timestamp 1698431365
transform 1 0 33936 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2599_
timestamp 1698431365
transform -1 0 40320 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2600_
timestamp 1698431365
transform -1 0 42336 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2601_
timestamp 1698431365
transform -1 0 38976 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2602_
timestamp 1698431365
transform 1 0 36960 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2603_
timestamp 1698431365
transform -1 0 37744 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2604_
timestamp 1698431365
transform -1 0 36624 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2605_
timestamp 1698431365
transform 1 0 31808 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2606_
timestamp 1698431365
transform 1 0 23408 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2607_
timestamp 1698431365
transform -1 0 30240 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2608_
timestamp 1698431365
transform -1 0 29792 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2609_
timestamp 1698431365
transform -1 0 30240 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2610_
timestamp 1698431365
transform 1 0 20944 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2611_
timestamp 1698431365
transform 1 0 17696 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2612_
timestamp 1698431365
transform -1 0 44800 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2613_
timestamp 1698431365
transform -1 0 44688 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2614_
timestamp 1698431365
transform 1 0 40880 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2615_
timestamp 1698431365
transform 1 0 39088 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2616_
timestamp 1698431365
transform -1 0 42896 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2617_
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2618_
timestamp 1698431365
transform -1 0 39424 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2619_
timestamp 1698431365
transform -1 0 39984 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2620_
timestamp 1698431365
transform 1 0 34720 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2621_
timestamp 1698431365
transform 1 0 33376 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2622_
timestamp 1698431365
transform -1 0 34832 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2623_
timestamp 1698431365
transform -1 0 36400 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2624_
timestamp 1698431365
transform -1 0 36176 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2625_
timestamp 1698431365
transform 1 0 30352 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2626_
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2627_
timestamp 1698431365
transform 1 0 20608 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2628_
timestamp 1698431365
transform 1 0 17360 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2629_
timestamp 1698431365
transform 1 0 18368 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2630_
timestamp 1698431365
transform -1 0 24752 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2631_
timestamp 1698431365
transform 1 0 21616 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2632_
timestamp 1698431365
transform -1 0 24752 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _2633_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2634_
timestamp 1698431365
transform -1 0 13888 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2635_
timestamp 1698431365
transform -1 0 13776 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2636_
timestamp 1698431365
transform 1 0 8624 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2637_
timestamp 1698431365
transform 1 0 5936 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2638_
timestamp 1698431365
transform 1 0 3696 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2639_
timestamp 1698431365
transform 1 0 3248 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2640_
timestamp 1698431365
transform 1 0 3472 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2641_
timestamp 1698431365
transform -1 0 12880 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2642_
timestamp 1698431365
transform 1 0 10416 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2643_
timestamp 1698431365
transform -1 0 11424 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _2644_
timestamp 1698431365
transform -1 0 10976 0 1 21952
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2645_
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2646_
timestamp 1698431365
transform 1 0 38304 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2647_
timestamp 1698431365
transform -1 0 42448 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2648_
timestamp 1698431365
transform -1 0 38192 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2649_
timestamp 1698431365
transform -1 0 38752 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2650_
timestamp 1698431365
transform 1 0 31808 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2651_
timestamp 1698431365
transform -1 0 41328 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2652_
timestamp 1698431365
transform 1 0 33376 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2653_
timestamp 1698431365
transform 1 0 33040 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2654_
timestamp 1698431365
transform 1 0 36288 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2655_
timestamp 1698431365
transform -1 0 48384 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2656_
timestamp 1698431365
transform -1 0 48384 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2657_
timestamp 1698431365
transform -1 0 48384 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2658_
timestamp 1698431365
transform 1 0 45136 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2659_
timestamp 1698431365
transform 1 0 43232 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2660_
timestamp 1698431365
transform 1 0 45136 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2661_
timestamp 1698431365
transform 1 0 45136 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2662_
timestamp 1698431365
transform 1 0 45136 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2663_
timestamp 1698431365
transform 1 0 29344 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2664_
timestamp 1698431365
transform -1 0 45024 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2665_
timestamp 1698431365
transform 1 0 39200 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2666_
timestamp 1698431365
transform 1 0 37744 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2667_
timestamp 1698431365
transform -1 0 45360 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2668_
timestamp 1698431365
transform 1 0 37296 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2669_
timestamp 1698431365
transform 1 0 40992 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2670_
timestamp 1698431365
transform -1 0 48384 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2671_
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2672_
timestamp 1698431365
transform -1 0 42784 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2673_
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2674_
timestamp 1698431365
transform 1 0 41216 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2675_
timestamp 1698431365
transform -1 0 48384 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2676_
timestamp 1698431365
transform -1 0 48048 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2677_
timestamp 1698431365
transform 1 0 41552 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2678_
timestamp 1698431365
transform 1 0 28336 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2679_
timestamp 1698431365
transform 1 0 24752 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2680_
timestamp 1698431365
transform 1 0 27104 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2681_
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2682_
timestamp 1698431365
transform 1 0 24304 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2683_
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2684_
timestamp 1698431365
transform 1 0 13440 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2685_
timestamp 1698431365
transform 1 0 15456 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2686_
timestamp 1698431365
transform 1 0 17472 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2687_
timestamp 1698431365
transform 1 0 13664 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2688_
timestamp 1698431365
transform 1 0 17696 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2689_
timestamp 1698431365
transform 1 0 17696 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2690_
timestamp 1698431365
transform 1 0 3584 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2691_
timestamp 1698431365
transform 1 0 2016 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2692_
timestamp 1698431365
transform 1 0 3248 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2693_
timestamp 1698431365
transform 1 0 2912 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2694_
timestamp 1698431365
transform 1 0 6832 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2695_
timestamp 1698431365
transform 1 0 5712 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2696_
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2697_
timestamp 1698431365
transform 1 0 23632 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2698_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21392 0 1 21952
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2699_
timestamp 1698431365
transform 1 0 20496 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2700_
timestamp 1698431365
transform 1 0 15680 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2701_
timestamp 1698431365
transform 1 0 15792 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2702_
timestamp 1698431365
transform 1 0 18592 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2703_
timestamp 1698431365
transform -1 0 18816 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2704_
timestamp 1698431365
transform -1 0 5040 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2705_
timestamp 1698431365
transform 1 0 1792 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _2706_
timestamp 1698431365
transform 1 0 2240 0 -1 18816
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2707_
timestamp 1698431365
transform -1 0 4816 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2708_
timestamp 1698431365
transform 1 0 8176 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _2709_
timestamp 1698431365
transform 1 0 12096 0 -1 20384
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2710_
timestamp 1698431365
transform 1 0 11872 0 -1 21952
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2711_
timestamp 1698431365
transform 1 0 8064 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2712_
timestamp 1698431365
transform -1 0 14112 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2713_
timestamp 1698431365
transform -1 0 16128 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2714_
timestamp 1698431365
transform 1 0 13664 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2715_
timestamp 1698431365
transform 1 0 38304 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2716_
timestamp 1698431365
transform 1 0 29904 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2717_
timestamp 1698431365
transform -1 0 34048 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2718_
timestamp 1698431365
transform 1 0 33600 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1260__A2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13552 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1268__I
timestamp 1698431365
transform -1 0 3808 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1270__A2
timestamp 1698431365
transform 1 0 16800 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1271__A1
timestamp 1698431365
transform 1 0 23184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1271__A2
timestamp 1698431365
transform 1 0 25312 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1272__I
timestamp 1698431365
transform 1 0 19040 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1277__A1
timestamp 1698431365
transform -1 0 15456 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1286__A3
timestamp 1698431365
transform -1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1292__A1
timestamp 1698431365
transform 1 0 35392 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1296__A3
timestamp 1698431365
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1297__A1
timestamp 1698431365
transform 1 0 36512 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1311__A2
timestamp 1698431365
transform -1 0 2240 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1315__A3
timestamp 1698431365
transform -1 0 3360 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1316__A1
timestamp 1698431365
transform 1 0 3584 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1317__B
timestamp 1698431365
transform -1 0 3360 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1330__B
timestamp 1698431365
transform 1 0 7616 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1338__A2
timestamp 1698431365
transform 1 0 27776 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1343__B
timestamp 1698431365
transform 1 0 19824 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1344__A1
timestamp 1698431365
transform -1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1345__B2
timestamp 1698431365
transform 1 0 25312 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1356__A1
timestamp 1698431365
transform -1 0 5936 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1356__A2
timestamp 1698431365
transform 1 0 14896 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1356__B
timestamp 1698431365
transform -1 0 5936 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1360__I
timestamp 1698431365
transform 1 0 18704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1370__A1
timestamp 1698431365
transform -1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1371__A1
timestamp 1698431365
transform 1 0 32256 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1375__A2
timestamp 1698431365
transform -1 0 29568 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1377__A2
timestamp 1698431365
transform -1 0 2800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1378__A3
timestamp 1698431365
transform 1 0 18368 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1379__B
timestamp 1698431365
transform 1 0 11536 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1391__A2
timestamp 1698431365
transform 1 0 10752 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1394__A2
timestamp 1698431365
transform -1 0 11760 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1394__A3
timestamp 1698431365
transform -1 0 2800 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1397__A2
timestamp 1698431365
transform -1 0 7504 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1398__B1
timestamp 1698431365
transform 1 0 11312 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1404__A3
timestamp 1698431365
transform -1 0 31472 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1409__A1
timestamp 1698431365
transform -1 0 15344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1431__A1
timestamp 1698431365
transform 1 0 25760 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1435__A1
timestamp 1698431365
transform -1 0 2352 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1437__A2
timestamp 1698431365
transform 1 0 12320 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1438__A1
timestamp 1698431365
transform -1 0 10976 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1438__B
timestamp 1698431365
transform -1 0 12656 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1439__A1
timestamp 1698431365
transform 1 0 27552 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1439__A3
timestamp 1698431365
transform 1 0 5040 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1440__A1
timestamp 1698431365
transform -1 0 13776 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1461__A1
timestamp 1698431365
transform 1 0 5712 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1512__A3
timestamp 1698431365
transform -1 0 16128 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1513__A2
timestamp 1698431365
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1520__A1
timestamp 1698431365
transform -1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1544__A1
timestamp 1698431365
transform -1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1551__I
timestamp 1698431365
transform -1 0 8736 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1557__A1
timestamp 1698431365
transform 1 0 24416 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1559__A1
timestamp 1698431365
transform -1 0 31920 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1574__I
timestamp 1698431365
transform 1 0 25760 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1580__A1
timestamp 1698431365
transform -1 0 8960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1606__A1
timestamp 1698431365
transform -1 0 11424 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1607__I
timestamp 1698431365
transform -1 0 12320 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1627__A2
timestamp 1698431365
transform 1 0 32480 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1633__A2
timestamp 1698431365
transform 1 0 29568 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1637__A1
timestamp 1698431365
transform 1 0 47376 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1641__I
timestamp 1698431365
transform -1 0 29456 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1642__I
timestamp 1698431365
transform 1 0 27552 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1643__I
timestamp 1698431365
transform 1 0 27440 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1644__I
timestamp 1698431365
transform -1 0 3136 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1645__A1
timestamp 1698431365
transform -1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1650__A1
timestamp 1698431365
transform -1 0 10304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1651__I
timestamp 1698431365
transform 1 0 28784 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1654__C
timestamp 1698431365
transform -1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__I
timestamp 1698431365
transform -1 0 21056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1657__I
timestamp 1698431365
transform 1 0 20048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__I
timestamp 1698431365
transform -1 0 10192 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1659__I
timestamp 1698431365
transform 1 0 4592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1660__I
timestamp 1698431365
transform -1 0 22848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__A1
timestamp 1698431365
transform -1 0 10528 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1663__I
timestamp 1698431365
transform 1 0 35840 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__I
timestamp 1698431365
transform 1 0 30464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A1
timestamp 1698431365
transform -1 0 14672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__I
timestamp 1698431365
transform 1 0 26992 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1670__A1
timestamp 1698431365
transform -1 0 14224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1672__I
timestamp 1698431365
transform -1 0 28560 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1677__A1
timestamp 1698431365
transform 1 0 28560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__C
timestamp 1698431365
transform 1 0 31248 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1680__A1
timestamp 1698431365
transform 1 0 26768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__I
timestamp 1698431365
transform 1 0 28112 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1683__A1
timestamp 1698431365
transform 1 0 29456 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1685__A1
timestamp 1698431365
transform 1 0 28336 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1687__A1
timestamp 1698431365
transform -1 0 25536 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__A1
timestamp 1698431365
transform 1 0 32480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1692__C
timestamp 1698431365
transform 1 0 30464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1694__A1
timestamp 1698431365
transform 1 0 29120 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1696__A1
timestamp 1698431365
transform 1 0 30800 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1697__I
timestamp 1698431365
transform -1 0 22512 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1698__I
timestamp 1698431365
transform -1 0 19488 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1699__B
timestamp 1698431365
transform 1 0 35952 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__A1
timestamp 1698431365
transform 1 0 36400 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1701__B
timestamp 1698431365
transform 1 0 34048 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1703__I
timestamp 1698431365
transform 1 0 44912 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1708__A1
timestamp 1698431365
transform 1 0 36624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1713__B
timestamp 1698431365
transform 1 0 26768 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1717__I
timestamp 1698431365
transform 1 0 24640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1728__B
timestamp 1698431365
transform -1 0 18480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1734__I
timestamp 1698431365
transform 1 0 23072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1735__B
timestamp 1698431365
transform 1 0 19936 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1752__I
timestamp 1698431365
transform -1 0 13216 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1760__B
timestamp 1698431365
transform -1 0 18368 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1763__B
timestamp 1698431365
transform 1 0 12544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1785__B
timestamp 1698431365
transform -1 0 12320 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__I
timestamp 1698431365
transform 1 0 5712 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1801__I
timestamp 1698431365
transform -1 0 14560 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1806__A1
timestamp 1698431365
transform -1 0 5936 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1818__A1
timestamp 1698431365
transform -1 0 15568 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1821__I
timestamp 1698431365
transform 1 0 35840 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1822__B
timestamp 1698431365
transform 1 0 16912 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1828__A2
timestamp 1698431365
transform 1 0 3696 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1829__A1
timestamp 1698431365
transform -1 0 2464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1830__A2
timestamp 1698431365
transform 1 0 2240 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1831__A2
timestamp 1698431365
transform 1 0 2688 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1834__I
timestamp 1698431365
transform 1 0 5264 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1841__A1
timestamp 1698431365
transform 1 0 7616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1861__I
timestamp 1698431365
transform 1 0 39984 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1866__A1
timestamp 1698431365
transform 1 0 9632 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1871__A1
timestamp 1698431365
transform 1 0 8960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1877__A1
timestamp 1698431365
transform 1 0 10752 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1879__I
timestamp 1698431365
transform -1 0 4144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1880__I
timestamp 1698431365
transform -1 0 35392 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1881__B
timestamp 1698431365
transform -1 0 11872 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1885__A2
timestamp 1698431365
transform -1 0 42000 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1887__A1
timestamp 1698431365
transform 1 0 41440 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1891__A1
timestamp 1698431365
transform 1 0 47488 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1894__A1
timestamp 1698431365
transform 1 0 48160 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1895__I
timestamp 1698431365
transform 1 0 41104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__I
timestamp 1698431365
transform 1 0 44912 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1902__A1
timestamp 1698431365
transform 1 0 42224 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1914__A1
timestamp 1698431365
transform 1 0 44016 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1968__I
timestamp 1698431365
transform -1 0 45136 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1970__A2
timestamp 1698431365
transform -1 0 46480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1973__A2
timestamp 1698431365
transform 1 0 46592 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__I
timestamp 1698431365
transform 1 0 40208 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1975__A2
timestamp 1698431365
transform 1 0 42336 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1978__A2
timestamp 1698431365
transform -1 0 45136 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1981__I
timestamp 1698431365
transform -1 0 15120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1982__I
timestamp 1698431365
transform 1 0 25760 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1984__A2
timestamp 1698431365
transform 1 0 40208 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1987__A1
timestamp 1698431365
transform 1 0 40992 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1989__B
timestamp 1698431365
transform 1 0 38640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1993__I
timestamp 1698431365
transform 1 0 37968 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__B
timestamp 1698431365
transform 1 0 39536 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1997__B
timestamp 1698431365
transform 1 0 37072 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2001__A1
timestamp 1698431365
transform 1 0 41104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2006__B
timestamp 1698431365
transform -1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2012__A1
timestamp 1698431365
transform 1 0 38528 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2016__B
timestamp 1698431365
transform 1 0 36400 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2018__I
timestamp 1698431365
transform 1 0 35952 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2023__A1
timestamp 1698431365
transform 1 0 35728 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2029__B
timestamp 1698431365
transform 1 0 33376 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2035__I
timestamp 1698431365
transform 1 0 36064 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2036__B
timestamp 1698431365
transform 1 0 29680 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2042__A1
timestamp 1698431365
transform 1 0 28560 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2047__B
timestamp 1698431365
transform 1 0 27776 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2052__A2
timestamp 1698431365
transform 1 0 26432 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2053__B
timestamp 1698431365
transform 1 0 28560 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2055__A2
timestamp 1698431365
transform 1 0 30464 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2056__A2
timestamp 1698431365
transform 1 0 26096 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2059__A1
timestamp 1698431365
transform 1 0 27440 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2062__C
timestamp 1698431365
transform 1 0 23408 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2064__I
timestamp 1698431365
transform 1 0 43456 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2065__A2
timestamp 1698431365
transform 1 0 43008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2071__A1
timestamp 1698431365
transform 1 0 40880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2072__B
timestamp 1698431365
transform 1 0 44128 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2073__I
timestamp 1698431365
transform -1 0 10080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2074__I
timestamp 1698431365
transform 1 0 37632 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2077__I
timestamp 1698431365
transform 1 0 32368 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2078__I
timestamp 1698431365
transform 1 0 34720 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2079__B
timestamp 1698431365
transform -1 0 40320 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2080__C
timestamp 1698431365
transform 1 0 43232 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2084__B
timestamp 1698431365
transform 1 0 44912 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2085__C
timestamp 1698431365
transform -1 0 39424 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2090__B
timestamp 1698431365
transform 1 0 40208 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2091__I
timestamp 1698431365
transform 1 0 32480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2100__I
timestamp 1698431365
transform 1 0 35168 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2110__A1
timestamp 1698431365
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2114__I
timestamp 1698431365
transform 1 0 37968 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2117__A1
timestamp 1698431365
transform 1 0 38416 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2119__A2
timestamp 1698431365
transform -1 0 40432 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2119__C
timestamp 1698431365
transform -1 0 39088 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2121__A1
timestamp 1698431365
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2122__I
timestamp 1698431365
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2123__A1
timestamp 1698431365
transform 1 0 34832 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2124__A2
timestamp 1698431365
transform 1 0 37744 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2125__B
timestamp 1698431365
transform 1 0 36960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2126__A1
timestamp 1698431365
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2129__A1
timestamp 1698431365
transform 1 0 38192 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2130__B
timestamp 1698431365
transform 1 0 36176 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2132__A2
timestamp 1698431365
transform 1 0 36624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2137__A1
timestamp 1698431365
transform 1 0 34832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2138__B
timestamp 1698431365
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2142__I
timestamp 1698431365
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2150__I
timestamp 1698431365
transform -1 0 23744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2166__I
timestamp 1698431365
transform -1 0 18480 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2173__A1
timestamp 1698431365
transform -1 0 23296 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2179__A1
timestamp 1698431365
transform 1 0 29680 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2181__A2
timestamp 1698431365
transform -1 0 26432 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2181__C
timestamp 1698431365
transform -1 0 27888 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2183__A1
timestamp 1698431365
transform 1 0 23856 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2184__A1
timestamp 1698431365
transform -1 0 23968 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2185__A2
timestamp 1698431365
transform -1 0 23072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2186__B
timestamp 1698431365
transform 1 0 23408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2188__A1
timestamp 1698431365
transform 1 0 22624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2189__A2
timestamp 1698431365
transform 1 0 24416 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2191__A1
timestamp 1698431365
transform 1 0 25872 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2192__I
timestamp 1698431365
transform 1 0 32704 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2193__A2
timestamp 1698431365
transform -1 0 3360 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2193__B
timestamp 1698431365
transform -1 0 3808 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2194__A2
timestamp 1698431365
transform -1 0 2464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2195__A2
timestamp 1698431365
transform -1 0 8176 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2200__A1
timestamp 1698431365
transform -1 0 12320 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2201__B
timestamp 1698431365
transform -1 0 11424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2202__I
timestamp 1698431365
transform -1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2210__I
timestamp 1698431365
transform -1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2218__I
timestamp 1698431365
transform -1 0 8512 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2229__A2
timestamp 1698431365
transform -1 0 5936 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2235__A1
timestamp 1698431365
transform -1 0 3248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2236__A2
timestamp 1698431365
transform -1 0 2800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2241__A1
timestamp 1698431365
transform -1 0 2240 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2243__A2
timestamp 1698431365
transform -1 0 3584 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2243__C
timestamp 1698431365
transform -1 0 4368 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2245__A1
timestamp 1698431365
transform -1 0 2912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2246__A1
timestamp 1698431365
transform -1 0 12432 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2247__A2
timestamp 1698431365
transform -1 0 6272 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2248__B
timestamp 1698431365
transform -1 0 9856 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2249__A1
timestamp 1698431365
transform -1 0 3920 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2252__A1
timestamp 1698431365
transform -1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2253__A1
timestamp 1698431365
transform 1 0 3472 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2253__B
timestamp 1698431365
transform 1 0 10416 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2254__A1
timestamp 1698431365
transform 1 0 3472 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2256__B
timestamp 1698431365
transform 1 0 38976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2260__A2
timestamp 1698431365
transform -1 0 29456 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2261__A2
timestamp 1698431365
transform 1 0 28560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2263__A1
timestamp 1698431365
transform 1 0 40320 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2269__B
timestamp 1698431365
transform 1 0 41440 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2276__A1
timestamp 1698431365
transform -1 0 40320 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2283__A1
timestamp 1698431365
transform -1 0 38864 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2288__I
timestamp 1698431365
transform 1 0 31360 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2289__B
timestamp 1698431365
transform 1 0 34384 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2297__A1
timestamp 1698431365
transform 1 0 40320 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2303__B
timestamp 1698431365
transform 1 0 35504 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2310__A1
timestamp 1698431365
transform 1 0 25760 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2315__B
timestamp 1698431365
transform -1 0 22512 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2321__A1
timestamp 1698431365
transform 1 0 32480 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2326__A1
timestamp 1698431365
transform -1 0 23968 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2329__C
timestamp 1698431365
transform -1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2334__C
timestamp 1698431365
transform 1 0 48048 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2345__B
timestamp 1698431365
transform 1 0 43008 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2348__A1
timestamp 1698431365
transform 1 0 46928 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2350__A2
timestamp 1698431365
transform -1 0 42112 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2353__A2
timestamp 1698431365
transform 1 0 43120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2354__A2
timestamp 1698431365
transform 1 0 39872 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2359__A2
timestamp 1698431365
transform 1 0 43120 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2360__A2
timestamp 1698431365
transform 1 0 40096 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2379__A2
timestamp 1698431365
transform -1 0 43568 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2380__A1
timestamp 1698431365
transform 1 0 42224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2381__I
timestamp 1698431365
transform 1 0 22736 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2385__I
timestamp 1698431365
transform 1 0 21952 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2390__B
timestamp 1698431365
transform -1 0 32704 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2391__A1
timestamp 1698431365
transform 1 0 30800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2392__I
timestamp 1698431365
transform -1 0 12656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2395__A1
timestamp 1698431365
transform 1 0 26432 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2398__A1
timestamp 1698431365
transform 1 0 29232 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2400__A1
timestamp 1698431365
transform 1 0 27776 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2403__A1
timestamp 1698431365
transform 1 0 27888 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2404__I
timestamp 1698431365
transform 1 0 27104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2408__A1
timestamp 1698431365
transform 1 0 25312 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2410__A2
timestamp 1698431365
transform -1 0 16128 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2415__A1
timestamp 1698431365
transform -1 0 15904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2416__I
timestamp 1698431365
transform 1 0 25984 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2418__A1
timestamp 1698431365
transform -1 0 19376 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2419__I
timestamp 1698431365
transform -1 0 3472 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2422__A1
timestamp 1698431365
transform -1 0 17472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2423__I
timestamp 1698431365
transform -1 0 2576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2426__A1
timestamp 1698431365
transform 1 0 6944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2428__A1
timestamp 1698431365
transform -1 0 19376 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2430__A1
timestamp 1698431365
transform -1 0 18928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2435__A1
timestamp 1698431365
transform -1 0 3472 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2438__A1
timestamp 1698431365
transform -1 0 3920 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2441__A1
timestamp 1698431365
transform -1 0 2128 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2443__A1
timestamp 1698431365
transform -1 0 4368 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2445__A1
timestamp 1698431365
transform -1 0 2128 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2447__B
timestamp 1698431365
transform -1 0 3024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2448__A1
timestamp 1698431365
transform -1 0 2016 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2452__A1
timestamp 1698431365
transform -1 0 24640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2452__A2
timestamp 1698431365
transform 1 0 26320 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2455__A1
timestamp 1698431365
transform -1 0 21056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2459__A1
timestamp 1698431365
transform 1 0 23856 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2459__C
timestamp 1698431365
transform 1 0 26544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2462__A1
timestamp 1698431365
transform 1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2464__A1
timestamp 1698431365
transform 1 0 24080 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2465__A1
timestamp 1698431365
transform -1 0 24528 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2466__A1
timestamp 1698431365
transform 1 0 20720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2470__A1
timestamp 1698431365
transform 1 0 23856 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2474__A1
timestamp 1698431365
transform -1 0 20496 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2475__A1
timestamp 1698431365
transform -1 0 8736 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2477__A1
timestamp 1698431365
transform 1 0 19376 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2477__C
timestamp 1698431365
transform -1 0 18368 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2479__A1
timestamp 1698431365
transform 1 0 2128 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2479__C
timestamp 1698431365
transform 1 0 35616 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2480__A1
timestamp 1698431365
transform -1 0 16576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2481__A1
timestamp 1698431365
transform 1 0 14784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2481__C
timestamp 1698431365
transform -1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2482__A2
timestamp 1698431365
transform 1 0 11984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2484__A1
timestamp 1698431365
transform 1 0 28000 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2485__I
timestamp 1698431365
transform -1 0 4704 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2486__I
timestamp 1698431365
transform -1 0 2912 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2488__A1
timestamp 1698431365
transform 1 0 2352 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2488__C
timestamp 1698431365
transform -1 0 2352 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2490__I
timestamp 1698431365
transform -1 0 3472 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2491__A1
timestamp 1698431365
transform 1 0 5040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2493__A1
timestamp 1698431365
transform -1 0 4256 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2495__A1
timestamp 1698431365
transform 1 0 3248 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2497__A1
timestamp 1698431365
transform -1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2501__A1
timestamp 1698431365
transform -1 0 2464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2502__A1
timestamp 1698431365
transform -1 0 2912 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2503__I
timestamp 1698431365
transform -1 0 8736 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2504__A1
timestamp 1698431365
transform -1 0 4704 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2504__C
timestamp 1698431365
transform -1 0 3248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2505__A1
timestamp 1698431365
transform -1 0 15120 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2506__A1
timestamp 1698431365
transform 1 0 5712 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2506__C
timestamp 1698431365
transform 1 0 5040 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2507__A1
timestamp 1698431365
transform -1 0 3024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2508__A1
timestamp 1698431365
transform 1 0 2800 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2508__C
timestamp 1698431365
transform -1 0 6720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2510__B
timestamp 1698431365
transform 1 0 4144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2511__A1
timestamp 1698431365
transform 1 0 6384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2512__B
timestamp 1698431365
transform -1 0 18592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2513__A1
timestamp 1698431365
transform 1 0 10416 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2514__C
timestamp 1698431365
transform -1 0 3248 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2516__A1
timestamp 1698431365
transform 1 0 37296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2519__B
timestamp 1698431365
transform 1 0 31248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2520__A1
timestamp 1698431365
transform 1 0 30352 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2522__A1
timestamp 1698431365
transform 1 0 35056 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2524__A1
timestamp 1698431365
transform 1 0 37072 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2525__C
timestamp 1698431365
transform 1 0 36288 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2526__CLK
timestamp 1698431365
transform 1 0 33488 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2526__D
timestamp 1698431365
transform 1 0 33936 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2527__CLK
timestamp 1698431365
transform -1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2528__CLK
timestamp 1698431365
transform -1 0 10976 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2529__CLK
timestamp 1698431365
transform -1 0 9632 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2530__CLK
timestamp 1698431365
transform -1 0 11872 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2531__CLK
timestamp 1698431365
transform 1 0 29904 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2532__CLK
timestamp 1698431365
transform 1 0 30128 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2533__CLK
timestamp 1698431365
transform 1 0 30688 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2534__CLK
timestamp 1698431365
transform 1 0 24080 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2535__CLK
timestamp 1698431365
transform 1 0 35728 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2536__CLK
timestamp 1698431365
transform 1 0 32032 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2537__CLK
timestamp 1698431365
transform 1 0 37072 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2538__CLK
timestamp 1698431365
transform 1 0 36288 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2541__CLK
timestamp 1698431365
transform 1 0 21392 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2542__CLK
timestamp 1698431365
transform 1 0 22288 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2543__CLK
timestamp 1698431365
transform 1 0 27776 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2544__CLK
timestamp 1698431365
transform -1 0 19936 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2545__CLK
timestamp 1698431365
transform 1 0 20496 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2546__CLK
timestamp 1698431365
transform 1 0 22288 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2547__CLK
timestamp 1698431365
transform 1 0 20496 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2548__CLK
timestamp 1698431365
transform 1 0 9632 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2549__CLK
timestamp 1698431365
transform 1 0 22288 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2550__CLK
timestamp 1698431365
transform 1 0 11984 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2551__CLK
timestamp 1698431365
transform 1 0 4592 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2552__CLK
timestamp 1698431365
transform -1 0 19040 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2553__CLK
timestamp 1698431365
transform 1 0 25088 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2554__CLK
timestamp 1698431365
transform 1 0 14560 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2555__CLK
timestamp 1698431365
transform 1 0 3136 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2556__CLK
timestamp 1698431365
transform 1 0 5040 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2557__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2558__CLK
timestamp 1698431365
transform 1 0 4480 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2559__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2560__CLK
timestamp 1698431365
transform 1 0 11312 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2561__CLK
timestamp 1698431365
transform 1 0 1792 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2562__CLK
timestamp 1698431365
transform 1 0 4144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2563__CLK
timestamp 1698431365
transform 1 0 3136 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2564__CLK
timestamp 1698431365
transform 1 0 8288 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2565__CLK
timestamp 1698431365
transform 1 0 5040 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2566__CLK
timestamp 1698431365
transform 1 0 1792 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2567__CLK
timestamp 1698431365
transform 1 0 9296 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2568__CLK
timestamp 1698431365
transform 1 0 8288 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2569__CLK
timestamp 1698431365
transform 1 0 7952 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2570__CLK
timestamp 1698431365
transform 1 0 10864 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2571__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2581__CLK
timestamp 1698431365
transform 1 0 44912 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2582__CLK
timestamp 1698431365
transform -1 0 45136 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2583__CLK
timestamp 1698431365
transform 1 0 45360 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2584__CLK
timestamp 1698431365
transform 1 0 45584 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2585__CLK
timestamp 1698431365
transform 1 0 44912 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2586__CLK
timestamp 1698431365
transform 1 0 42784 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2587__CLK
timestamp 1698431365
transform 1 0 44912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2588__CLK
timestamp 1698431365
transform 1 0 44912 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2594__CLK
timestamp 1698431365
transform 1 0 44128 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2595__CLK
timestamp 1698431365
transform 1 0 40880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2605__CLK
timestamp 1698431365
transform -1 0 35504 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2606__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2607__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2608__CLK
timestamp 1698431365
transform 1 0 30016 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2609__CLK
timestamp 1698431365
transform 1 0 31360 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2610__CLK
timestamp 1698431365
transform 1 0 20048 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2611__CLK
timestamp 1698431365
transform 1 0 21840 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2612__CLK
timestamp 1698431365
transform 1 0 45696 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2613__CLK
timestamp 1698431365
transform 1 0 44912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2614__CLK
timestamp 1698431365
transform 1 0 44128 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2615__CLK
timestamp 1698431365
transform 1 0 43008 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2616__CLK
timestamp 1698431365
transform -1 0 43904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2617__CLK
timestamp 1698431365
transform 1 0 38864 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2618__CLK
timestamp 1698431365
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2620__CLK
timestamp 1698431365
transform 1 0 38192 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2623__CLK
timestamp 1698431365
transform 1 0 37184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2624__CLK
timestamp 1698431365
transform -1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2625__CLK
timestamp 1698431365
transform 1 0 35616 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2626__CLK
timestamp 1698431365
transform -1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2627__CLK
timestamp 1698431365
transform -1 0 28672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2628__CLK
timestamp 1698431365
transform 1 0 26208 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2629__CLK
timestamp 1698431365
transform -1 0 21952 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2630__CLK
timestamp 1698431365
transform -1 0 21504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2633__CLK
timestamp 1698431365
transform 1 0 2128 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2634__CLK
timestamp 1698431365
transform 1 0 9856 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2635__CLK
timestamp 1698431365
transform -1 0 7392 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2636__CLK
timestamp 1698431365
transform -1 0 6944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2637__CLK
timestamp 1698431365
transform -1 0 6496 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2638__CLK
timestamp 1698431365
transform 1 0 5264 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2639__CLK
timestamp 1698431365
transform 1 0 3472 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2640__CLK
timestamp 1698431365
transform 1 0 2800 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2641__CLK
timestamp 1698431365
transform 1 0 2464 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2642__CLK
timestamp 1698431365
transform 1 0 3696 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2643__CLK
timestamp 1698431365
transform 1 0 3024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2644__CLK
timestamp 1698431365
transform 1 0 10976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2650__CLK
timestamp 1698431365
transform 1 0 35056 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2651__CLK
timestamp 1698431365
transform 1 0 39872 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2652__CLK
timestamp 1698431365
transform 1 0 35952 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2653__CLK
timestamp 1698431365
transform 1 0 27328 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2654__CLK
timestamp 1698431365
transform 1 0 39088 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2655__CLK
timestamp 1698431365
transform 1 0 22848 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2656__CLK
timestamp 1698431365
transform -1 0 22064 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2657__CLK
timestamp 1698431365
transform 1 0 25200 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2658__CLK
timestamp 1698431365
transform 1 0 40320 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2661__CLK
timestamp 1698431365
transform 1 0 47824 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2662__CLK
timestamp 1698431365
transform 1 0 45360 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2663__CLK
timestamp 1698431365
transform 1 0 32032 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2663__D
timestamp 1698431365
transform 1 0 32480 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2667__CLK
timestamp 1698431365
transform 1 0 44912 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2668__CLK
timestamp 1698431365
transform 1 0 38192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2669__CLK
timestamp 1698431365
transform -1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2670__CLK
timestamp 1698431365
transform 1 0 28560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2671__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2672__CLK
timestamp 1698431365
transform 1 0 23296 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2673__CLK
timestamp 1698431365
transform 1 0 26320 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2674__CLK
timestamp 1698431365
transform 1 0 26768 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2675__CLK
timestamp 1698431365
transform 1 0 40992 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2676__CLK
timestamp 1698431365
transform 1 0 48160 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2678__CLK
timestamp 1698431365
transform 1 0 36848 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2679__CLK
timestamp 1698431365
transform 1 0 28560 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2680__CLK
timestamp 1698431365
transform 1 0 33600 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2681__CLK
timestamp 1698431365
transform 1 0 31920 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2682__CLK
timestamp 1698431365
transform 1 0 28224 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2684__CLK
timestamp 1698431365
transform 1 0 17696 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2685__CLK
timestamp 1698431365
transform -1 0 18928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2686__CLK
timestamp 1698431365
transform 1 0 21392 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2687__CLK
timestamp 1698431365
transform 1 0 8064 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2690__CLK
timestamp 1698431365
transform 1 0 5040 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2691__CLK
timestamp 1698431365
transform 1 0 4592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2692__CLK
timestamp 1698431365
transform 1 0 4592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2693__CLK
timestamp 1698431365
transform -1 0 2016 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2694__CLK
timestamp 1698431365
transform 1 0 2352 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2695__CLK
timestamp 1698431365
transform -1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2700__CLK
timestamp 1698431365
transform -1 0 19152 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2701__CLK
timestamp 1698431365
transform -1 0 6272 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2702__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2704__CLK
timestamp 1698431365
transform 1 0 1792 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2705__CLK
timestamp 1698431365
transform 1 0 1904 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2706__CLK
timestamp 1698431365
transform 1 0 2240 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2707__CLK
timestamp 1698431365
transform 1 0 1792 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2708__CLK
timestamp 1698431365
transform 1 0 2576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2709__CLK
timestamp 1698431365
transform 1 0 2016 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2710__CLK
timestamp 1698431365
transform 1 0 5488 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2711__CLK
timestamp 1698431365
transform 1 0 4592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2712__CLK
timestamp 1698431365
transform 1 0 2128 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2713__CLK
timestamp 1698431365
transform 1 0 4032 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2714__CLK
timestamp 1698431365
transform 1 0 16352 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2716__CLK
timestamp 1698431365
transform 1 0 36064 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 25536 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_0_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 19264 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_1_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 18816 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_2_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 21616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_3_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 24752 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_4_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 15792 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_5_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 15344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_6_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 15792 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_7_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 20720 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_8_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_9_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 37744 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_10_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 39984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_11_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 40992 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_12_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 35952 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_13_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 33824 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_14_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 38080 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_15_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 42672 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 41328 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 40880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 48384 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 47712 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 45136 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 47936 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 44016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform 1 0 1792 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 1792 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output15_I
timestamp 1698431365
transform 1 0 30912 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output16_I
timestamp 1698431365
transform -1 0 23072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_rebuffer10_I
timestamp 1698431365
transform -1 0 16352 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_rebuffer20_I
timestamp 1698431365
transform -1 0 12656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_0_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16240 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_1_0_wb_clk_i
timestamp 1698431365
transform 1 0 14112 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_2_0_wb_clk_i
timestamp 1698431365
transform -1 0 21280 0 -1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_3_0_wb_clk_i
timestamp 1698431365
transform 1 0 19376 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_4_0_wb_clk_i
timestamp 1698431365
transform -1 0 15568 0 -1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_5_0_wb_clk_i
timestamp 1698431365
transform -1 0 15120 0 -1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_6_0_wb_clk_i
timestamp 1698431365
transform 1 0 18032 0 -1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_7_0_wb_clk_i
timestamp 1698431365
transform -1 0 20496 0 -1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_8_0_wb_clk_i
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_9_0_wb_clk_i
timestamp 1698431365
transform -1 0 39760 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_10_0_wb_clk_i
timestamp 1698431365
transform -1 0 42672 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_11_0_wb_clk_i
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_12_0_wb_clk_i
timestamp 1698431365
transform 1 0 36960 0 -1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_13_0_wb_clk_i
timestamp 1698431365
transform 1 0 34048 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_14_0_wb_clk_i
timestamp 1698431365
transform 1 0 40096 0 1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_15_0_wb_clk_i
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_36 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_46 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6496 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_50
timestamp 1698431365
transform 1 0 6944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_58 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7840 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_64
timestamp 1698431365
transform 1 0 8512 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_74
timestamp 1698431365
transform 1 0 9632 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_78
timestamp 1698431365
transform 1 0 10080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_82
timestamp 1698431365
transform 1 0 10528 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_86
timestamp 1698431365
transform 1 0 10976 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_90
timestamp 1698431365
transform 1 0 11424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_94
timestamp 1698431365
transform 1 0 11872 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_98
timestamp 1698431365
transform 1 0 12320 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_108
timestamp 1698431365
transform 1 0 13440 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_112 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_115
timestamp 1698431365
transform 1 0 14224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_119
timestamp 1698431365
transform 1 0 14672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_123
timestamp 1698431365
transform 1 0 15120 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_127
timestamp 1698431365
transform 1 0 15568 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_130
timestamp 1698431365
transform 1 0 15904 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_144
timestamp 1698431365
transform 1 0 17472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_148
timestamp 1698431365
transform 1 0 17920 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_150
timestamp 1698431365
transform 1 0 18144 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_153
timestamp 1698431365
transform 1 0 18480 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_157
timestamp 1698431365
transform 1 0 18928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_165
timestamp 1698431365
transform 1 0 19824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698431365
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698431365
transform 1 0 21056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_180
timestamp 1698431365
transform 1 0 21504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_188
timestamp 1698431365
transform 1 0 22400 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_192
timestamp 1698431365
transform 1 0 22848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_196
timestamp 1698431365
transform 1 0 23296 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_200
timestamp 1698431365
transform 1 0 23744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_235
timestamp 1698431365
transform 1 0 27664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698431365
transform 1 0 27888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_244 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28672 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_260
timestamp 1698431365
transform 1 0 30464 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_268
timestamp 1698431365
transform 1 0 31360 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_290
timestamp 1698431365
transform 1 0 33824 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_298
timestamp 1698431365
transform 1 0 34720 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_302
timestamp 1698431365
transform 1 0 35168 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_337
timestamp 1698431365
transform 1 0 39088 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_339
timestamp 1698431365
transform 1 0 39312 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_371
timestamp 1698431365
transform 1 0 42896 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_373
timestamp 1698431365
transform 1 0 43120 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_376
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_380
timestamp 1698431365
transform 1 0 43904 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_388
timestamp 1698431365
transform 1 0 44800 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_391
timestamp 1698431365
transform 1 0 45136 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_399
timestamp 1698431365
transform 1 0 46032 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_403
timestamp 1698431365
transform 1 0 46480 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_405
timestamp 1698431365
transform 1 0 46704 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_410
timestamp 1698431365
transform 1 0 47264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_2
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_34
timestamp 1698431365
transform 1 0 5152 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_37
timestamp 1698431365
transform 1 0 5488 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_201
timestamp 1698431365
transform 1 0 23856 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_205
timestamp 1698431365
transform 1 0 24304 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698431365
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_216
timestamp 1698431365
transform 1 0 25536 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_220
timestamp 1698431365
transform 1 0 25984 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_224
timestamp 1698431365
transform 1 0 26432 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_226
timestamp 1698431365
transform 1 0 26656 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_229
timestamp 1698431365
transform 1 0 26992 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_260
timestamp 1698431365
transform 1 0 30464 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_264
timestamp 1698431365
transform 1 0 30912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698431365
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_344
timestamp 1698431365
transform 1 0 39872 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_348
timestamp 1698431365
transform 1 0 40320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_387
timestamp 1698431365
transform 1 0 44688 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_18
timestamp 1698431365
transform 1 0 3360 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_26
timestamp 1698431365
transform 1 0 4256 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_28
timestamp 1698431365
transform 1 0 4480 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_31
timestamp 1698431365
transform 1 0 4816 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_41
timestamp 1698431365
transform 1 0 5936 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_43
timestamp 1698431365
transform 1 0 6160 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_64
timestamp 1698431365
transform 1 0 8512 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_102
timestamp 1698431365
transform 1 0 12768 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_104
timestamp 1698431365
transform 1 0 12992 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_119
timestamp 1698431365
transform 1 0 14672 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_123
timestamp 1698431365
transform 1 0 15120 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_153
timestamp 1698431365
transform 1 0 18480 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_157
timestamp 1698431365
transform 1 0 18928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_161
timestamp 1698431365
transform 1 0 19376 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_174
timestamp 1698431365
transform 1 0 20832 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_181
timestamp 1698431365
transform 1 0 21616 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_183
timestamp 1698431365
transform 1 0 21840 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_255
timestamp 1698431365
transform 1 0 29904 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_304
timestamp 1698431365
transform 1 0 35392 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_312
timestamp 1698431365
transform 1 0 36288 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_314
timestamp 1698431365
transform 1 0 36512 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_321
timestamp 1698431365
transform 1 0 37296 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_329
timestamp 1698431365
transform 1 0 38192 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_333
timestamp 1698431365
transform 1 0 38640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_370
timestamp 1698431365
transform 1 0 42784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_374
timestamp 1698431365
transform 1 0 43232 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_384
timestamp 1698431365
transform 1 0 44352 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_391
timestamp 1698431365
transform 1 0 45136 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_395
timestamp 1698431365
transform 1 0 45584 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_416
timestamp 1698431365
transform 1 0 47936 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_18
timestamp 1698431365
transform 1 0 3360 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_93
timestamp 1698431365
transform 1 0 11760 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_123
timestamp 1698431365
transform 1 0 15120 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_151
timestamp 1698431365
transform 1 0 18256 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_153
timestamp 1698431365
transform 1 0 18480 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_170
timestamp 1698431365
transform 1 0 20384 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_198
timestamp 1698431365
transform 1 0 23520 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_226
timestamp 1698431365
transform 1 0 26656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_228
timestamp 1698431365
transform 1 0 26880 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_253
timestamp 1698431365
transform 1 0 29680 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_275
timestamp 1698431365
transform 1 0 32144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_277
timestamp 1698431365
transform 1 0 32368 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_300
timestamp 1698431365
transform 1 0 34944 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_304
timestamp 1698431365
transform 1 0 35392 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_318
timestamp 1698431365
transform 1 0 36960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_322
timestamp 1698431365
transform 1 0 37408 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_326
timestamp 1698431365
transform 1 0 37856 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_334
timestamp 1698431365
transform 1 0 38752 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_344
timestamp 1698431365
transform 1 0 39872 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_348
timestamp 1698431365
transform 1 0 40320 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_382
timestamp 1698431365
transform 1 0 44128 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_388
timestamp 1698431365
transform 1 0 44800 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_390
timestamp 1698431365
transform 1 0 45024 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_10
timestamp 1698431365
transform 1 0 2464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_12
timestamp 1698431365
transform 1 0 2688 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_15
timestamp 1698431365
transform 1 0 3024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_19
timestamp 1698431365
transform 1 0 3472 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_23
timestamp 1698431365
transform 1 0 3920 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_27
timestamp 1698431365
transform 1 0 4368 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_31
timestamp 1698431365
transform 1 0 4816 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_55
timestamp 1698431365
transform 1 0 7504 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_97
timestamp 1698431365
transform 1 0 12208 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_158
timestamp 1698431365
transform 1 0 19040 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_160
timestamp 1698431365
transform 1 0 19264 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_181
timestamp 1698431365
transform 1 0 21616 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_190
timestamp 1698431365
transform 1 0 22624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_194
timestamp 1698431365
transform 1 0 23072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_239
timestamp 1698431365
transform 1 0 28112 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_243
timestamp 1698431365
transform 1 0 28560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_253
timestamp 1698431365
transform 1 0 29680 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_265
timestamp 1698431365
transform 1 0 31024 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_290
timestamp 1698431365
transform 1 0 33824 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_297
timestamp 1698431365
transform 1 0 34608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_301
timestamp 1698431365
transform 1 0 35056 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_314
timestamp 1698431365
transform 1 0 36512 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_351
timestamp 1698431365
transform 1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_355
timestamp 1698431365
transform 1 0 41104 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_395
timestamp 1698431365
transform 1 0 45584 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_397
timestamp 1698431365
transform 1 0 45808 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_416
timestamp 1698431365
transform 1 0 47936 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_6
timestamp 1698431365
transform 1 0 2016 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_10
timestamp 1698431365
transform 1 0 2464 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_13
timestamp 1698431365
transform 1 0 2800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_62
timestamp 1698431365
transform 1 0 8288 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_125
timestamp 1698431365
transform 1 0 15344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_127
timestamp 1698431365
transform 1 0 15568 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_132
timestamp 1698431365
transform 1 0 16128 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_150
timestamp 1698431365
transform 1 0 18144 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_154
timestamp 1698431365
transform 1 0 18592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_158
timestamp 1698431365
transform 1 0 19040 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_180
timestamp 1698431365
transform 1 0 21504 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_182
timestamp 1698431365
transform 1 0 21728 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_195
timestamp 1698431365
transform 1 0 23184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_199
timestamp 1698431365
transform 1 0 23632 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_209
timestamp 1698431365
transform 1 0 24752 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_220
timestamp 1698431365
transform 1 0 25984 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_279
timestamp 1698431365
transform 1 0 32592 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_296
timestamp 1698431365
transform 1 0 34496 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_300
timestamp 1698431365
transform 1 0 34944 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_323
timestamp 1698431365
transform 1 0 37520 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_340
timestamp 1698431365
transform 1 0 39424 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_372
timestamp 1698431365
transform 1 0 43008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_376
timestamp 1698431365
transform 1 0 43456 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_393
timestamp 1698431365
transform 1 0 45360 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_397
timestamp 1698431365
transform 1 0 45808 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_401
timestamp 1698431365
transform 1 0 46256 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_403
timestamp 1698431365
transform 1 0 46480 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_6
timestamp 1698431365
transform 1 0 2016 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_10
timestamp 1698431365
transform 1 0 2464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_14
timestamp 1698431365
transform 1 0 2912 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_18
timestamp 1698431365
transform 1 0 3360 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_22
timestamp 1698431365
transform 1 0 3808 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_26
timestamp 1698431365
transform 1 0 4256 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_41
timestamp 1698431365
transform 1 0 5936 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_43
timestamp 1698431365
transform 1 0 6160 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_76
timestamp 1698431365
transform 1 0 9856 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_172
timestamp 1698431365
transform 1 0 20608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_174
timestamp 1698431365
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_182
timestamp 1698431365
transform 1 0 21728 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_186
timestamp 1698431365
transform 1 0 22176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_241
timestamp 1698431365
transform 1 0 28336 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_261
timestamp 1698431365
transform 1 0 30576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_265
timestamp 1698431365
transform 1 0 31024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_269
timestamp 1698431365
transform 1 0 31472 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_273
timestamp 1698431365
transform 1 0 31920 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_345
timestamp 1698431365
transform 1 0 39984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_349
timestamp 1698431365
transform 1 0 40432 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_351
timestamp 1698431365
transform 1 0 40656 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_380
timestamp 1698431365
transform 1 0 43904 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_384
timestamp 1698431365
transform 1 0 44352 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_4
timestamp 1698431365
transform 1 0 1792 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_7
timestamp 1698431365
transform 1 0 2128 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_11
timestamp 1698431365
transform 1 0 2576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_15
timestamp 1698431365
transform 1 0 3024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_48
timestamp 1698431365
transform 1 0 6720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_50
timestamp 1698431365
transform 1 0 6944 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_69
timestamp 1698431365
transform 1 0 9072 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_79
timestamp 1698431365
transform 1 0 10192 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_125
timestamp 1698431365
transform 1 0 15344 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_129
timestamp 1698431365
transform 1 0 15792 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_132
timestamp 1698431365
transform 1 0 16128 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_136
timestamp 1698431365
transform 1 0 16576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_148
timestamp 1698431365
transform 1 0 17920 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_189
timestamp 1698431365
transform 1 0 22512 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_193
timestamp 1698431365
transform 1 0 22960 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_198
timestamp 1698431365
transform 1 0 23520 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_200
timestamp 1698431365
transform 1 0 23744 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_203
timestamp 1698431365
transform 1 0 24080 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_205
timestamp 1698431365
transform 1 0 24304 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_208
timestamp 1698431365
transform 1 0 24640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_216
timestamp 1698431365
transform 1 0 25536 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_222
timestamp 1698431365
transform 1 0 26208 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_226
timestamp 1698431365
transform 1 0 26656 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_233
timestamp 1698431365
transform 1 0 27440 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_237
timestamp 1698431365
transform 1 0 27888 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_241
timestamp 1698431365
transform 1 0 28336 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_245
timestamp 1698431365
transform 1 0 28784 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_247
timestamp 1698431365
transform 1 0 29008 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_258
timestamp 1698431365
transform 1 0 30240 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_276
timestamp 1698431365
transform 1 0 32256 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_313
timestamp 1698431365
transform 1 0 36400 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_317
timestamp 1698431365
transform 1 0 36848 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_321
timestamp 1698431365
transform 1 0 37296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_339
timestamp 1698431365
transform 1 0 39312 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_341
timestamp 1698431365
transform 1 0 39536 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_357
timestamp 1698431365
transform 1 0 41328 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_394
timestamp 1698431365
transform 1 0 45472 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_398
timestamp 1698431365
transform 1 0 45920 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_400
timestamp 1698431365
transform 1 0 46144 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_418
timestamp 1698431365
transform 1 0 48160 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_4
timestamp 1698431365
transform 1 0 1792 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_7
timestamp 1698431365
transform 1 0 2128 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_11
timestamp 1698431365
transform 1 0 2576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_15
timestamp 1698431365
transform 1 0 3024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_19
timestamp 1698431365
transform 1 0 3472 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_23
timestamp 1698431365
transform 1 0 3920 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_27
timestamp 1698431365
transform 1 0 4368 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_31
timestamp 1698431365
transform 1 0 4816 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_41
timestamp 1698431365
transform 1 0 5936 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_44
timestamp 1698431365
transform 1 0 6272 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_48
timestamp 1698431365
transform 1 0 6720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_65
timestamp 1698431365
transform 1 0 8624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_67
timestamp 1698431365
transform 1 0 8848 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_73
timestamp 1698431365
transform 1 0 9520 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_79
timestamp 1698431365
transform 1 0 10192 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_83
timestamp 1698431365
transform 1 0 10640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_85
timestamp 1698431365
transform 1 0 10864 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_88
timestamp 1698431365
transform 1 0 11200 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_90
timestamp 1698431365
transform 1 0 11424 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_93
timestamp 1698431365
transform 1 0 11760 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_97
timestamp 1698431365
transform 1 0 12208 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_109
timestamp 1698431365
transform 1 0 13552 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_115
timestamp 1698431365
transform 1 0 14224 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_119
timestamp 1698431365
transform 1 0 14672 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_122
timestamp 1698431365
transform 1 0 15008 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_155
timestamp 1698431365
transform 1 0 18704 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_159
timestamp 1698431365
transform 1 0 19152 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_163
timestamp 1698431365
transform 1 0 19600 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_170
timestamp 1698431365
transform 1 0 20384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_172
timestamp 1698431365
transform 1 0 20608 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_179
timestamp 1698431365
transform 1 0 21392 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_244
timestamp 1698431365
transform 1 0 28672 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_305
timestamp 1698431365
transform 1 0 35504 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_325
timestamp 1698431365
transform 1 0 37744 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_378
timestamp 1698431365
transform 1 0 43680 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_8
timestamp 1698431365
transform 1 0 2240 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_12
timestamp 1698431365
transform 1 0 2688 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_16
timestamp 1698431365
transform 1 0 3136 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_57
timestamp 1698431365
transform 1 0 7728 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_59
timestamp 1698431365
transform 1 0 7952 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_62
timestamp 1698431365
transform 1 0 8288 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_103
timestamp 1698431365
transform 1 0 12880 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_128
timestamp 1698431365
transform 1 0 15680 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_144
timestamp 1698431365
transform 1 0 17472 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_167
timestamp 1698431365
transform 1 0 20048 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_204
timestamp 1698431365
transform 1 0 24192 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_208
timestamp 1698431365
transform 1 0 24640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_228
timestamp 1698431365
transform 1 0 26880 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_259
timestamp 1698431365
transform 1 0 30352 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_268
timestamp 1698431365
transform 1 0 31360 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_272
timestamp 1698431365
transform 1 0 31808 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_275
timestamp 1698431365
transform 1 0 32144 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_279
timestamp 1698431365
transform 1 0 32592 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_286
timestamp 1698431365
transform 1 0 33376 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_290
timestamp 1698431365
transform 1 0 33824 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_297
timestamp 1698431365
transform 1 0 34608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_301
timestamp 1698431365
transform 1 0 35056 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_316
timestamp 1698431365
transform 1 0 36736 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_320
timestamp 1698431365
transform 1 0 37184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_340
timestamp 1698431365
transform 1 0 39424 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_394
timestamp 1698431365
transform 1 0 45472 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_398
timestamp 1698431365
transform 1 0 45920 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_412
timestamp 1698431365
transform 1 0 47488 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_84
timestamp 1698431365
transform 1 0 10752 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_103
timestamp 1698431365
transform 1 0 12880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_143
timestamp 1698431365
transform 1 0 17360 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_173
timestamp 1698431365
transform 1 0 20720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_199
timestamp 1698431365
transform 1 0 23632 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_203
timestamp 1698431365
transform 1 0 24080 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_207
timestamp 1698431365
transform 1 0 24528 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_217
timestamp 1698431365
transform 1 0 25648 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_221
timestamp 1698431365
transform 1 0 26096 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_225
timestamp 1698431365
transform 1 0 26544 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_234
timestamp 1698431365
transform 1 0 27552 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_238
timestamp 1698431365
transform 1 0 28000 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_242
timestamp 1698431365
transform 1 0 28448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_244
timestamp 1698431365
transform 1 0 28672 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_251
timestamp 1698431365
transform 1 0 29456 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_255
timestamp 1698431365
transform 1 0 29904 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_259
timestamp 1698431365
transform 1 0 30352 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_325
timestamp 1698431365
transform 1 0 37744 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_329
timestamp 1698431365
transform 1 0 38192 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_333
timestamp 1698431365
transform 1 0 38640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_337
timestamp 1698431365
transform 1 0 39088 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_345
timestamp 1698431365
transform 1 0 39984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_370
timestamp 1698431365
transform 1 0 42784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_374
timestamp 1698431365
transform 1 0 43232 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_378
timestamp 1698431365
transform 1 0 43680 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_382
timestamp 1698431365
transform 1 0 44128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_384
timestamp 1698431365
transform 1 0 44352 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_415
timestamp 1698431365
transform 1 0 47824 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_419
timestamp 1698431365
transform 1 0 48272 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_6
timestamp 1698431365
transform 1 0 2016 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_10
timestamp 1698431365
transform 1 0 2464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_43
timestamp 1698431365
transform 1 0 6160 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_61
timestamp 1698431365
transform 1 0 8176 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_63
timestamp 1698431365
transform 1 0 8400 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_88
timestamp 1698431365
transform 1 0 11200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_110
timestamp 1698431365
transform 1 0 13664 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_129
timestamp 1698431365
transform 1 0 15792 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_131
timestamp 1698431365
transform 1 0 16016 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_230
timestamp 1698431365
transform 1 0 27104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_232
timestamp 1698431365
transform 1 0 27328 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_257
timestamp 1698431365
transform 1 0 30128 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_259
timestamp 1698431365
transform 1 0 30352 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_277
timestamp 1698431365
transform 1 0 32368 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_279
timestamp 1698431365
transform 1 0 32592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_290
timestamp 1698431365
transform 1 0 33824 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_345
timestamp 1698431365
transform 1 0 39984 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_349
timestamp 1698431365
transform 1 0 40432 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_364
timestamp 1698431365
transform 1 0 42112 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_368
timestamp 1698431365
transform 1 0 42560 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_372
timestamp 1698431365
transform 1 0 43008 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_380
timestamp 1698431365
transform 1 0 43904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_384
timestamp 1698431365
transform 1 0 44352 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_388
timestamp 1698431365
transform 1 0 44800 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_4
timestamp 1698431365
transform 1 0 1792 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_7
timestamp 1698431365
transform 1 0 2128 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_11
timestamp 1698431365
transform 1 0 2576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_15
timestamp 1698431365
transform 1 0 3024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_19
timestamp 1698431365
transform 1 0 3472 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_23
timestamp 1698431365
transform 1 0 3920 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_27
timestamp 1698431365
transform 1 0 4368 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_31
timestamp 1698431365
transform 1 0 4816 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_78
timestamp 1698431365
transform 1 0 10080 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_102
timestamp 1698431365
transform 1 0 12768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1698431365
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_109
timestamp 1698431365
transform 1 0 13552 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_144
timestamp 1698431365
transform 1 0 17472 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_179
timestamp 1698431365
transform 1 0 21392 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_201
timestamp 1698431365
transform 1 0 23856 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_234
timestamp 1698431365
transform 1 0 27552 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_236
timestamp 1698431365
transform 1 0 27776 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_276
timestamp 1698431365
transform 1 0 32256 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_280
timestamp 1698431365
transform 1 0 32704 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_282
timestamp 1698431365
transform 1 0 32928 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_314
timestamp 1698431365
transform 1 0 36512 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_321
timestamp 1698431365
transform 1 0 37296 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_323
timestamp 1698431365
transform 1 0 37520 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_382
timestamp 1698431365
transform 1 0 44128 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_384
timestamp 1698431365
transform 1 0 44352 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_393
timestamp 1698431365
transform 1 0 45360 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_395
timestamp 1698431365
transform 1 0 45584 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_401
timestamp 1698431365
transform 1 0 46256 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_410
timestamp 1698431365
transform 1 0 47264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_6
timestamp 1698431365
transform 1 0 2016 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_9
timestamp 1698431365
transform 1 0 2352 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_13
timestamp 1698431365
transform 1 0 2800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_118
timestamp 1698431365
transform 1 0 14560 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_206
timestamp 1698431365
transform 1 0 24416 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_214
timestamp 1698431365
transform 1 0 25312 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_223
timestamp 1698431365
transform 1 0 26320 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_227
timestamp 1698431365
transform 1 0 26768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_231
timestamp 1698431365
transform 1 0 27216 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_235
timestamp 1698431365
transform 1 0 27664 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_239
timestamp 1698431365
transform 1 0 28112 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_243
timestamp 1698431365
transform 1 0 28560 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_247
timestamp 1698431365
transform 1 0 29008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_251
timestamp 1698431365
transform 1 0 29456 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_261
timestamp 1698431365
transform 1 0 30576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_265
timestamp 1698431365
transform 1 0 31024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_277
timestamp 1698431365
transform 1 0 32368 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698431365
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_327
timestamp 1698431365
transform 1 0 37968 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_345
timestamp 1698431365
transform 1 0 39984 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_349
timestamp 1698431365
transform 1 0 40432 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_356
timestamp 1698431365
transform 1 0 41216 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_363
timestamp 1698431365
transform 1 0 42000 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_371
timestamp 1698431365
transform 1 0 42896 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_383
timestamp 1698431365
transform 1 0 44240 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_391
timestamp 1698431365
transform 1 0 45136 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_399
timestamp 1698431365
transform 1 0 46032 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_416
timestamp 1698431365
transform 1 0 47936 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_6
timestamp 1698431365
transform 1 0 2016 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_10
timestamp 1698431365
transform 1 0 2464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_14
timestamp 1698431365
transform 1 0 2912 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_18
timestamp 1698431365
transform 1 0 3360 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_22
timestamp 1698431365
transform 1 0 3808 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_26
timestamp 1698431365
transform 1 0 4256 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_113
timestamp 1698431365
transform 1 0 14000 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_130
timestamp 1698431365
transform 1 0 15904 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_132
timestamp 1698431365
transform 1 0 16128 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_144
timestamp 1698431365
transform 1 0 17472 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_206
timestamp 1698431365
transform 1 0 24416 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_228
timestamp 1698431365
transform 1 0 26880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_232
timestamp 1698431365
transform 1 0 27328 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_236
timestamp 1698431365
transform 1 0 27776 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_240
timestamp 1698431365
transform 1 0 28224 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_255
timestamp 1698431365
transform 1 0 29904 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_306
timestamp 1698431365
transform 1 0 35616 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_310
timestamp 1698431365
transform 1 0 36064 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_314
timestamp 1698431365
transform 1 0 36512 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_323
timestamp 1698431365
transform 1 0 37520 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_327
timestamp 1698431365
transform 1 0 37968 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_331
timestamp 1698431365
transform 1 0 38416 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_333
timestamp 1698431365
transform 1 0 38640 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_345
timestamp 1698431365
transform 1 0 39984 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_355
timestamp 1698431365
transform 1 0 41104 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_6
timestamp 1698431365
transform 1 0 2016 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_9
timestamp 1698431365
transform 1 0 2352 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_13
timestamp 1698431365
transform 1 0 2800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_17
timestamp 1698431365
transform 1 0 3248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_69
timestamp 1698431365
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_74
timestamp 1698431365
transform 1 0 9632 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_102
timestamp 1698431365
transform 1 0 12768 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_179
timestamp 1698431365
transform 1 0 21392 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698431365
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_278
timestamp 1698431365
transform 1 0 32480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_307
timestamp 1698431365
transform 1 0 35728 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_311
timestamp 1698431365
transform 1 0 36176 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_315
timestamp 1698431365
transform 1 0 36624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_319
timestamp 1698431365
transform 1 0 37072 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_323
timestamp 1698431365
transform 1 0 37520 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_327
timestamp 1698431365
transform 1 0 37968 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_331
timestamp 1698431365
transform 1 0 38416 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_335
timestamp 1698431365
transform 1 0 38864 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_339
timestamp 1698431365
transform 1 0 39312 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_347
timestamp 1698431365
transform 1 0 40208 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_349
timestamp 1698431365
transform 1 0 40432 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_378
timestamp 1698431365
transform 1 0 43680 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_385
timestamp 1698431365
transform 1 0 44464 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_395
timestamp 1698431365
transform 1 0 45584 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_402
timestamp 1698431365
transform 1 0 46368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_404
timestamp 1698431365
transform 1 0 46592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_6
timestamp 1698431365
transform 1 0 2016 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_9
timestamp 1698431365
transform 1 0 2352 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_13
timestamp 1698431365
transform 1 0 2800 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_17
timestamp 1698431365
transform 1 0 3248 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_21
timestamp 1698431365
transform 1 0 3696 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_39
timestamp 1698431365
transform 1 0 5712 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_50
timestamp 1698431365
transform 1 0 6944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_60
timestamp 1698431365
transform 1 0 8064 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_90
timestamp 1698431365
transform 1 0 11424 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_92
timestamp 1698431365
transform 1 0 11648 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_103
timestamp 1698431365
transform 1 0 12880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_189
timestamp 1698431365
transform 1 0 22512 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_191
timestamp 1698431365
transform 1 0 22736 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_223
timestamp 1698431365
transform 1 0 26320 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_231
timestamp 1698431365
transform 1 0 27216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_255
timestamp 1698431365
transform 1 0 29904 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_265
timestamp 1698431365
transform 1 0 31024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_277
timestamp 1698431365
transform 1 0 32368 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_321
timestamp 1698431365
transform 1 0 37296 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_375
timestamp 1698431365
transform 1 0 43344 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_381
timestamp 1698431365
transform 1 0 44016 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_18
timestamp 1698431365
transform 1 0 3360 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_35
timestamp 1698431365
transform 1 0 5264 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698431365
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_160
timestamp 1698431365
transform 1 0 19264 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_220
timestamp 1698431365
transform 1 0 25984 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_246
timestamp 1698431365
transform 1 0 28896 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698431365
transform 1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698431365
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_308
timestamp 1698431365
transform 1 0 35840 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_349
timestamp 1698431365
transform 1 0 40432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_418
timestamp 1698431365
transform 1 0 48160 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_11
timestamp 1698431365
transform 1 0 2576 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_15
timestamp 1698431365
transform 1 0 3024 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_26
timestamp 1698431365
transform 1 0 4256 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_39
timestamp 1698431365
transform 1 0 5712 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_191
timestamp 1698431365
transform 1 0 22736 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_203
timestamp 1698431365
transform 1 0 24080 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_253
timestamp 1698431365
transform 1 0 29680 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_299
timestamp 1698431365
transform 1 0 34832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_303
timestamp 1698431365
transform 1 0 35280 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_312
timestamp 1698431365
transform 1 0 36288 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_314
timestamp 1698431365
transform 1 0 36512 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_379
timestamp 1698431365
transform 1 0 43792 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_383
timestamp 1698431365
transform 1 0 44240 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_410
timestamp 1698431365
transform 1 0 47264 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_417
timestamp 1698431365
transform 1 0 48048 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_419
timestamp 1698431365
transform 1 0 48272 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_109
timestamp 1698431365
transform 1 0 13552 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698431365
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_182
timestamp 1698431365
transform 1 0 21728 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_184
timestamp 1698431365
transform 1 0 21952 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_249
timestamp 1698431365
transform 1 0 29232 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_317
timestamp 1698431365
transform 1 0 36848 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_321
timestamp 1698431365
transform 1 0 37296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_323
timestamp 1698431365
transform 1 0 37520 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_332
timestamp 1698431365
transform 1 0 38528 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_412
timestamp 1698431365
transform 1 0 47488 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_31
timestamp 1698431365
transform 1 0 4816 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_47
timestamp 1698431365
transform 1 0 6608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_49
timestamp 1698431365
transform 1 0 6832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_60
timestamp 1698431365
transform 1 0 8064 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_90
timestamp 1698431365
transform 1 0 11424 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698431365
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_242
timestamp 1698431365
transform 1 0 28448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698431365
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_302
timestamp 1698431365
transform 1 0 35168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_306
timestamp 1698431365
transform 1 0 35616 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_310
timestamp 1698431365
transform 1 0 36064 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698431365
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_375
timestamp 1698431365
transform 1 0 43344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_6
timestamp 1698431365
transform 1 0 2016 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_69
timestamp 1698431365
transform 1 0 9072 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_89
timestamp 1698431365
transform 1 0 11312 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_217
timestamp 1698431365
transform 1 0 25648 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_267
timestamp 1698431365
transform 1 0 31248 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_300
timestamp 1698431365
transform 1 0 34944 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_304
timestamp 1698431365
transform 1 0 35392 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_308
timestamp 1698431365
transform 1 0 35840 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_312
timestamp 1698431365
transform 1 0 36288 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_316
timestamp 1698431365
transform 1 0 36736 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_318
timestamp 1698431365
transform 1 0 36960 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_339
timestamp 1698431365
transform 1 0 39312 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_343
timestamp 1698431365
transform 1 0 39760 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_347
timestamp 1698431365
transform 1 0 40208 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_349
timestamp 1698431365
transform 1 0 40432 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_356
timestamp 1698431365
transform 1 0 41216 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_358
timestamp 1698431365
transform 1 0 41440 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_398
timestamp 1698431365
transform 1 0 45920 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_400
timestamp 1698431365
transform 1 0 46144 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_418
timestamp 1698431365
transform 1 0 48160 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_33
timestamp 1698431365
transform 1 0 5040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_90
timestamp 1698431365
transform 1 0 11424 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_193
timestamp 1698431365
transform 1 0 22960 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_232
timestamp 1698431365
transform 1 0 27328 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698431365
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_280
timestamp 1698431365
transform 1 0 32704 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_282
timestamp 1698431365
transform 1 0 32928 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_323
timestamp 1698431365
transform 1 0 37520 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_333
timestamp 1698431365
transform 1 0 38640 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_372
timestamp 1698431365
transform 1 0 43008 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_380
timestamp 1698431365
transform 1 0 43904 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_382
timestamp 1698431365
transform 1 0 44128 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_387
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_33
timestamp 1698431365
transform 1 0 5040 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_81
timestamp 1698431365
transform 1 0 10416 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_83
timestamp 1698431365
transform 1 0 10640 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698431365
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_192
timestamp 1698431365
transform 1 0 22848 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_194
timestamp 1698431365
transform 1 0 23072 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_257
timestamp 1698431365
transform 1 0 30128 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_266
timestamp 1698431365
transform 1 0 31136 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_290
timestamp 1698431365
transform 1 0 33824 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_328
timestamp 1698431365
transform 1 0 38080 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_332
timestamp 1698431365
transform 1 0 38528 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_345
timestamp 1698431365
transform 1 0 39984 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_349
timestamp 1698431365
transform 1 0 40432 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_358
timestamp 1698431365
transform 1 0 41440 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_363
timestamp 1698431365
transform 1 0 42000 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_367
timestamp 1698431365
transform 1 0 42448 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_371
timestamp 1698431365
transform 1 0 42896 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_402
timestamp 1698431365
transform 1 0 46368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_47
timestamp 1698431365
transform 1 0 6608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_49
timestamp 1698431365
transform 1 0 6832 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_94
timestamp 1698431365
transform 1 0 11872 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_96
timestamp 1698431365
transform 1 0 12096 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_121
timestamp 1698431365
transform 1 0 14896 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_163
timestamp 1698431365
transform 1 0 19600 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_172
timestamp 1698431365
transform 1 0 20608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698431365
transform 1 0 20832 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_241
timestamp 1698431365
transform 1 0 28336 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_305
timestamp 1698431365
transform 1 0 35504 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_353
timestamp 1698431365
transform 1 0 40880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_357
timestamp 1698431365
transform 1 0 41328 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_384
timestamp 1698431365
transform 1 0 44352 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_417
timestamp 1698431365
transform 1 0 48048 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_419
timestamp 1698431365
transform 1 0 48272 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_38
timestamp 1698431365
transform 1 0 5600 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_86
timestamp 1698431365
transform 1 0 10976 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_183
timestamp 1698431365
transform 1 0 21840 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_185
timestamp 1698431365
transform 1 0 22064 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_222
timestamp 1698431365
transform 1 0 26208 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_276
timestamp 1698431365
transform 1 0 32256 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_298
timestamp 1698431365
transform 1 0 34720 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_300
timestamp 1698431365
transform 1 0 34944 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_309
timestamp 1698431365
transform 1 0 35952 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_313
timestamp 1698431365
transform 1 0 36400 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_317
timestamp 1698431365
transform 1 0 36848 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_321
timestamp 1698431365
transform 1 0 37296 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_325
timestamp 1698431365
transform 1 0 37744 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_340
timestamp 1698431365
transform 1 0 39424 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_348
timestamp 1698431365
transform 1 0 40320 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_387
timestamp 1698431365
transform 1 0 44688 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_403
timestamp 1698431365
transform 1 0 46480 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_51
timestamp 1698431365
transform 1 0 7056 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_53
timestamp 1698431365
transform 1 0 7280 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_102
timestamp 1698431365
transform 1 0 12768 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_104
timestamp 1698431365
transform 1 0 12992 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_158
timestamp 1698431365
transform 1 0 19040 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_160
timestamp 1698431365
transform 1 0 19264 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_192
timestamp 1698431365
transform 1 0 22848 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_216
timestamp 1698431365
transform 1 0 25536 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_218
timestamp 1698431365
transform 1 0 25760 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_266
timestamp 1698431365
transform 1 0 31136 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_278
timestamp 1698431365
transform 1 0 32480 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698431365
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_331
timestamp 1698431365
transform 1 0 38416 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_339
timestamp 1698431365
transform 1 0 39312 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_343
timestamp 1698431365
transform 1 0 39760 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_353
timestamp 1698431365
transform 1 0 40880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_357
timestamp 1698431365
transform 1 0 41328 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_378
timestamp 1698431365
transform 1 0 43680 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_382
timestamp 1698431365
transform 1 0 44128 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_384
timestamp 1698431365
transform 1 0 44352 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_42
timestamp 1698431365
transform 1 0 6048 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_80
timestamp 1698431365
transform 1 0 10304 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_186
timestamp 1698431365
transform 1 0 22176 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_188
timestamp 1698431365
transform 1 0 22400 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_262
timestamp 1698431365
transform 1 0 30688 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_276
timestamp 1698431365
transform 1 0 32256 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_303
timestamp 1698431365
transform 1 0 35280 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_360
timestamp 1698431365
transform 1 0 41664 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_418
timestamp 1698431365
transform 1 0 48160 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_31
timestamp 1698431365
transform 1 0 4816 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_218
timestamp 1698431365
transform 1 0 25760 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_292
timestamp 1698431365
transform 1 0 34048 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_307
timestamp 1698431365
transform 1 0 35728 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_311
timestamp 1698431365
transform 1 0 36176 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_325
timestamp 1698431365
transform 1 0 37744 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_333
timestamp 1698431365
transform 1 0 38640 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_357
timestamp 1698431365
transform 1 0 41328 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_364
timestamp 1698431365
transform 1 0 42112 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_372
timestamp 1698431365
transform 1 0 43008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_374
timestamp 1698431365
transform 1 0 43232 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_377
timestamp 1698431365
transform 1 0 43568 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_381
timestamp 1698431365
transform 1 0 44016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_399
timestamp 1698431365
transform 1 0 46032 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_416
timestamp 1698431365
transform 1 0 47936 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_33
timestamp 1698431365
transform 1 0 5040 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_74
timestamp 1698431365
transform 1 0 9632 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_138
timestamp 1698431365
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_207
timestamp 1698431365
transform 1 0 24528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698431365
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698431365
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_290
timestamp 1698431365
transform 1 0 33824 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_338
timestamp 1698431365
transform 1 0 39200 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_343
timestamp 1698431365
transform 1 0 39760 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_347
timestamp 1698431365
transform 1 0 40208 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_349
timestamp 1698431365
transform 1 0 40432 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_360
timestamp 1698431365
transform 1 0 41664 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_382
timestamp 1698431365
transform 1 0 44128 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_88
timestamp 1698431365
transform 1 0 11200 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_90
timestamp 1698431365
transform 1 0 11424 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_236
timestamp 1698431365
transform 1 0 27776 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_255
timestamp 1698431365
transform 1 0 29904 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_269
timestamp 1698431365
transform 1 0 31472 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_273
timestamp 1698431365
transform 1 0 31920 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_303
timestamp 1698431365
transform 1 0 35280 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698431365
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_355
timestamp 1698431365
transform 1 0 41104 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_387
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_31
timestamp 1698431365
transform 1 0 4816 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_51
timestamp 1698431365
transform 1 0 7056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_108
timestamp 1698431365
transform 1 0 13440 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_135
timestamp 1698431365
transform 1 0 16464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_137
timestamp 1698431365
transform 1 0 16688 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_225
timestamp 1698431365
transform 1 0 26544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698431365
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_295
timestamp 1698431365
transform 1 0 34384 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_330
timestamp 1698431365
transform 1 0 38304 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_334
timestamp 1698431365
transform 1 0 38752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698431365
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_356
timestamp 1698431365
transform 1 0 41216 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_389
timestamp 1698431365
transform 1 0 44912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_391
timestamp 1698431365
transform 1 0 45136 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_410
timestamp 1698431365
transform 1 0 47264 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_25
timestamp 1698431365
transform 1 0 4144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_57
timestamp 1698431365
transform 1 0 7728 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_59
timestamp 1698431365
transform 1 0 7952 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_75
timestamp 1698431365
transform 1 0 9744 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_155
timestamp 1698431365
transform 1 0 18704 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_157
timestamp 1698431365
transform 1 0 18928 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_232
timestamp 1698431365
transform 1 0 27328 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698431365
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_291
timestamp 1698431365
transform 1 0 33936 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_300
timestamp 1698431365
transform 1 0 34944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_310
timestamp 1698431365
transform 1 0 36064 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_312
timestamp 1698431365
transform 1 0 36288 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_325
timestamp 1698431365
transform 1 0 37744 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_327
timestamp 1698431365
transform 1 0 37968 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_359
timestamp 1698431365
transform 1 0 41552 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_365
timestamp 1698431365
transform 1 0 42224 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_383
timestamp 1698431365
transform 1 0 44240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_387
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_12
timestamp 1698431365
transform 1 0 2688 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_28
timestamp 1698431365
transform 1 0 4480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_68
timestamp 1698431365
transform 1 0 8960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_84
timestamp 1698431365
transform 1 0 10752 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_192
timestamp 1698431365
transform 1 0 22848 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_232
timestamp 1698431365
transform 1 0 27328 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_250
timestamp 1698431365
transform 1 0 29344 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_274
timestamp 1698431365
transform 1 0 32032 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_278
timestamp 1698431365
transform 1 0 32480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_373
timestamp 1698431365
transform 1 0 43120 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_403
timestamp 1698431365
transform 1 0 46480 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_412
timestamp 1698431365
transform 1 0 47488 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_416
timestamp 1698431365
transform 1 0 47936 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_20
timestamp 1698431365
transform 1 0 3584 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_69
timestamp 1698431365
transform 1 0 9072 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_91
timestamp 1698431365
transform 1 0 11536 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_163
timestamp 1698431365
transform 1 0 19600 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_185
timestamp 1698431365
transform 1 0 22064 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_211
timestamp 1698431365
transform 1 0 24976 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_225
timestamp 1698431365
transform 1 0 26544 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_227
timestamp 1698431365
transform 1 0 26768 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_240
timestamp 1698431365
transform 1 0 28224 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_242
timestamp 1698431365
transform 1 0 28448 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_251
timestamp 1698431365
transform 1 0 29456 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_257
timestamp 1698431365
transform 1 0 30128 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_290
timestamp 1698431365
transform 1 0 33824 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_294
timestamp 1698431365
transform 1 0 34272 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_296
timestamp 1698431365
transform 1 0 34496 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_305
timestamp 1698431365
transform 1 0 35504 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_309
timestamp 1698431365
transform 1 0 35952 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_382
timestamp 1698431365
transform 1 0 44128 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_384
timestamp 1698431365
transform 1 0 44352 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_415
timestamp 1698431365
transform 1 0 47824 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_419
timestamp 1698431365
transform 1 0 48272 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_37
timestamp 1698431365
transform 1 0 5488 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_39
timestamp 1698431365
transform 1 0 5712 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_69
timestamp 1698431365
transform 1 0 9072 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_127
timestamp 1698431365
transform 1 0 15568 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_139
timestamp 1698431365
transform 1 0 16912 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_193
timestamp 1698431365
transform 1 0 22960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_222
timestamp 1698431365
transform 1 0 26208 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_235
timestamp 1698431365
transform 1 0 27664 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_245
timestamp 1698431365
transform 1 0 28784 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_249
timestamp 1698431365
transform 1 0 29232 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_349
timestamp 1698431365
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_405
timestamp 1698431365
transform 1 0 46704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_409
timestamp 1698431365
transform 1 0 47152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_413
timestamp 1698431365
transform 1 0 47600 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_417
timestamp 1698431365
transform 1 0 48048 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_28
timestamp 1698431365
transform 1 0 4480 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_60
timestamp 1698431365
transform 1 0 8064 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_87
timestamp 1698431365
transform 1 0 11088 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_102
timestamp 1698431365
transform 1 0 12768 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_104
timestamp 1698431365
transform 1 0 12992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_120
timestamp 1698431365
transform 1 0 14784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_122
timestamp 1698431365
transform 1 0 15008 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_192
timestamp 1698431365
transform 1 0 22848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_211
timestamp 1698431365
transform 1 0 24976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_213
timestamp 1698431365
transform 1 0 25200 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_219
timestamp 1698431365
transform 1 0 25872 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_319
timestamp 1698431365
transform 1 0 37072 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_334
timestamp 1698431365
transform 1 0 38752 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_367
timestamp 1698431365
transform 1 0 42448 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_371
timestamp 1698431365
transform 1 0 42896 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_383
timestamp 1698431365
transform 1 0 44240 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_393
timestamp 1698431365
transform 1 0 45360 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_411
timestamp 1698431365
transform 1 0 47376 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_25
timestamp 1698431365
transform 1 0 4144 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_144
timestamp 1698431365
transform 1 0 17472 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_177
timestamp 1698431365
transform 1 0 21168 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_225
timestamp 1698431365
transform 1 0 26544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_227
timestamp 1698431365
transform 1 0 26768 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_234
timestamp 1698431365
transform 1 0 27552 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_238
timestamp 1698431365
transform 1 0 28000 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_240
timestamp 1698431365
transform 1 0 28224 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_254
timestamp 1698431365
transform 1 0 29792 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_272
timestamp 1698431365
transform 1 0 31808 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_276
timestamp 1698431365
transform 1 0 32256 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_305
timestamp 1698431365
transform 1 0 35504 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_315
timestamp 1698431365
transform 1 0 36624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_317
timestamp 1698431365
transform 1 0 36848 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_344
timestamp 1698431365
transform 1 0 39872 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_348
timestamp 1698431365
transform 1 0 40320 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_360
timestamp 1698431365
transform 1 0 41664 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_390
timestamp 1698431365
transform 1 0 45024 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_12
timestamp 1698431365
transform 1 0 2688 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_49
timestamp 1698431365
transform 1 0 6832 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_56
timestamp 1698431365
transform 1 0 7616 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_87
timestamp 1698431365
transform 1 0 11088 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_97
timestamp 1698431365
transform 1 0 12208 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_123
timestamp 1698431365
transform 1 0 15120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_166
timestamp 1698431365
transform 1 0 19936 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_168
timestamp 1698431365
transform 1 0 20160 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_225
timestamp 1698431365
transform 1 0 26544 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_242
timestamp 1698431365
transform 1 0 28448 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_244
timestamp 1698431365
transform 1 0 28672 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_255
timestamp 1698431365
transform 1 0 29904 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_301
timestamp 1698431365
transform 1 0 35056 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_305
timestamp 1698431365
transform 1 0 35504 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_312
timestamp 1698431365
transform 1 0 36288 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_314
timestamp 1698431365
transform 1 0 36512 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_336
timestamp 1698431365
transform 1 0 38976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_367
timestamp 1698431365
transform 1 0 42448 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_371
timestamp 1698431365
transform 1 0 42896 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_382
timestamp 1698431365
transform 1 0 44128 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_384
timestamp 1698431365
transform 1 0 44352 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_391
timestamp 1698431365
transform 1 0 45136 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_395
timestamp 1698431365
transform 1 0 45584 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_418
timestamp 1698431365
transform 1 0 48160 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_43
timestamp 1698431365
transform 1 0 6160 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_54
timestamp 1698431365
transform 1 0 7392 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_69
timestamp 1698431365
transform 1 0 9072 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_95
timestamp 1698431365
transform 1 0 11984 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_97
timestamp 1698431365
transform 1 0 12208 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_130
timestamp 1698431365
transform 1 0 15904 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_139
timestamp 1698431365
transform 1 0 16912 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_166
timestamp 1698431365
transform 1 0 19936 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_196
timestamp 1698431365
transform 1 0 23296 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_220
timestamp 1698431365
transform 1 0 25984 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_277
timestamp 1698431365
transform 1 0 32368 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_279
timestamp 1698431365
transform 1 0 32592 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_290
timestamp 1698431365
transform 1 0 33824 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_349
timestamp 1698431365
transform 1 0 40432 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_356
timestamp 1698431365
transform 1 0 41216 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_360
timestamp 1698431365
transform 1 0 41664 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_393
timestamp 1698431365
transform 1 0 45360 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_413
timestamp 1698431365
transform 1 0 47600 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_417
timestamp 1698431365
transform 1 0 48048 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_419
timestamp 1698431365
transform 1 0 48272 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_6
timestamp 1698431365
transform 1 0 2016 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_18
timestamp 1698431365
transform 1 0 3360 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_20
timestamp 1698431365
transform 1 0 3584 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_23
timestamp 1698431365
transform 1 0 3920 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_27
timestamp 1698431365
transform 1 0 4368 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_31
timestamp 1698431365
transform 1 0 4816 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_50
timestamp 1698431365
transform 1 0 6944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_63
timestamp 1698431365
transform 1 0 8400 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_82
timestamp 1698431365
transform 1 0 10528 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_102
timestamp 1698431365
transform 1 0 12768 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_104
timestamp 1698431365
transform 1 0 12992 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_117
timestamp 1698431365
transform 1 0 14448 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_140
timestamp 1698431365
transform 1 0 17024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_158
timestamp 1698431365
transform 1 0 19040 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_195
timestamp 1698431365
transform 1 0 23184 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_226
timestamp 1698431365
transform 1 0 26656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_255
timestamp 1698431365
transform 1 0 29904 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_257
timestamp 1698431365
transform 1 0 30128 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_273
timestamp 1698431365
transform 1 0 31920 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_275
timestamp 1698431365
transform 1 0 32144 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_284
timestamp 1698431365
transform 1 0 33152 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_288
timestamp 1698431365
transform 1 0 33600 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_292
timestamp 1698431365
transform 1 0 34048 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_297
timestamp 1698431365
transform 1 0 34608 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_314
timestamp 1698431365
transform 1 0 36512 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_323
timestamp 1698431365
transform 1 0 37520 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_363
timestamp 1698431365
transform 1 0 42000 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_365
timestamp 1698431365
transform 1 0 42224 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_376
timestamp 1698431365
transform 1 0 43456 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_378
timestamp 1698431365
transform 1 0 43680 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_387
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_31
timestamp 1698431365
transform 1 0 4816 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_37
timestamp 1698431365
transform 1 0 5488 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_61
timestamp 1698431365
transform 1 0 8176 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_69
timestamp 1698431365
transform 1 0 9072 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_118
timestamp 1698431365
transform 1 0 14560 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_120
timestamp 1698431365
transform 1 0 14784 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_133
timestamp 1698431365
transform 1 0 16240 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_183
timestamp 1698431365
transform 1 0 21840 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_185
timestamp 1698431365
transform 1 0 22064 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_204
timestamp 1698431365
transform 1 0 24192 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_208
timestamp 1698431365
transform 1 0 24640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_216
timestamp 1698431365
transform 1 0 25536 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_220
timestamp 1698431365
transform 1 0 25984 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_250
timestamp 1698431365
transform 1 0 29344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_252
timestamp 1698431365
transform 1 0 29568 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_278
timestamp 1698431365
transform 1 0 32480 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_342
timestamp 1698431365
transform 1 0 39648 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698431365
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_354
timestamp 1698431365
transform 1 0 40992 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_371
timestamp 1698431365
transform 1 0 42896 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_375
timestamp 1698431365
transform 1 0 43344 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_384
timestamp 1698431365
transform 1 0 44352 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_390
timestamp 1698431365
transform 1 0 45024 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_6
timestamp 1698431365
transform 1 0 2016 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_10
timestamp 1698431365
transform 1 0 2464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_14
timestamp 1698431365
transform 1 0 2912 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_59
timestamp 1698431365
transform 1 0 7952 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_68
timestamp 1698431365
transform 1 0 8960 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_102
timestamp 1698431365
transform 1 0 12768 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_104
timestamp 1698431365
transform 1 0 12992 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_174
timestamp 1698431365
transform 1 0 20832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_206
timestamp 1698431365
transform 1 0 24416 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_210
timestamp 1698431365
transform 1 0 24864 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_214
timestamp 1698431365
transform 1 0 25312 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_218
timestamp 1698431365
transform 1 0 25760 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_239
timestamp 1698431365
transform 1 0 28112 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_255
timestamp 1698431365
transform 1 0 29904 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_257
timestamp 1698431365
transform 1 0 30128 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_304
timestamp 1698431365
transform 1 0 35392 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_330
timestamp 1698431365
transform 1 0 38304 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_344
timestamp 1698431365
transform 1 0 39872 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_348
timestamp 1698431365
transform 1 0 40320 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_350
timestamp 1698431365
transform 1 0 40544 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_371
timestamp 1698431365
transform 1 0 42896 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_402
timestamp 1698431365
transform 1 0 46368 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_419
timestamp 1698431365
transform 1 0 48272 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_52
timestamp 1698431365
transform 1 0 7168 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_137
timestamp 1698431365
transform 1 0 16688 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_139
timestamp 1698431365
transform 1 0 16912 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_146
timestamp 1698431365
transform 1 0 17696 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_150
timestamp 1698431365
transform 1 0 18144 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_153
timestamp 1698431365
transform 1 0 18480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_185
timestamp 1698431365
transform 1 0 22064 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_189
timestamp 1698431365
transform 1 0 22512 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_202
timestamp 1698431365
transform 1 0 23968 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_220
timestamp 1698431365
transform 1 0 25984 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_222
timestamp 1698431365
transform 1 0 26208 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_225
timestamp 1698431365
transform 1 0 26544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_258
timestamp 1698431365
transform 1 0 30240 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_260
timestamp 1698431365
transform 1 0 30464 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_276
timestamp 1698431365
transform 1 0 32256 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_286
timestamp 1698431365
transform 1 0 33376 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_289
timestamp 1698431365
transform 1 0 33712 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_313
timestamp 1698431365
transform 1 0 36400 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_315
timestamp 1698431365
transform 1 0 36624 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_387
timestamp 1698431365
transform 1 0 44688 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_417
timestamp 1698431365
transform 1 0 48048 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_419
timestamp 1698431365
transform 1 0 48272 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_6
timestamp 1698431365
transform 1 0 2016 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_9
timestamp 1698431365
transform 1 0 2352 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_13
timestamp 1698431365
transform 1 0 2800 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_15
timestamp 1698431365
transform 1 0 3024 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_31
timestamp 1698431365
transform 1 0 4816 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_41
timestamp 1698431365
transform 1 0 5936 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_43
timestamp 1698431365
transform 1 0 6160 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_52
timestamp 1698431365
transform 1 0 7168 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_58
timestamp 1698431365
transform 1 0 7840 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_76
timestamp 1698431365
transform 1 0 9856 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_78
timestamp 1698431365
transform 1 0 10080 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_89
timestamp 1698431365
transform 1 0 11312 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_101
timestamp 1698431365
transform 1 0 12656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_140
timestamp 1698431365
transform 1 0 17024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_171
timestamp 1698431365
transform 1 0 20496 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_183
timestamp 1698431365
transform 1 0 21840 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_185
timestamp 1698431365
transform 1 0 22064 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_210
timestamp 1698431365
transform 1 0 24864 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_212
timestamp 1698431365
transform 1 0 25088 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_244
timestamp 1698431365
transform 1 0 28672 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_271
timestamp 1698431365
transform 1 0 31696 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_301
timestamp 1698431365
transform 1 0 35056 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_327
timestamp 1698431365
transform 1 0 37968 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_331
timestamp 1698431365
transform 1 0 38416 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_335
timestamp 1698431365
transform 1 0 38864 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_339
timestamp 1698431365
transform 1 0 39312 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_343
timestamp 1698431365
transform 1 0 39760 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698431365
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_383
timestamp 1698431365
transform 1 0 44240 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_410
timestamp 1698431365
transform 1 0 47264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_6
timestamp 1698431365
transform 1 0 2016 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_8
timestamp 1698431365
transform 1 0 2240 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_34
timestamp 1698431365
transform 1 0 5152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_64
timestamp 1698431365
transform 1 0 8512 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_68
timestamp 1698431365
transform 1 0 8960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_77
timestamp 1698431365
transform 1 0 9968 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_79
timestamp 1698431365
transform 1 0 10192 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_90
timestamp 1698431365
transform 1 0 11424 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_94
timestamp 1698431365
transform 1 0 11872 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_97
timestamp 1698431365
transform 1 0 12208 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_119
timestamp 1698431365
transform 1 0 14672 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_139
timestamp 1698431365
transform 1 0 16912 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_150
timestamp 1698431365
transform 1 0 18144 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_154
timestamp 1698431365
transform 1 0 18592 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_158
timestamp 1698431365
transform 1 0 19040 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_162
timestamp 1698431365
transform 1 0 19488 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_209
timestamp 1698431365
transform 1 0 24752 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_238
timestamp 1698431365
transform 1 0 28000 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_242
timestamp 1698431365
transform 1 0 28448 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_269
timestamp 1698431365
transform 1 0 31472 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_273
timestamp 1698431365
transform 1 0 31920 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_276
timestamp 1698431365
transform 1 0 32256 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_294
timestamp 1698431365
transform 1 0 34272 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_296
timestamp 1698431365
transform 1 0 34496 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_305
timestamp 1698431365
transform 1 0 35504 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_312
timestamp 1698431365
transform 1 0 36288 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_348
timestamp 1698431365
transform 1 0 40320 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_356
timestamp 1698431365
transform 1 0 41216 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_369
timestamp 1698431365
transform 1 0 42672 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_390
timestamp 1698431365
transform 1 0 45024 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_31
timestamp 1698431365
transform 1 0 4816 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_72
timestamp 1698431365
transform 1 0 9408 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_82
timestamp 1698431365
transform 1 0 10528 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_96
timestamp 1698431365
transform 1 0 12096 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_164
timestamp 1698431365
transform 1 0 19712 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_168
timestamp 1698431365
transform 1 0 20160 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_189
timestamp 1698431365
transform 1 0 22512 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_214
timestamp 1698431365
transform 1 0 25312 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_216
timestamp 1698431365
transform 1 0 25536 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_229
timestamp 1698431365
transform 1 0 26992 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_231
timestamp 1698431365
transform 1 0 27216 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_234
timestamp 1698431365
transform 1 0 27552 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_242
timestamp 1698431365
transform 1 0 28448 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_244
timestamp 1698431365
transform 1 0 28672 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_259
timestamp 1698431365
transform 1 0 30352 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_292
timestamp 1698431365
transform 1 0 34048 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_294
timestamp 1698431365
transform 1 0 34272 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_297
timestamp 1698431365
transform 1 0 34608 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_303
timestamp 1698431365
transform 1 0 35280 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_307
timestamp 1698431365
transform 1 0 35728 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_327
timestamp 1698431365
transform 1 0 37968 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_6
timestamp 1698431365
transform 1 0 2016 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_31
timestamp 1698431365
transform 1 0 4816 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_35
timestamp 1698431365
transform 1 0 5264 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_43
timestamp 1698431365
transform 1 0 6160 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_47
timestamp 1698431365
transform 1 0 6608 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_61
timestamp 1698431365
transform 1 0 8176 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_63
timestamp 1698431365
transform 1 0 8400 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_66
timestamp 1698431365
transform 1 0 8736 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_98
timestamp 1698431365
transform 1 0 12320 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_102
timestamp 1698431365
transform 1 0 12768 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_106
timestamp 1698431365
transform 1 0 13216 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_111
timestamp 1698431365
transform 1 0 13776 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_115
timestamp 1698431365
transform 1 0 14224 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_118
timestamp 1698431365
transform 1 0 14560 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_122
timestamp 1698431365
transform 1 0 15008 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_125
timestamp 1698431365
transform 1 0 15344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_129
timestamp 1698431365
transform 1 0 15792 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_131
timestamp 1698431365
transform 1 0 16016 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_134
timestamp 1698431365
transform 1 0 16352 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_208
timestamp 1698431365
transform 1 0 24640 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_227
timestamp 1698431365
transform 1 0 26768 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_328
timestamp 1698431365
transform 1 0 38080 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_418
timestamp 1698431365
transform 1 0 48160 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_32
timestamp 1698431365
transform 1 0 4928 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_41
timestamp 1698431365
transform 1 0 5936 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_45
timestamp 1698431365
transform 1 0 6384 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_69
timestamp 1698431365
transform 1 0 9072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_73
timestamp 1698431365
transform 1 0 9520 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_80
timestamp 1698431365
transform 1 0 10304 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_94
timestamp 1698431365
transform 1 0 11872 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_104
timestamp 1698431365
transform 1 0 12992 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_116
timestamp 1698431365
transform 1 0 14336 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_120
timestamp 1698431365
transform 1 0 14784 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_124
timestamp 1698431365
transform 1 0 15232 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_133
timestamp 1698431365
transform 1 0 16240 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_149
timestamp 1698431365
transform 1 0 18032 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_152
timestamp 1698431365
transform 1 0 18368 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_156
timestamp 1698431365
transform 1 0 18816 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_163
timestamp 1698431365
transform 1 0 19600 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_173
timestamp 1698431365
transform 1 0 20720 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_185
timestamp 1698431365
transform 1 0 22064 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_189
timestamp 1698431365
transform 1 0 22512 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_191
timestamp 1698431365
transform 1 0 22736 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_194
timestamp 1698431365
transform 1 0 23072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_198
timestamp 1698431365
transform 1 0 23520 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_213
timestamp 1698431365
transform 1 0 25200 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_217
timestamp 1698431365
transform 1 0 25648 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_240
timestamp 1698431365
transform 1 0 28224 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_242
timestamp 1698431365
transform 1 0 28448 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_251
timestamp 1698431365
transform 1 0 29456 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_262
timestamp 1698431365
transform 1 0 30688 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_264
timestamp 1698431365
transform 1 0 30912 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_276
timestamp 1698431365
transform 1 0 32256 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_319
timestamp 1698431365
transform 1 0 37072 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_335
timestamp 1698431365
transform 1 0 38864 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_60
timestamp 1698431365
transform 1 0 8064 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_64
timestamp 1698431365
transform 1 0 8512 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_68
timestamp 1698431365
transform 1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_87
timestamp 1698431365
transform 1 0 11088 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_89
timestamp 1698431365
transform 1 0 11312 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_146
timestamp 1698431365
transform 1 0 17696 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_217
timestamp 1698431365
transform 1 0 25648 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_219
timestamp 1698431365
transform 1 0 25872 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_254
timestamp 1698431365
transform 1 0 29792 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_290
timestamp 1698431365
transform 1 0 33824 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_331
timestamp 1698431365
transform 1 0 38416 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_10
timestamp 1698431365
transform 1 0 2464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_33
timestamp 1698431365
transform 1 0 5040 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_47
timestamp 1698431365
transform 1 0 6608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_60
timestamp 1698431365
transform 1 0 8064 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_62
timestamp 1698431365
transform 1 0 8288 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_69
timestamp 1698431365
transform 1 0 9072 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_136
timestamp 1698431365
transform 1 0 16576 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_138
timestamp 1698431365
transform 1 0 16800 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_141
timestamp 1698431365
transform 1 0 17136 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_173
timestamp 1698431365
transform 1 0 20720 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_201
timestamp 1698431365
transform 1 0 23856 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_203
timestamp 1698431365
transform 1 0 24080 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_209
timestamp 1698431365
transform 1 0 24752 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_211
timestamp 1698431365
transform 1 0 24976 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_216
timestamp 1698431365
transform 1 0 25536 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_233
timestamp 1698431365
transform 1 0 27440 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_242
timestamp 1698431365
transform 1 0 28448 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_244
timestamp 1698431365
transform 1 0 28672 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_313
timestamp 1698431365
transform 1 0 36400 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_334
timestamp 1698431365
transform 1 0 38752 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_370
timestamp 1698431365
transform 1 0 42784 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_413
timestamp 1698431365
transform 1 0 47600 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_6
timestamp 1698431365
transform 1 0 2016 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_14
timestamp 1698431365
transform 1 0 2912 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_24
timestamp 1698431365
transform 1 0 4032 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_50
timestamp 1698431365
transform 1 0 6944 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_68
timestamp 1698431365
transform 1 0 8960 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_82
timestamp 1698431365
transform 1 0 10528 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_86
timestamp 1698431365
transform 1 0 10976 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_90
timestamp 1698431365
transform 1 0 11424 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_94
timestamp 1698431365
transform 1 0 11872 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_116
timestamp 1698431365
transform 1 0 14336 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_139
timestamp 1698431365
transform 1 0 16912 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_171
timestamp 1698431365
transform 1 0 20496 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_179
timestamp 1698431365
transform 1 0 21392 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_185
timestamp 1698431365
transform 1 0 22064 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_194
timestamp 1698431365
transform 1 0 23072 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_196
timestamp 1698431365
transform 1 0 23296 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_209
timestamp 1698431365
transform 1 0 24752 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_219
timestamp 1698431365
transform 1 0 25872 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_231
timestamp 1698431365
transform 1 0 27216 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_295
timestamp 1698431365
transform 1 0 34384 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_342
timestamp 1698431365
transform 1 0 39648 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_32
timestamp 1698431365
transform 1 0 4928 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_46
timestamp 1698431365
transform 1 0 6496 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_109
timestamp 1698431365
transform 1 0 13552 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_165
timestamp 1698431365
transform 1 0 19824 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_169
timestamp 1698431365
transform 1 0 20272 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_173
timestamp 1698431365
transform 1 0 20720 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_181
timestamp 1698431365
transform 1 0 21616 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_185
timestamp 1698431365
transform 1 0 22064 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_189
timestamp 1698431365
transform 1 0 22512 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_191
timestamp 1698431365
transform 1 0 22736 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_222
timestamp 1698431365
transform 1 0 26208 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_243
timestamp 1698431365
transform 1 0 28560 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_249
timestamp 1698431365
transform 1 0 29232 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_305
timestamp 1698431365
transform 1 0 35504 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_355
timestamp 1698431365
transform 1 0 41104 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_419
timestamp 1698431365
transform 1 0 48272 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_10
timestamp 1698431365
transform 1 0 2464 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_12
timestamp 1698431365
transform 1 0 2688 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_21
timestamp 1698431365
transform 1 0 3696 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_29
timestamp 1698431365
transform 1 0 4592 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_65
timestamp 1698431365
transform 1 0 8624 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_67
timestamp 1698431365
transform 1 0 8848 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_109
timestamp 1698431365
transform 1 0 13552 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_142
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_209
timestamp 1698431365
transform 1 0 24752 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_212
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_218
timestamp 1698431365
transform 1 0 25760 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_258
timestamp 1698431365
transform 1 0 30240 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_262
timestamp 1698431365
transform 1 0 30688 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_266
timestamp 1698431365
transform 1 0 31136 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_270
timestamp 1698431365
transform 1 0 31584 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_349
timestamp 1698431365
transform 1 0 40432 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_18
timestamp 1698431365
transform 1 0 3360 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_20
timestamp 1698431365
transform 1 0 3584 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_25
timestamp 1698431365
transform 1 0 4144 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_33
timestamp 1698431365
transform 1 0 5040 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_40
timestamp 1698431365
transform 1 0 5824 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_48
timestamp 1698431365
transform 1 0 6720 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_53
timestamp 1698431365
transform 1 0 7280 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_57
timestamp 1698431365
transform 1 0 7728 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_61
timestamp 1698431365
transform 1 0 8176 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_67
timestamp 1698431365
transform 1 0 8848 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_76
timestamp 1698431365
transform 1 0 9856 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_81
timestamp 1698431365
transform 1 0 10416 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_87
timestamp 1698431365
transform 1 0 11088 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_95
timestamp 1698431365
transform 1 0 11984 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_97
timestamp 1698431365
transform 1 0 12208 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_133
timestamp 1698431365
transform 1 0 16240 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_135
timestamp 1698431365
transform 1 0 16464 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_142
timestamp 1698431365
transform 1 0 17248 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_172
timestamp 1698431365
transform 1 0 20608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_174
timestamp 1698431365
transform 1 0 20832 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_201
timestamp 1698431365
transform 1 0 23856 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_203
timestamp 1698431365
transform 1 0 24080 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_236
timestamp 1698431365
transform 1 0 27776 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_240
timestamp 1698431365
transform 1 0 28224 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_303
timestamp 1698431365
transform 1 0 35280 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_305
timestamp 1698431365
transform 1 0 35504 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_418
timestamp 1698431365
transform 1 0 48160 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input1
timestamp 1698431365
transform 1 0 44800 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 48384 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input3
timestamp 1698431365
transform -1 0 48384 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform -1 0 48384 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input5
timestamp 1698431365
transform -1 0 48384 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform -1 0 48384 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform -1 0 48384 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform -1 0 48384 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input9
timestamp 1698431365
transform -1 0 48384 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input10
timestamp 1698431365
transform -1 0 48384 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input11
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input12
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698431365
transform -1 0 20384 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698431365
transform -1 0 27328 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698431365
transform -1 0 31808 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698431365
transform 1 0 32592 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698431365
transform 1 0 35840 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698431365
transform -1 0 37968 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698431365
transform -1 0 39760 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698431365
transform -1 0 42560 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698431365
transform -1 0 43680 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698431365
transform 1 0 43456 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698431365
transform 1 0 45472 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output27
timestamp 1698431365
transform -1 0 16576 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output28
timestamp 1698431365
transform 1 0 17808 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_55 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 48608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 48608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 48608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 48608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 48608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 48608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 48608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 48608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 48608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 48608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 48608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 48608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 48608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 48608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 48608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 48608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 48608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 48608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 48608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 48608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 48608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 48608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 48608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_78
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 48608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_79
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 48608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_80
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 48608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_81
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 48608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 48608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 48608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 48608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 48608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_86
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 48608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_87
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 48608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_88
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 48608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_89
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 48608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_90
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 48608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_91
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 48608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_92
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 48608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_93
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 48608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_94
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 48608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_95
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 48608 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_96
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 48608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_97
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 48608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_98
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 48608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_99
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 48608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_100
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 48608 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_101
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 48608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_102
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 48608 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_103
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 48608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_104
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 48608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_105
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 48608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_106
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 48608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_107
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 48608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_108
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 48608 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_109
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 48608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer1
timestamp 1698431365
transform 1 0 16352 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer2
timestamp 1698431365
transform -1 0 48272 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer3
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  rebuffer4
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer5
timestamp 1698431365
transform 1 0 11424 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer6
timestamp 1698431365
transform 1 0 11536 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer7
timestamp 1698431365
transform 1 0 33152 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer8
timestamp 1698431365
transform -1 0 10752 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer9
timestamp 1698431365
transform -1 0 27552 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer10
timestamp 1698431365
transform -1 0 17024 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer11
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer12
timestamp 1698431365
transform -1 0 16240 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer13
timestamp 1698431365
transform 1 0 31808 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  rebuffer14
timestamp 1698431365
transform 1 0 35168 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer15
timestamp 1698431365
transform -1 0 32704 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dlya_2  rebuffer16 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  rebuffer17
timestamp 1698431365
transform 1 0 32256 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer18
timestamp 1698431365
transform -1 0 16912 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  rebuffer19
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  rebuffer20
timestamp 1698431365
transform 1 0 14896 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  rebuffer21
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_110 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_111
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_112
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_113
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_114
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_115
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_116
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_117
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_118
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_119
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_120
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_121
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_122
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_123
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_124
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_125
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_126
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_127
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_128
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_129
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_130
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_131
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_132
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_133
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_134
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_135
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_136
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_137
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_138
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_139
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_140
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_141
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_142
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_143
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_144
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_145
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_146
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_147
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_148
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_149
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_150
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_151
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_152
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_153
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_154
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_155
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_156
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_157
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_158
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_159
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_160
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_161
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_162
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_163
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_164
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_165
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_166
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_167
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_168
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_169
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_170
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_171
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_172
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_173
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_174
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_175
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_176
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_177
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_178
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_179
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_180
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_181
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_182
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_183
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_184
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_185
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_186
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_187
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_188
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_189
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_190
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_191
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_192
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_193
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_194
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_195
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_196
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_197
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_198
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_199
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_200
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_201
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_202
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_203
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_204
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_205
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_206
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_207
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_208
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_209
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_210
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_211
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_212
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_213
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_214
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_215
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_216
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_217
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_218
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_219
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_220
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_221
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_222
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_223
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_224
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_225
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_226
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_227
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_228
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_229
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_230
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_231
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_232
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_233
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_234
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_235
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_236
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_237
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_238
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_239
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_240
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_241
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_242
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_243
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_244
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_245
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_246
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_247
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_248
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_249
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_250
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_251
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_252
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_253
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_254
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_255
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_256
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_257
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_258
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_259
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_260
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_261
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_262
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_263
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_264
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_265
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_266
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_267
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_268
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_269
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_270
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_271
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_272
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_273
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_274
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_275
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_276
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_277
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_278
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_279
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_280
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_281
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_282
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_283
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_284
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_285
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_286
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_287
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_288
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_289
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_290
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_291
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_292
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_293
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_294
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_295
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_296
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_297
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_298
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_299
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_300
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_301
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_302
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_303
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_304
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_305
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_306
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_307
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_308
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_309
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_310
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_311
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_312
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_313
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_314
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_315
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_316
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_317
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_318
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_319
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_320
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_321
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_322
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_323
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_324
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_325
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_326
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_327
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_328
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_329
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_330
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_331
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_332
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_333
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_334
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_335
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_336
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_337
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_338
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_339
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_340
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_341
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_342
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_343
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_344
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_345
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_346
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_347
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_348
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_349
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_350
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_351
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_352
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_353
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_354
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_355
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_356
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_357
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_358
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_359
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_360
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_361
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_362
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_363
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_364
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_365
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_366
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_367
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_368
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_369
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_370
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_371
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_372
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_373
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_374
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_375
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_376
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_377
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_378
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_379
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_380
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_381
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_382
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_383
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_384
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_385
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_386
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_387
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_388
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_389
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_390
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_391
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_392
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_393
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_394
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_395
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_396
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_397
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_398
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_399
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_400
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_401
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_402
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_403
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_404
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_405
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_406
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_407
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_408
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_409
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_410
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_411
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_412
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_413
timestamp 1698431365
transform 1 0 5152 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_414
timestamp 1698431365
transform 1 0 8960 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_415
timestamp 1698431365
transform 1 0 12768 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_416
timestamp 1698431365
transform 1 0 16576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_417
timestamp 1698431365
transform 1 0 20384 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_418
timestamp 1698431365
transform 1 0 24192 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_419
timestamp 1698431365
transform 1 0 28000 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_420
timestamp 1698431365
transform 1 0 31808 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_421
timestamp 1698431365
transform 1 0 35616 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_422
timestamp 1698431365
transform 1 0 39424 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_423
timestamp 1698431365
transform 1 0 43232 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_424
timestamp 1698431365
transform 1 0 47040 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_29 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4144 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_30
timestamp 1698431365
transform -1 0 5824 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_31
timestamp 1698431365
transform -1 0 7280 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_32
timestamp 1698431365
transform -1 0 8848 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_33
timestamp 1698431365
transform -1 0 10416 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_34
timestamp 1698431365
transform -1 0 11984 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_35
timestamp 1698431365
transform 1 0 12320 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_36
timestamp 1698431365
transform -1 0 17248 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_37
timestamp 1698431365
transform 1 0 23072 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_38
timestamp 1698431365
transform -1 0 26992 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_39
timestamp 1698431365
transform -1 0 27776 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_40
timestamp 1698431365
transform 1 0 28448 0 1 45472
box -86 -86 534 870
<< labels >>
flabel metal3 s 49200 42112 50000 42224 0 FreeSans 448 0 0 0 custom_settings[0]
port 0 nsew signal input
flabel metal3 s 49200 47040 50000 47152 0 FreeSans 448 0 0 0 custom_settings[1]
port 1 nsew signal input
flabel metal3 s 49200 2688 50000 2800 0 FreeSans 448 0 0 0 io_in_1[0]
port 2 nsew signal input
flabel metal3 s 49200 7616 50000 7728 0 FreeSans 448 0 0 0 io_in_1[1]
port 3 nsew signal input
flabel metal3 s 49200 12544 50000 12656 0 FreeSans 448 0 0 0 io_in_1[2]
port 4 nsew signal input
flabel metal3 s 49200 17472 50000 17584 0 FreeSans 448 0 0 0 io_in_1[3]
port 5 nsew signal input
flabel metal3 s 49200 22400 50000 22512 0 FreeSans 448 0 0 0 io_in_1[4]
port 6 nsew signal input
flabel metal3 s 49200 27328 50000 27440 0 FreeSans 448 0 0 0 io_in_1[5]
port 7 nsew signal input
flabel metal3 s 49200 32256 50000 32368 0 FreeSans 448 0 0 0 io_in_1[6]
port 8 nsew signal input
flabel metal3 s 49200 37184 50000 37296 0 FreeSans 448 0 0 0 io_in_1[7]
port 9 nsew signal input
flabel metal3 s 0 41440 800 41552 0 FreeSans 448 0 0 0 io_in_2
port 10 nsew signal input
flabel metal2 s 3584 49200 3696 50000 0 FreeSans 448 90 0 0 io_out[0]
port 11 nsew signal tristate
flabel metal2 s 19264 49200 19376 50000 0 FreeSans 448 90 0 0 io_out[10]
port 12 nsew signal tristate
flabel metal2 s 20832 49200 20944 50000 0 FreeSans 448 90 0 0 io_out[11]
port 13 nsew signal tristate
flabel metal2 s 22400 49200 22512 50000 0 FreeSans 448 90 0 0 io_out[12]
port 14 nsew signal tristate
flabel metal2 s 23968 49200 24080 50000 0 FreeSans 448 90 0 0 io_out[13]
port 15 nsew signal tristate
flabel metal2 s 25536 49200 25648 50000 0 FreeSans 448 90 0 0 io_out[14]
port 16 nsew signal tristate
flabel metal2 s 27104 49200 27216 50000 0 FreeSans 448 90 0 0 io_out[15]
port 17 nsew signal tristate
flabel metal2 s 28672 49200 28784 50000 0 FreeSans 448 90 0 0 io_out[16]
port 18 nsew signal tristate
flabel metal2 s 30240 49200 30352 50000 0 FreeSans 448 90 0 0 io_out[17]
port 19 nsew signal tristate
flabel metal2 s 31808 49200 31920 50000 0 FreeSans 448 90 0 0 io_out[18]
port 20 nsew signal tristate
flabel metal2 s 33376 49200 33488 50000 0 FreeSans 448 90 0 0 io_out[19]
port 21 nsew signal tristate
flabel metal2 s 5152 49200 5264 50000 0 FreeSans 448 90 0 0 io_out[1]
port 22 nsew signal tristate
flabel metal2 s 34944 49200 35056 50000 0 FreeSans 448 90 0 0 io_out[20]
port 23 nsew signal tristate
flabel metal2 s 36512 49200 36624 50000 0 FreeSans 448 90 0 0 io_out[21]
port 24 nsew signal tristate
flabel metal2 s 38080 49200 38192 50000 0 FreeSans 448 90 0 0 io_out[22]
port 25 nsew signal tristate
flabel metal2 s 39648 49200 39760 50000 0 FreeSans 448 90 0 0 io_out[23]
port 26 nsew signal tristate
flabel metal2 s 41216 49200 41328 50000 0 FreeSans 448 90 0 0 io_out[24]
port 27 nsew signal tristate
flabel metal2 s 42784 49200 42896 50000 0 FreeSans 448 90 0 0 io_out[25]
port 28 nsew signal tristate
flabel metal2 s 44352 49200 44464 50000 0 FreeSans 448 90 0 0 io_out[26]
port 29 nsew signal tristate
flabel metal2 s 45920 49200 46032 50000 0 FreeSans 448 90 0 0 io_out[27]
port 30 nsew signal tristate
flabel metal2 s 6720 49200 6832 50000 0 FreeSans 448 90 0 0 io_out[2]
port 31 nsew signal tristate
flabel metal2 s 8288 49200 8400 50000 0 FreeSans 448 90 0 0 io_out[3]
port 32 nsew signal tristate
flabel metal2 s 9856 49200 9968 50000 0 FreeSans 448 90 0 0 io_out[4]
port 33 nsew signal tristate
flabel metal2 s 11424 49200 11536 50000 0 FreeSans 448 90 0 0 io_out[5]
port 34 nsew signal tristate
flabel metal2 s 12992 49200 13104 50000 0 FreeSans 448 90 0 0 io_out[6]
port 35 nsew signal tristate
flabel metal2 s 14560 49200 14672 50000 0 FreeSans 448 90 0 0 io_out[7]
port 36 nsew signal tristate
flabel metal2 s 16128 49200 16240 50000 0 FreeSans 448 90 0 0 io_out[8]
port 37 nsew signal tristate
flabel metal2 s 17696 49200 17808 50000 0 FreeSans 448 90 0 0 io_out[9]
port 38 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 rst_n
port 39 nsew signal input
flabel metal4 s 4448 3076 4768 46316 0 FreeSans 1280 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 35168 3076 35488 46316 0 FreeSans 1280 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 19808 3076 20128 46316 0 FreeSans 1280 90 0 0 vss
port 41 nsew ground bidirectional
flabel metal3 s 0 8288 800 8400 0 FreeSans 448 0 0 0 wb_clk_i
port 42 nsew signal input
rlabel metal1 24976 46256 24976 46256 0 vdd
rlabel metal1 24976 45472 24976 45472 0 vss
rlabel metal2 43176 36736 43176 36736 0 _0000_
rlabel metal3 16240 8120 16240 8120 0 _0001_
rlabel metal2 16184 5264 16184 5264 0 _0002_
rlabel metal2 16072 4704 16072 4704 0 _0003_
rlabel metal2 16296 7000 16296 7000 0 _0004_
rlabel metal2 28840 7616 28840 7616 0 _0005_
rlabel metal2 27272 5488 27272 5488 0 _0006_
rlabel metal2 28168 5096 28168 5096 0 _0007_
rlabel metal3 25816 6664 25816 6664 0 _0008_
rlabel metal2 31584 11480 31584 11480 0 _0009_
rlabel metal2 29736 9464 29736 9464 0 _0010_
rlabel metal2 30856 9464 30856 9464 0 _0011_
rlabel metal2 31864 15148 31864 15148 0 _0012_
rlabel metal2 34328 27440 34328 27440 0 _0013_
rlabel metal2 35112 23128 35112 23128 0 _0014_
rlabel metal3 25424 28616 25424 28616 0 _0015_
rlabel metal2 21000 34608 21000 34608 0 _0016_
rlabel metal3 19824 31640 19824 31640 0 _0017_
rlabel metal2 18200 36008 18200 36008 0 _0018_
rlabel metal3 19880 37912 19880 37912 0 _0019_
rlabel metal2 21448 40040 21448 40040 0 _0020_
rlabel metal3 19544 43400 19544 43400 0 _0021_
rlabel metal2 15176 39088 15176 39088 0 _0022_
rlabel metal2 17752 40656 17752 40656 0 _0023_
rlabel metal2 9576 30184 9576 30184 0 _0024_
rlabel metal2 10136 33600 10136 33600 0 _0025_
rlabel metal2 17640 33992 17640 33992 0 _0026_
rlabel metal2 16408 37800 16408 37800 0 _0027_
rlabel metal2 11984 36232 11984 36232 0 _0028_
rlabel metal3 4256 37128 4256 37128 0 _0029_
rlabel metal2 2520 40152 2520 40152 0 _0030_
rlabel metal3 4256 41272 4256 41272 0 _0031_
rlabel metal2 2632 44464 2632 44464 0 _0032_
rlabel metal2 15960 41552 15960 41552 0 _0033_
rlabel metal2 14840 44352 14840 44352 0 _0034_
rlabel metal2 2464 25592 2464 25592 0 _0035_
rlabel metal2 3920 27944 3920 27944 0 _0036_
rlabel metal2 2520 31416 2520 31416 0 _0037_
rlabel metal2 8232 32704 8232 32704 0 _0038_
rlabel metal2 2520 34272 2520 34272 0 _0039_
rlabel metal2 2520 36008 2520 36008 0 _0040_
rlabel metal2 5992 39256 5992 39256 0 _0041_
rlabel metal2 5768 42000 5768 42000 0 _0042_
rlabel metal2 5656 45416 5656 45416 0 _0043_
rlabel metal2 10248 44688 10248 44688 0 _0044_
rlabel metal2 13048 45528 13048 45528 0 _0045_
rlabel metal2 42560 26152 42560 26152 0 _0046_
rlabel metal3 42504 27160 42504 27160 0 _0047_
rlabel metal2 46088 27384 46088 27384 0 _0048_
rlabel metal2 46088 24640 46088 24640 0 _0049_
rlabel metal2 43120 24136 43120 24136 0 _0050_
rlabel metal2 44072 21728 44072 21728 0 _0051_
rlabel metal3 43008 23016 43008 23016 0 _0052_
rlabel metal2 42392 18424 42392 18424 0 _0053_
rlabel metal2 43568 13944 43568 13944 0 _0054_
rlabel metal3 43568 6552 43568 6552 0 _0055_
rlabel metal2 46088 4648 46088 4648 0 _0056_
rlabel metal3 46536 5992 46536 5992 0 _0057_
rlabel metal2 46088 8400 46088 8400 0 _0058_
rlabel metal2 46088 9968 46088 9968 0 _0059_
rlabel metal3 44352 10696 44352 10696 0 _0060_
rlabel metal2 46088 12320 46088 12320 0 _0061_
rlabel metal2 46984 14168 46984 14168 0 _0062_
rlabel metal2 46088 16520 46088 16520 0 _0063_
rlabel metal2 46872 18928 46872 18928 0 _0064_
rlabel metal2 46144 18648 46144 18648 0 _0065_
rlabel metal2 44968 17192 44968 17192 0 _0066_
rlabel metal2 41776 16184 41776 16184 0 _0067_
rlabel metal3 42448 13048 42448 13048 0 _0068_
rlabel metal2 38472 13048 38472 13048 0 _0069_
rlabel metal2 39816 15960 39816 15960 0 _0070_
rlabel metal2 37800 19376 37800 19376 0 _0071_
rlabel metal3 36344 21448 36344 21448 0 _0072_
rlabel metal2 39256 22456 39256 22456 0 _0073_
rlabel metal2 41384 21112 41384 21112 0 _0074_
rlabel metal2 38024 24304 38024 24304 0 _0075_
rlabel metal2 37688 26684 37688 26684 0 _0076_
rlabel metal2 36792 28056 36792 28056 0 _0077_
rlabel metal2 34664 31416 34664 31416 0 _0078_
rlabel metal2 32760 33488 32760 33488 0 _0079_
rlabel metal2 27272 35280 27272 35280 0 _0080_
rlabel metal3 28784 37352 28784 37352 0 _0081_
rlabel metal2 27944 41552 27944 41552 0 _0082_
rlabel metal2 28112 42504 28112 42504 0 _0083_
rlabel metal3 24024 44968 24024 44968 0 _0084_
rlabel metal2 21336 44744 21336 44744 0 _0085_
rlabel metal2 42504 8456 42504 8456 0 _0086_
rlabel metal2 43736 4648 43736 4648 0 _0087_
rlabel metal2 41272 5152 41272 5152 0 _0088_
rlabel metal2 40040 5432 40040 5432 0 _0089_
rlabel metal2 41944 3864 41944 3864 0 _0090_
rlabel metal2 36792 4368 36792 4368 0 _0091_
rlabel metal2 38472 4648 38472 4648 0 _0092_
rlabel metal2 39032 12320 39032 12320 0 _0093_
rlabel metal2 35504 12712 35504 12712 0 _0094_
rlabel metal2 35336 15736 35336 15736 0 _0095_
rlabel metal2 33544 22008 33544 22008 0 _0096_
rlabel metal2 34440 8456 34440 8456 0 _0097_
rlabel metal2 35224 4648 35224 4648 0 _0098_
rlabel metal2 31304 4760 31304 4760 0 _0099_
rlabel metal2 25368 3864 25368 3864 0 _0100_
rlabel metal2 22120 3976 22120 3976 0 _0101_
rlabel metal2 19544 3976 19544 3976 0 _0102_
rlabel metal3 19264 8344 19264 8344 0 _0103_
rlabel metal2 23856 9912 23856 9912 0 _0104_
rlabel metal2 22624 12264 22624 12264 0 _0105_
rlabel metal2 23744 14728 23744 14728 0 _0106_
rlabel metal2 2688 17080 2688 17080 0 _0107_
rlabel metal3 13720 8904 13720 8904 0 _0108_
rlabel metal2 13160 3976 13160 3976 0 _0109_
rlabel metal2 10248 4816 10248 4816 0 _0110_
rlabel metal2 7560 3976 7560 3976 0 _0111_
rlabel metal2 5656 5544 5656 5544 0 _0112_
rlabel metal3 4928 7560 4928 7560 0 _0113_
rlabel metal2 4872 8680 4872 8680 0 _0114_
rlabel metal2 11928 10752 11928 10752 0 _0115_
rlabel metal2 12152 13328 12152 13328 0 _0116_
rlabel metal3 12040 15960 12040 15960 0 _0117_
rlabel metal2 10024 23688 10024 23688 0 _0118_
rlabel metal2 37464 29848 37464 29848 0 _0119_
rlabel metal2 39144 28280 39144 28280 0 _0120_
rlabel metal2 41440 31864 41440 31864 0 _0121_
rlabel metal2 37240 31136 37240 31136 0 _0122_
rlabel metal2 37352 35336 37352 35336 0 _0123_
rlabel metal2 34440 37688 34440 37688 0 _0124_
rlabel metal2 40152 39088 40152 39088 0 _0125_
rlabel metal2 36008 40824 36008 40824 0 _0126_
rlabel metal2 39368 43512 39368 43512 0 _0127_
rlabel metal2 37800 43456 37800 43456 0 _0128_
rlabel metal2 47376 41944 47376 41944 0 _0129_
rlabel metal2 43288 43120 43288 43120 0 _0130_
rlabel metal3 46144 45192 46144 45192 0 _0131_
rlabel metal3 42000 36232 42000 36232 0 _0132_
rlabel metal2 44184 29792 44184 29792 0 _0133_
rlabel metal2 46032 28728 46032 28728 0 _0134_
rlabel metal2 45864 34552 45864 34552 0 _0135_
rlabel metal2 46088 32872 46088 32872 0 _0136_
rlabel metal2 47096 40152 47096 40152 0 _0137_
rlabel metal2 44296 31808 44296 31808 0 _0138_
rlabel metal2 40152 33544 40152 33544 0 _0139_
rlabel metal2 38696 35056 38696 35056 0 _0140_
rlabel metal2 44408 34440 44408 34440 0 _0141_
rlabel metal2 38584 36848 38584 36848 0 _0142_
rlabel metal3 41384 37912 41384 37912 0 _0143_
rlabel metal2 47432 39312 47432 39312 0 _0144_
rlabel metal2 41720 41104 41720 41104 0 _0145_
rlabel metal3 41272 39032 41272 39032 0 _0146_
rlabel metal2 42280 39032 42280 39032 0 _0147_
rlabel metal2 46984 41384 46984 41384 0 _0148_
rlabel metal2 44856 36064 44856 36064 0 _0149_
rlabel metal2 47096 37632 47096 37632 0 _0150_
rlabel metal2 42504 20496 42504 20496 0 _0151_
rlabel metal2 29288 14896 29288 14896 0 _0152_
rlabel metal2 25704 9968 25704 9968 0 _0153_
rlabel metal2 28056 11536 28056 11536 0 _0154_
rlabel metal3 29064 13048 29064 13048 0 _0155_
rlabel metal3 25256 12992 25256 12992 0 _0156_
rlabel metal2 25928 15400 25928 15400 0 _0157_
rlabel metal2 15064 11256 15064 11256 0 _0158_
rlabel metal3 17584 9912 17584 9912 0 _0159_
rlabel metal2 18368 11368 18368 11368 0 _0160_
rlabel metal2 15176 12600 15176 12600 0 _0161_
rlabel metal2 18648 12992 18648 12992 0 _0162_
rlabel metal2 17752 14168 17752 14168 0 _0163_
rlabel metal2 4536 10920 4536 10920 0 _0164_
rlabel metal2 2968 11032 2968 11032 0 _0165_
rlabel metal2 4200 14056 4200 14056 0 _0166_
rlabel metal3 5040 12264 5040 12264 0 _0167_
rlabel metal2 7784 13496 7784 13496 0 _0168_
rlabel metal2 8456 16184 8456 16184 0 _0169_
rlabel metal3 25368 18312 25368 18312 0 _0170_
rlabel metal2 24640 19320 24640 19320 0 _0171_
rlabel metal2 22344 21840 22344 21840 0 _0172_
rlabel metal2 21336 19600 21336 19600 0 _0173_
rlabel metal2 16632 21952 16632 21952 0 _0174_
rlabel metal2 16744 22792 16744 22792 0 _0175_
rlabel metal2 19544 22792 19544 22792 0 _0176_
rlabel metal2 17864 20272 17864 20272 0 _0177_
rlabel metal3 4872 19320 4872 19320 0 _0178_
rlabel metal2 2744 19712 2744 19712 0 _0179_
rlabel metal2 3304 16688 3304 16688 0 _0180_
rlabel metal2 3864 18704 3864 18704 0 _0181_
rlabel metal3 8456 19096 8456 19096 0 _0182_
rlabel metal2 12992 19320 12992 19320 0 _0183_
rlabel metal2 12936 18424 12936 18424 0 _0184_
rlabel metal3 8400 17528 8400 17528 0 _0185_
rlabel metal3 13888 16744 13888 16744 0 _0186_
rlabel metal2 15176 15148 15176 15148 0 _0187_
rlabel metal3 13216 18424 13216 18424 0 _0188_
rlabel metal2 36176 17528 36176 17528 0 _0189_
rlabel metal2 30856 17304 30856 17304 0 _0190_
rlabel metal2 31528 18872 31528 18872 0 _0191_
rlabel metal2 34664 18032 34664 18032 0 _0192_
rlabel metal2 6440 37800 6440 37800 0 _0193_
rlabel metal2 40488 29176 40488 29176 0 _0194_
rlabel metal2 7336 40376 7336 40376 0 _0195_
rlabel metal3 7896 38808 7896 38808 0 _0196_
rlabel metal3 9296 41160 9296 41160 0 _0197_
rlabel metal2 8904 41944 8904 41944 0 _0198_
rlabel metal2 7952 42840 7952 42840 0 _0199_
rlabel metal2 9464 41888 9464 41888 0 _0200_
rlabel metal2 8680 43400 8680 43400 0 _0201_
rlabel metal2 9128 45080 9128 45080 0 _0202_
rlabel metal2 8232 44464 8232 44464 0 _0203_
rlabel metal2 8792 43680 8792 43680 0 _0204_
rlabel metal2 7896 44184 7896 44184 0 _0205_
rlabel metal2 10920 44128 10920 44128 0 _0206_
rlabel metal2 10528 44184 10528 44184 0 _0207_
rlabel metal2 12880 43736 12880 43736 0 _0208_
rlabel metal2 10920 23968 10920 23968 0 _0209_
rlabel metal2 13608 43288 13608 43288 0 _0210_
rlabel metal2 13216 43736 13216 43736 0 _0211_
rlabel metal2 43288 26320 43288 26320 0 _0212_
rlabel metal2 40488 24024 40488 24024 0 _0213_
rlabel metal2 42896 26376 42896 26376 0 _0214_
rlabel metal2 42168 24752 42168 24752 0 _0215_
rlabel metal2 46200 26040 46200 26040 0 _0216_
rlabel metal2 45192 25424 45192 25424 0 _0217_
rlabel metal3 46256 25480 46256 25480 0 _0218_
rlabel metal2 46984 25256 46984 25256 0 _0219_
rlabel metal2 41160 20664 41160 20664 0 _0220_
rlabel metal2 43512 24304 43512 24304 0 _0221_
rlabel metal2 45080 22624 45080 22624 0 _0222_
rlabel metal2 9296 2968 9296 2968 0 _0223_
rlabel metal2 42280 23296 42280 23296 0 _0224_
rlabel metal2 44016 22344 44016 22344 0 _0225_
rlabel metal2 44576 22232 44576 22232 0 _0226_
rlabel metal2 43624 22512 43624 22512 0 _0227_
rlabel metal2 41720 21056 41720 21056 0 _0228_
rlabel metal2 42840 21168 42840 21168 0 _0229_
rlabel metal2 44744 18704 44744 18704 0 _0230_
rlabel metal3 43792 15288 43792 15288 0 _0231_
rlabel metal2 42728 15960 42728 15960 0 _0232_
rlabel metal2 43400 18032 43400 18032 0 _0233_
rlabel metal2 43176 15232 43176 15232 0 _0234_
rlabel metal2 43400 17584 43400 17584 0 _0235_
rlabel metal2 43736 14112 43736 14112 0 _0236_
rlabel metal2 45080 16632 45080 16632 0 _0237_
rlabel metal3 46648 6552 46648 6552 0 _0238_
rlabel metal2 44744 7224 44744 7224 0 _0239_
rlabel metal2 43960 14112 43960 14112 0 _0240_
rlabel metal2 47544 5824 47544 5824 0 _0241_
rlabel metal2 45080 6832 45080 6832 0 _0242_
rlabel metal2 44744 6384 44744 6384 0 _0243_
rlabel metal3 47432 5096 47432 5096 0 _0244_
rlabel metal2 46480 5096 46480 5096 0 _0245_
rlabel metal3 47432 6664 47432 6664 0 _0246_
rlabel metal2 47320 6944 47320 6944 0 _0247_
rlabel metal2 46648 8344 46648 8344 0 _0248_
rlabel metal3 46928 11256 46928 11256 0 _0249_
rlabel metal2 47096 8904 47096 8904 0 _0250_
rlabel metal2 46536 13384 46536 13384 0 _0251_
rlabel metal2 47712 11368 47712 11368 0 _0252_
rlabel metal2 46816 10808 46816 10808 0 _0253_
rlabel metal2 46088 10864 46088 10864 0 _0254_
rlabel metal2 45752 11480 45752 11480 0 _0255_
rlabel metal2 45416 12040 45416 12040 0 _0256_
rlabel metal2 47208 11144 47208 11144 0 _0257_
rlabel metal2 47208 12152 47208 12152 0 _0258_
rlabel metal3 47432 13720 47432 13720 0 _0259_
rlabel metal3 47432 15288 47432 15288 0 _0260_
rlabel metal2 47768 15064 47768 15064 0 _0261_
rlabel metal2 47208 18368 47208 18368 0 _0262_
rlabel metal2 45976 16464 45976 16464 0 _0263_
rlabel metal2 47768 16184 47768 16184 0 _0264_
rlabel metal2 47208 16184 47208 16184 0 _0265_
rlabel metal2 47096 19152 47096 19152 0 _0266_
rlabel metal2 46760 18032 46760 18032 0 _0267_
rlabel metal2 46256 18424 46256 18424 0 _0268_
rlabel metal2 46424 18144 46424 18144 0 _0269_
rlabel metal3 45416 17528 45416 17528 0 _0270_
rlabel metal2 43512 16856 43512 16856 0 _0271_
rlabel metal2 39032 18200 39032 18200 0 _0272_
rlabel metal2 41720 16016 41720 16016 0 _0273_
rlabel metal2 42392 16128 42392 16128 0 _0274_
rlabel via2 47544 23240 47544 23240 0 _0275_
rlabel metal2 47208 21616 47208 21616 0 _0276_
rlabel metal2 46984 20832 46984 20832 0 _0277_
rlabel metal2 47544 20776 47544 20776 0 _0278_
rlabel metal2 47656 24136 47656 24136 0 _0279_
rlabel metal2 48216 23016 48216 23016 0 _0280_
rlabel metal2 22344 11256 22344 11256 0 _0281_
rlabel metal2 41888 12264 41888 12264 0 _0282_
rlabel metal2 41160 24584 41160 24584 0 _0283_
rlabel metal2 47544 21896 47544 21896 0 _0284_
rlabel metal3 41496 16744 41496 16744 0 _0285_
rlabel metal3 25928 14112 25928 14112 0 _0286_
rlabel metal3 20440 1288 20440 1288 0 _0287_
rlabel metal2 26320 5880 26320 5880 0 _0288_
rlabel metal2 21448 8232 21448 8232 0 _0289_
rlabel metal2 38696 13664 38696 13664 0 _0290_
rlabel metal2 39592 14392 39592 14392 0 _0291_
rlabel metal2 39984 16632 39984 16632 0 _0292_
rlabel metal3 40096 15512 40096 15512 0 _0293_
rlabel metal2 39704 15624 39704 15624 0 _0294_
rlabel metal2 38528 20104 38528 20104 0 _0295_
rlabel metal3 38724 20104 38724 20104 0 _0296_
rlabel metal2 41384 8288 41384 8288 0 _0297_
rlabel metal2 38136 18424 38136 18424 0 _0298_
rlabel metal2 37688 21616 37688 21616 0 _0299_
rlabel metal3 36848 21672 36848 21672 0 _0300_
rlabel metal2 38248 22008 38248 22008 0 _0301_
rlabel via2 39032 22232 39032 22232 0 _0302_
rlabel metal2 40600 22736 40600 22736 0 _0303_
rlabel metal3 40376 21448 40376 21448 0 _0304_
rlabel metal2 38248 25144 38248 25144 0 _0305_
rlabel metal2 37912 24640 37912 24640 0 _0306_
rlabel metal2 36456 26208 36456 26208 0 _0307_
rlabel metal3 37240 26264 37240 26264 0 _0308_
rlabel metal2 37576 26264 37576 26264 0 _0309_
rlabel metal3 38668 26488 38668 26488 0 _0310_
rlabel metal2 37912 26376 37912 26376 0 _0311_
rlabel metal2 35728 28616 35728 28616 0 _0312_
rlabel metal2 35336 28560 35336 28560 0 _0313_
rlabel metal3 36512 28616 36512 28616 0 _0314_
rlabel metal2 35448 15568 35448 15568 0 _0315_
rlabel metal3 35560 28840 35560 28840 0 _0316_
rlabel metal2 35728 29400 35728 29400 0 _0317_
rlabel metal2 34888 31752 34888 31752 0 _0318_
rlabel metal2 34776 31920 34776 31920 0 _0319_
rlabel metal3 32872 30856 32872 30856 0 _0320_
rlabel metal2 32648 31248 32648 31248 0 _0321_
rlabel metal2 32760 34944 32760 34944 0 _0322_
rlabel metal3 32872 34888 32872 34888 0 _0323_
rlabel metal2 32984 34384 32984 34384 0 _0324_
rlabel metal2 33544 34384 33544 34384 0 _0325_
rlabel metal2 30072 35840 30072 35840 0 _0326_
rlabel metal2 30408 35280 30408 35280 0 _0327_
rlabel metal2 29176 35728 29176 35728 0 _0328_
rlabel metal3 28112 36344 28112 36344 0 _0329_
rlabel metal2 32984 22904 32984 22904 0 _0330_
rlabel metal3 28504 35784 28504 35784 0 _0331_
rlabel metal3 26852 35560 26852 35560 0 _0332_
rlabel metal2 28056 35952 28056 35952 0 _0333_
rlabel metal2 26264 38724 26264 38724 0 _0334_
rlabel metal2 28000 37912 28000 37912 0 _0335_
rlabel metal2 25592 38752 25592 38752 0 _0336_
rlabel metal2 27384 38808 27384 38808 0 _0337_
rlabel metal2 27160 40376 27160 40376 0 _0338_
rlabel metal2 27496 41272 27496 41272 0 _0339_
rlabel metal2 27216 40600 27216 40600 0 _0340_
rlabel metal2 26432 42168 26432 42168 0 _0341_
rlabel metal3 26488 42616 26488 42616 0 _0342_
rlabel metal2 26712 42896 26712 42896 0 _0343_
rlabel metal2 27832 43960 27832 43960 0 _0344_
rlabel metal2 28168 43232 28168 43232 0 _0345_
rlabel metal2 25256 43904 25256 43904 0 _0346_
rlabel metal2 25648 43624 25648 43624 0 _0347_
rlabel metal2 25480 44576 25480 44576 0 _0348_
rlabel metal2 26040 44632 26040 44632 0 _0349_
rlabel metal3 25088 43512 25088 43512 0 _0350_
rlabel metal3 24696 43624 24696 43624 0 _0351_
rlabel metal2 24360 43456 24360 43456 0 _0352_
rlabel metal3 18872 1624 18872 1624 0 _0353_
rlabel metal2 42672 8232 42672 8232 0 _0354_
rlabel metal3 19544 2296 19544 2296 0 _0355_
rlabel metal2 42280 9800 42280 9800 0 _0356_
rlabel metal2 38696 10024 38696 10024 0 _0357_
rlabel metal2 39704 9296 39704 9296 0 _0358_
rlabel metal2 40936 9520 40936 9520 0 _0359_
rlabel metal3 41720 8232 41720 8232 0 _0360_
rlabel metal2 23688 2856 23688 2856 0 _0361_
rlabel metal2 41272 7616 41272 7616 0 _0362_
rlabel metal2 40376 8008 40376 8008 0 _0363_
rlabel metal2 42840 7784 42840 7784 0 _0364_
rlabel metal3 17696 1400 17696 1400 0 _0365_
rlabel metal2 34496 2632 34496 2632 0 _0366_
rlabel metal3 40600 7672 40600 7672 0 _0367_
rlabel metal2 42504 5824 42504 5824 0 _0368_
rlabel metal2 40040 8680 40040 8680 0 _0369_
rlabel metal2 39816 7840 39816 7840 0 _0370_
rlabel metal2 41944 7728 41944 7728 0 _0371_
rlabel metal2 41160 5936 41160 5936 0 _0372_
rlabel metal2 38584 9912 38584 9912 0 _0373_
rlabel metal2 38864 8232 38864 8232 0 _0374_
rlabel metal3 39088 7672 39088 7672 0 _0375_
rlabel metal2 39480 7112 39480 7112 0 _0376_
rlabel metal3 37184 6552 37184 6552 0 _0377_
rlabel metal2 39592 6216 39592 6216 0 _0378_
rlabel metal2 38136 8344 38136 8344 0 _0379_
rlabel metal3 38024 7224 38024 7224 0 _0380_
rlabel metal2 33544 6776 33544 6776 0 _0381_
rlabel metal2 38808 7112 38808 7112 0 _0382_
rlabel metal2 39592 4928 39592 4928 0 _0383_
rlabel metal2 36456 6048 36456 6048 0 _0384_
rlabel metal2 36848 7560 36848 7560 0 _0385_
rlabel metal2 35896 7840 35896 7840 0 _0386_
rlabel metal2 35840 5880 35840 5880 0 _0387_
rlabel metal2 37128 5488 37128 5488 0 _0388_
rlabel metal3 35784 10696 35784 10696 0 _0389_
rlabel metal2 35112 7560 35112 7560 0 _0390_
rlabel metal2 35448 6720 35448 6720 0 _0391_
rlabel metal2 35504 11928 35504 11928 0 _0392_
rlabel metal2 35448 6888 35448 6888 0 _0393_
rlabel metal2 36064 5208 36064 5208 0 _0394_
rlabel metal3 37016 11592 37016 11592 0 _0395_
rlabel metal2 23352 11312 23352 11312 0 _0396_
rlabel metal2 34776 11816 34776 11816 0 _0397_
rlabel metal3 34832 11368 34832 11368 0 _0398_
rlabel metal2 34888 11760 34888 11760 0 _0399_
rlabel metal3 35224 12152 35224 12152 0 _0400_
rlabel metal2 34104 13384 34104 13384 0 _0401_
rlabel metal3 34776 12936 34776 12936 0 _0402_
rlabel metal2 22960 6440 22960 6440 0 _0403_
rlabel metal2 34608 13160 34608 13160 0 _0404_
rlabel metal2 35560 13216 35560 13216 0 _0405_
rlabel metal2 33768 20776 33768 20776 0 _0406_
rlabel metal2 34104 14896 34104 14896 0 _0407_
rlabel metal2 35056 15288 35056 15288 0 _0408_
rlabel metal2 33208 21952 33208 21952 0 _0409_
rlabel metal2 34552 9408 34552 9408 0 _0410_
rlabel metal2 29904 6104 29904 6104 0 _0411_
rlabel metal2 23128 7896 23128 7896 0 _0412_
rlabel metal2 26488 7728 26488 7728 0 _0413_
rlabel metal2 32312 7728 32312 7728 0 _0414_
rlabel metal3 34832 8120 34832 8120 0 _0415_
rlabel metal3 32312 6664 32312 6664 0 _0416_
rlabel metal2 32200 5488 32200 5488 0 _0417_
rlabel metal2 33152 5880 33152 5880 0 _0418_
rlabel metal2 24808 5208 24808 5208 0 _0419_
rlabel metal2 35112 5432 35112 5432 0 _0420_
rlabel metal2 31752 6440 31752 6440 0 _0421_
rlabel metal2 24416 6104 24416 6104 0 _0422_
rlabel metal2 31976 4536 31976 4536 0 _0423_
rlabel metal2 31416 4816 31416 4816 0 _0424_
rlabel metal3 20720 4984 20720 4984 0 _0425_
rlabel metal3 24696 7560 24696 7560 0 _0426_
rlabel metal3 24752 5880 24752 5880 0 _0427_
rlabel metal2 22344 5824 22344 5824 0 _0428_
rlabel metal2 18648 5936 18648 5936 0 _0429_
rlabel metal2 24304 5320 24304 5320 0 _0430_
rlabel metal2 25200 4424 25200 4424 0 _0431_
rlabel metal2 22120 6272 22120 6272 0 _0432_
rlabel metal2 20216 5824 20216 5824 0 _0433_
rlabel metal2 22176 5320 22176 5320 0 _0434_
rlabel metal2 22232 3696 22232 3696 0 _0435_
rlabel metal2 19992 5992 19992 5992 0 _0436_
rlabel metal2 19768 7672 19768 7672 0 _0437_
rlabel metal3 19432 5320 19432 5320 0 _0438_
rlabel metal2 19992 4928 19992 4928 0 _0439_
rlabel metal2 19656 4368 19656 4368 0 _0440_
rlabel metal2 21784 8568 21784 8568 0 _0441_
rlabel metal2 19544 8568 19544 8568 0 _0442_
rlabel metal3 20216 7224 20216 7224 0 _0443_
rlabel metal3 21336 10696 21336 10696 0 _0444_
rlabel metal2 20384 7448 20384 7448 0 _0445_
rlabel metal3 20104 7560 20104 7560 0 _0446_
rlabel metal2 23352 9688 23352 9688 0 _0447_
rlabel metal2 21952 11144 21952 11144 0 _0448_
rlabel metal2 23240 11592 23240 11592 0 _0449_
rlabel metal2 23296 10696 23296 10696 0 _0450_
rlabel metal3 22064 10584 22064 10584 0 _0451_
rlabel metal3 22400 13720 22400 13720 0 _0452_
rlabel metal2 23352 13776 23352 13776 0 _0453_
rlabel metal2 22232 12208 22232 12208 0 _0454_
rlabel metal2 22456 12880 22456 12880 0 _0455_
rlabel metal2 25760 17640 25760 17640 0 _0456_
rlabel metal3 12264 2856 12264 2856 0 _0457_
rlabel metal2 22120 16184 22120 16184 0 _0458_
rlabel metal2 23184 14392 23184 14392 0 _0459_
rlabel metal3 21000 23352 21000 23352 0 _0460_
rlabel metal2 3640 17192 3640 17192 0 _0461_
rlabel metal2 14280 9352 14280 9352 0 _0462_
rlabel metal2 12208 6664 12208 6664 0 _0463_
rlabel metal2 9800 7784 9800 7784 0 _0464_
rlabel metal3 10640 7672 10640 7672 0 _0465_
rlabel metal2 12824 8456 12824 8456 0 _0466_
rlabel metal3 15008 9016 15008 9016 0 _0467_
rlabel metal2 8680 5488 8680 5488 0 _0468_
rlabel metal3 14000 6104 14000 6104 0 _0469_
rlabel metal2 12656 5656 12656 5656 0 _0470_
rlabel metal2 13552 5320 13552 5320 0 _0471_
rlabel metal2 13272 4256 13272 4256 0 _0472_
rlabel metal3 10584 5880 10584 5880 0 _0473_
rlabel metal2 8568 6160 8568 6160 0 _0474_
rlabel metal3 10360 6104 10360 6104 0 _0475_
rlabel metal2 10360 5656 10360 5656 0 _0476_
rlabel metal2 10360 3976 10360 3976 0 _0477_
rlabel metal2 10024 8344 10024 8344 0 _0478_
rlabel metal3 8848 6440 8848 6440 0 _0479_
rlabel metal3 6664 6104 6664 6104 0 _0480_
rlabel metal2 8008 6328 8008 6328 0 _0481_
rlabel metal3 8120 5992 8120 5992 0 _0482_
rlabel metal2 7672 4536 7672 4536 0 _0483_
rlabel metal3 6776 6440 6776 6440 0 _0484_
rlabel metal3 7560 7560 7560 7560 0 _0485_
rlabel metal2 7336 5544 7336 5544 0 _0486_
rlabel metal2 5768 5264 5768 5264 0 _0487_
rlabel metal2 7000 7840 7000 7840 0 _0488_
rlabel metal2 7336 9352 7336 9352 0 _0489_
rlabel metal2 7112 8232 7112 8232 0 _0490_
rlabel metal3 6944 8120 6944 8120 0 _0491_
rlabel metal3 10192 12936 10192 12936 0 _0492_
rlabel metal2 7672 9352 7672 9352 0 _0493_
rlabel metal2 7448 8848 7448 8848 0 _0494_
rlabel metal2 8568 11424 8568 11424 0 _0495_
rlabel metal2 8904 9296 8904 9296 0 _0496_
rlabel metal2 4984 8624 4984 8624 0 _0497_
rlabel metal2 12824 10640 12824 10640 0 _0498_
rlabel metal2 9240 11368 9240 11368 0 _0499_
rlabel metal2 13160 11872 13160 11872 0 _0500_
rlabel metal3 11648 11256 11648 11256 0 _0501_
rlabel metal2 11816 11200 11816 11200 0 _0502_
rlabel metal2 11816 12432 11816 12432 0 _0503_
rlabel metal2 11536 15288 11536 15288 0 _0504_
rlabel metal2 13048 12320 13048 12320 0 _0505_
rlabel metal2 12096 12376 12096 12376 0 _0506_
rlabel metal2 9632 21560 9632 21560 0 _0507_
rlabel metal3 10360 14616 10360 14616 0 _0508_
rlabel metal3 12656 15176 12656 15176 0 _0509_
rlabel metal2 9744 21784 9744 21784 0 _0510_
rlabel metal2 39928 28896 39928 28896 0 _0511_
rlabel metal2 37800 29568 37800 29568 0 _0512_
rlabel metal2 40264 29344 40264 29344 0 _0513_
rlabel metal2 29400 28728 29400 28728 0 _0514_
rlabel metal2 31640 29456 31640 29456 0 _0515_
rlabel metal2 42112 28504 42112 28504 0 _0516_
rlabel metal2 39032 28168 39032 28168 0 _0517_
rlabel metal3 42224 29288 42224 29288 0 _0518_
rlabel metal2 41720 28784 41720 28784 0 _0519_
rlabel metal2 41160 31024 41160 31024 0 _0520_
rlabel metal2 38808 33544 38808 33544 0 _0521_
rlabel metal2 41496 32704 41496 32704 0 _0522_
rlabel metal3 40600 32648 40600 32648 0 _0523_
rlabel metal2 38304 33096 38304 33096 0 _0524_
rlabel metal2 37912 33208 37912 33208 0 _0525_
rlabel metal2 38360 33712 38360 33712 0 _0526_
rlabel metal2 38808 35784 38808 35784 0 _0527_
rlabel metal2 37352 32312 37352 32312 0 _0528_
rlabel metal2 36120 33264 36120 33264 0 _0529_
rlabel metal2 36176 33544 36176 33544 0 _0530_
rlabel metal2 35000 35336 35000 35336 0 _0531_
rlabel metal2 35896 34160 35896 34160 0 _0532_
rlabel metal2 36344 34720 36344 34720 0 _0533_
rlabel metal3 35448 36344 35448 36344 0 _0534_
rlabel metal2 37016 35504 37016 35504 0 _0535_
rlabel metal2 39592 36176 39592 36176 0 _0536_
rlabel metal2 35000 38724 35000 38724 0 _0537_
rlabel metal2 34776 38724 34776 38724 0 _0538_
rlabel metal2 24024 42336 24024 42336 0 _0539_
rlabel metal2 34944 38360 34944 38360 0 _0540_
rlabel metal2 40768 24696 40768 24696 0 _0541_
rlabel metal2 37240 37520 37240 37520 0 _0542_
rlabel metal2 37184 39592 37184 39592 0 _0543_
rlabel metal2 36624 38808 36624 38808 0 _0544_
rlabel metal3 36904 38752 36904 38752 0 _0545_
rlabel metal2 39648 38696 39648 38696 0 _0546_
rlabel metal2 37800 40768 37800 40768 0 _0547_
rlabel metal2 38024 40376 38024 40376 0 _0548_
rlabel metal2 36232 40600 36232 40600 0 _0549_
rlabel metal2 39032 43288 39032 43288 0 _0550_
rlabel metal2 35896 40992 35896 40992 0 _0551_
rlabel metal2 36456 40768 36456 40768 0 _0552_
rlabel metal2 38696 41272 38696 41272 0 _0553_
rlabel metal2 38024 41272 38024 41272 0 _0554_
rlabel metal2 38472 41496 38472 41496 0 _0555_
rlabel metal2 38696 41888 38696 41888 0 _0556_
rlabel metal2 38808 42616 38808 42616 0 _0557_
rlabel metal2 39928 44632 39928 44632 0 _0558_
rlabel metal3 35952 42616 35952 42616 0 _0559_
rlabel metal3 38920 42112 38920 42112 0 _0560_
rlabel metal2 40152 44128 40152 44128 0 _0561_
rlabel metal2 39816 44632 39816 44632 0 _0562_
rlabel metal2 38808 42168 38808 42168 0 _0563_
rlabel metal2 39648 41944 39648 41944 0 _0564_
rlabel metal2 43512 41608 43512 41608 0 _0565_
rlabel metal2 44184 42504 44184 42504 0 _0566_
rlabel metal3 47880 40376 47880 40376 0 _0567_
rlabel metal3 45472 42504 45472 42504 0 _0568_
rlabel metal2 46872 37296 46872 37296 0 _0569_
rlabel metal2 43512 42616 43512 42616 0 _0570_
rlabel metal2 44632 44408 44632 44408 0 _0571_
rlabel metal2 44408 45248 44408 45248 0 _0572_
rlabel metal2 45752 34552 45752 34552 0 _0573_
rlabel metal2 44856 36512 44856 36512 0 _0574_
rlabel metal2 45472 29960 45472 29960 0 _0575_
rlabel metal2 45304 30632 45304 30632 0 _0576_
rlabel metal2 46872 29792 46872 29792 0 _0577_
rlabel metal2 47432 33152 47432 33152 0 _0578_
rlabel metal2 46144 34104 46144 34104 0 _0579_
rlabel metal3 46872 33208 46872 33208 0 _0580_
rlabel metal2 43288 39200 43288 39200 0 _0581_
rlabel metal2 44184 31416 44184 31416 0 _0582_
rlabel metal2 46256 31752 46256 31752 0 _0583_
rlabel metal2 44408 31304 44408 31304 0 _0584_
rlabel metal2 41720 37520 41720 37520 0 _0585_
rlabel metal2 41048 34608 41048 34608 0 _0586_
rlabel metal2 39144 34776 39144 34776 0 _0587_
rlabel metal3 40376 35896 40376 35896 0 _0588_
rlabel metal2 43064 36680 43064 36680 0 _0589_
rlabel metal2 43400 40096 43400 40096 0 _0590_
rlabel metal2 42560 35000 42560 35000 0 _0591_
rlabel metal2 39256 36400 39256 36400 0 _0592_
rlabel metal2 42056 39648 42056 39648 0 _0593_
rlabel metal2 41048 37520 41048 37520 0 _0594_
rlabel metal2 44296 39200 44296 39200 0 _0595_
rlabel metal2 46312 41160 46312 41160 0 _0596_
rlabel metal2 41776 39592 41776 39592 0 _0597_
rlabel metal2 40208 41832 40208 41832 0 _0598_
rlabel metal2 40936 40376 40936 40376 0 _0599_
rlabel metal2 40824 39928 40824 39928 0 _0600_
rlabel metal3 46480 40376 46480 40376 0 _0601_
rlabel metal2 43904 39368 43904 39368 0 _0602_
rlabel metal3 46928 40488 46928 40488 0 _0603_
rlabel metal2 23128 16856 23128 16856 0 _0604_
rlabel metal3 18760 10752 18760 10752 0 _0605_
rlabel metal3 19096 15960 19096 15960 0 _0606_
rlabel metal2 17080 15680 17080 15680 0 _0607_
rlabel metal2 23576 19096 23576 19096 0 _0608_
rlabel metal2 19432 16800 19432 16800 0 _0609_
rlabel metal3 22344 15848 22344 15848 0 _0610_
rlabel metal2 28056 13216 28056 13216 0 _0611_
rlabel metal3 27944 16072 27944 16072 0 _0612_
rlabel metal2 29736 14616 29736 14616 0 _0613_
rlabel metal2 17192 11648 17192 11648 0 _0614_
rlabel metal2 29064 12208 29064 12208 0 _0615_
rlabel metal2 26936 10920 26936 10920 0 _0616_
rlabel metal3 25928 14280 25928 14280 0 _0617_
rlabel metal3 28840 12152 28840 12152 0 _0618_
rlabel metal2 28616 12600 28616 12600 0 _0619_
rlabel metal2 16632 14000 16632 14000 0 _0620_
rlabel metal2 26488 13048 26488 13048 0 _0621_
rlabel metal3 25312 17640 25312 17640 0 _0622_
rlabel metal2 1960 12432 1960 12432 0 _0623_
rlabel metal2 25144 12600 25144 12600 0 _0624_
rlabel metal2 26376 15736 26376 15736 0 _0625_
rlabel metal2 15456 17528 15456 17528 0 _0626_
rlabel metal2 17976 16464 17976 16464 0 _0627_
rlabel metal2 16912 15848 16912 15848 0 _0628_
rlabel metal2 17640 12040 17640 12040 0 _0629_
rlabel metal3 17024 10808 17024 10808 0 _0630_
rlabel metal2 15512 10640 15512 10640 0 _0631_
rlabel metal2 24248 19040 24248 19040 0 _0632_
rlabel metal3 18536 10584 18536 10584 0 _0633_
rlabel metal2 1064 17528 1064 17528 0 _0634_
rlabel metal3 16128 12376 16128 12376 0 _0635_
rlabel metal2 18200 12320 18200 12320 0 _0636_
rlabel metal2 17976 19320 17976 19320 0 _0637_
rlabel metal2 9576 12432 9576 12432 0 _0638_
rlabel metal2 15624 12208 15624 12208 0 _0639_
rlabel metal2 18648 12544 18648 12544 0 _0640_
rlabel metal2 19768 12376 19768 12376 0 _0641_
rlabel metal3 17528 15456 17528 15456 0 _0642_
rlabel metal2 5544 14616 5544 14616 0 _0643_
rlabel metal3 6496 15400 6496 15400 0 _0644_
rlabel metal3 6552 11368 6552 11368 0 _0645_
rlabel metal2 7112 14224 7112 14224 0 _0646_
rlabel metal2 7448 11144 7448 11144 0 _0647_
rlabel metal3 6328 14280 6328 14280 0 _0648_
rlabel metal3 6552 14392 6552 14392 0 _0649_
rlabel metal2 6664 13216 6664 13216 0 _0650_
rlabel metal2 8008 13608 8008 13608 0 _0651_
rlabel metal3 18256 16856 18256 16856 0 _0652_
rlabel metal3 8344 15288 8344 15288 0 _0653_
rlabel metal2 2632 15512 2632 15512 0 _0654_
rlabel metal2 21336 14280 21336 14280 0 _0655_
rlabel metal2 23912 14616 23912 14616 0 _0656_
rlabel metal2 23912 14112 23912 14112 0 _0657_
rlabel metal3 18928 17640 18928 17640 0 _0658_
rlabel metal2 21224 13160 21224 13160 0 _0659_
rlabel metal2 21672 18312 21672 18312 0 _0660_
rlabel metal3 22008 19208 22008 19208 0 _0661_
rlabel metal2 22792 19152 22792 19152 0 _0662_
rlabel metal2 24360 19096 24360 19096 0 _0663_
rlabel metal2 24360 20552 24360 20552 0 _0664_
rlabel metal3 21336 21560 21336 21560 0 _0665_
rlabel metal3 21336 17864 21336 17864 0 _0666_
rlabel metal2 23800 18480 23800 18480 0 _0667_
rlabel metal2 19880 18144 19880 18144 0 _0668_
rlabel metal3 14336 10808 14336 10808 0 _0669_
rlabel metal3 20664 18312 20664 18312 0 _0670_
rlabel metal2 22400 17640 22400 17640 0 _0671_
rlabel metal2 19096 19936 19096 19936 0 _0672_
rlabel metal2 19096 22512 19096 22512 0 _0673_
rlabel metal2 16744 20384 16744 20384 0 _0674_
rlabel metal2 17416 14672 17416 14672 0 _0675_
rlabel metal2 1400 16968 1400 16968 0 _0676_
rlabel metal3 16688 23576 16688 23576 0 _0677_
rlabel metal2 18424 19712 18424 19712 0 _0678_
rlabel metal2 18816 16744 18816 16744 0 _0679_
rlabel metal2 18312 18928 18312 18928 0 _0680_
rlabel metal2 9520 2744 9520 2744 0 _0681_
rlabel metal2 5992 16632 5992 16632 0 _0682_
rlabel metal2 4872 13496 4872 13496 0 _0683_
rlabel metal3 5096 16632 5096 16632 0 _0684_
rlabel metal2 5208 16800 5208 16800 0 _0685_
rlabel metal2 6776 16016 6776 16016 0 _0686_
rlabel metal3 5992 15960 5992 15960 0 _0687_
rlabel metal2 4648 16296 4648 16296 0 _0688_
rlabel metal3 17584 14504 17584 14504 0 _0689_
rlabel metal3 15820 14728 15820 14728 0 _0690_
rlabel metal2 7896 18256 7896 18256 0 _0691_
rlabel metal2 10528 16184 10528 16184 0 _0692_
rlabel metal3 7840 17976 7840 17976 0 _0693_
rlabel metal2 10808 17808 10808 17808 0 _0694_
rlabel metal2 3192 14448 3192 14448 0 _0695_
rlabel metal3 13328 16296 13328 16296 0 _0696_
rlabel metal2 7560 16324 7560 16324 0 _0697_
rlabel metal2 11816 17584 11816 17584 0 _0698_
rlabel metal3 13552 14392 13552 14392 0 _0699_
rlabel metal3 16632 16744 16632 16744 0 _0700_
rlabel metal3 12936 17752 12936 17752 0 _0701_
rlabel metal2 33096 18704 33096 18704 0 _0702_
rlabel metal2 31192 18088 31192 18088 0 _0703_
rlabel metal3 31696 16856 31696 16856 0 _0704_
rlabel metal2 31864 19152 31864 19152 0 _0705_
rlabel metal2 34104 18032 34104 18032 0 _0706_
rlabel metal3 33936 17528 33936 17528 0 _0707_
rlabel metal2 1512 19600 1512 19600 0 _0708_
rlabel metal2 23240 27440 23240 27440 0 _0709_
rlabel metal2 21224 20104 21224 20104 0 _0710_
rlabel metal3 18368 28728 18368 28728 0 _0711_
rlabel metal3 21336 25592 21336 25592 0 _0712_
rlabel metal2 22680 24976 22680 24976 0 _0713_
rlabel metal2 23240 25984 23240 25984 0 _0714_
rlabel metal2 15512 24472 15512 24472 0 _0715_
rlabel metal2 21168 26712 21168 26712 0 _0716_
rlabel metal2 19992 24864 19992 24864 0 _0717_
rlabel metal3 19656 26040 19656 26040 0 _0718_
rlabel metal2 23576 34160 23576 34160 0 _0719_
rlabel metal2 25872 35560 25872 35560 0 _0720_
rlabel metal3 23744 27048 23744 27048 0 _0721_
rlabel metal3 24472 27160 24472 27160 0 _0722_
rlabel metal3 20440 19992 20440 19992 0 _0723_
rlabel metal3 21000 23912 21000 23912 0 _0724_
rlabel metal2 19544 25200 19544 25200 0 _0725_
rlabel metal3 17360 28504 17360 28504 0 _0726_
rlabel metal2 22792 28952 22792 28952 0 _0727_
rlabel metal2 29400 27552 29400 27552 0 _0728_
rlabel metal3 30016 19208 30016 19208 0 _0729_
rlabel metal2 26040 20664 26040 20664 0 _0730_
rlabel metal2 30128 20888 30128 20888 0 _0731_
rlabel metal2 24584 21448 24584 21448 0 _0732_
rlabel metal2 25480 21784 25480 21784 0 _0733_
rlabel metal2 43064 17808 43064 17808 0 _0734_
rlabel metal2 25032 25704 25032 25704 0 _0735_
rlabel metal2 32088 20440 32088 20440 0 _0736_
rlabel metal2 25592 20832 25592 20832 0 _0737_
rlabel metal3 31808 21560 31808 21560 0 _0738_
rlabel metal2 39704 19096 39704 19096 0 _0739_
rlabel metal2 29624 24080 29624 24080 0 _0740_
rlabel metal2 28504 20832 28504 20832 0 _0741_
rlabel metal2 27496 26320 27496 26320 0 _0742_
rlabel metal2 27272 26208 27272 26208 0 _0743_
rlabel metal2 24696 17080 24696 17080 0 _0744_
rlabel metal2 26264 22848 26264 22848 0 _0745_
rlabel metal2 25480 21336 25480 21336 0 _0746_
rlabel metal2 24584 23688 24584 23688 0 _0747_
rlabel metal3 28896 27048 28896 27048 0 _0748_
rlabel metal2 31080 28728 31080 28728 0 _0749_
rlabel metal2 16632 23296 16632 23296 0 _0750_
rlabel metal2 17640 24304 17640 24304 0 _0751_
rlabel metal3 12768 20776 12768 20776 0 _0752_
rlabel via2 11704 23464 11704 23464 0 _0753_
rlabel metal2 10584 19880 10584 19880 0 _0754_
rlabel metal3 7112 18200 7112 18200 0 _0755_
rlabel metal2 12600 25200 12600 25200 0 _0756_
rlabel metal3 11928 26152 11928 26152 0 _0757_
rlabel metal3 17192 21336 17192 21336 0 _0758_
rlabel metal3 11984 26264 11984 26264 0 _0759_
rlabel metal2 17528 26544 17528 26544 0 _0760_
rlabel metal3 13832 26376 13832 26376 0 _0761_
rlabel metal2 15624 24192 15624 24192 0 _0762_
rlabel metal2 3192 15960 3192 15960 0 _0763_
rlabel metal3 10192 24024 10192 24024 0 _0764_
rlabel metal2 18760 37184 18760 37184 0 _0765_
rlabel metal2 11648 24136 11648 24136 0 _0766_
rlabel metal2 6664 24696 6664 24696 0 _0767_
rlabel metal2 2856 23296 2856 23296 0 _0768_
rlabel metal2 6216 24472 6216 24472 0 _0769_
rlabel metal2 7000 25872 7000 25872 0 _0770_
rlabel metal3 5992 19880 5992 19880 0 _0771_
rlabel metal2 6440 25592 6440 25592 0 _0772_
rlabel metal2 6104 28056 6104 28056 0 _0773_
rlabel metal2 10248 20720 10248 20720 0 _0774_
rlabel metal2 9464 25256 9464 25256 0 _0775_
rlabel metal2 9016 25200 9016 25200 0 _0776_
rlabel metal2 4984 16800 4984 16800 0 _0777_
rlabel metal2 1344 15288 1344 15288 0 _0778_
rlabel metal3 6832 26376 6832 26376 0 _0779_
rlabel metal2 1960 18592 1960 18592 0 _0780_
rlabel metal2 2408 24528 2408 24528 0 _0781_
rlabel metal2 8400 22792 8400 22792 0 _0782_
rlabel metal2 3192 23128 3192 23128 0 _0783_
rlabel metal2 8680 28616 8680 28616 0 _0784_
rlabel metal2 16408 25592 16408 25592 0 _0785_
rlabel metal2 27832 28336 27832 28336 0 _0786_
rlabel metal2 29848 29288 29848 29288 0 _0787_
rlabel metal3 30800 26264 30800 26264 0 _0788_
rlabel metal2 32200 26320 32200 26320 0 _0789_
rlabel metal2 32872 28840 32872 28840 0 _0790_
rlabel metal3 30856 29960 30856 29960 0 _0791_
rlabel metal3 21448 26264 21448 26264 0 _0792_
rlabel metal2 21560 25984 21560 25984 0 _0793_
rlabel metal2 22904 26432 22904 26432 0 _0794_
rlabel metal2 30744 21168 30744 21168 0 _0795_
rlabel metal2 30856 23576 30856 23576 0 _0796_
rlabel metal2 31304 26096 31304 26096 0 _0797_
rlabel metal2 30408 23184 30408 23184 0 _0798_
rlabel metal2 31192 24640 31192 24640 0 _0799_
rlabel metal2 30296 24304 30296 24304 0 _0800_
rlabel metal2 31864 25424 31864 25424 0 _0801_
rlabel metal3 30296 29512 30296 29512 0 _0802_
rlabel metal3 24248 27664 24248 27664 0 _0803_
rlabel metal2 15288 20104 15288 20104 0 _0804_
rlabel metal2 16296 26096 16296 26096 0 _0805_
rlabel metal2 18536 21616 18536 21616 0 _0806_
rlabel metal3 18368 21784 18368 21784 0 _0807_
rlabel metal3 17472 27944 17472 27944 0 _0808_
rlabel metal3 18816 24696 18816 24696 0 _0809_
rlabel metal2 17472 24920 17472 24920 0 _0810_
rlabel metal3 1960 30072 1960 30072 0 _0811_
rlabel metal2 7952 16184 7952 16184 0 _0812_
rlabel metal2 5208 27776 5208 27776 0 _0813_
rlabel metal2 7784 20496 7784 20496 0 _0814_
rlabel metal2 3080 25144 3080 25144 0 _0815_
rlabel metal2 2744 22624 2744 22624 0 _0816_
rlabel metal2 6328 22232 6328 22232 0 _0817_
rlabel metal2 10136 28448 10136 28448 0 _0818_
rlabel metal2 12936 29232 12936 29232 0 _0819_
rlabel metal2 32704 30184 32704 30184 0 _0820_
rlabel metal2 31640 31024 31640 31024 0 _0821_
rlabel metal2 32312 24864 32312 24864 0 _0822_
rlabel metal2 29960 24976 29960 24976 0 _0823_
rlabel metal2 31416 30520 31416 30520 0 _0824_
rlabel metal2 8680 23184 8680 23184 0 _0825_
rlabel metal2 17976 34328 17976 34328 0 _0826_
rlabel metal2 16072 26572 16072 26572 0 _0827_
rlabel metal2 15736 26600 15736 26600 0 _0828_
rlabel metal2 16520 26264 16520 26264 0 _0829_
rlabel metal2 17752 34608 17752 34608 0 _0830_
rlabel metal2 2632 24416 2632 24416 0 _0831_
rlabel metal2 2128 27160 2128 27160 0 _0832_
rlabel metal2 1792 22456 1792 22456 0 _0833_
rlabel metal2 6664 25704 6664 25704 0 _0834_
rlabel metal2 6776 29288 6776 29288 0 _0835_
rlabel metal3 6888 30184 6888 30184 0 _0836_
rlabel metal2 6216 29176 6216 29176 0 _0837_
rlabel metal4 1736 30912 1736 30912 0 _0838_
rlabel metal3 7000 28336 7000 28336 0 _0839_
rlabel metal3 16408 27720 16408 27720 0 _0840_
rlabel metal2 15064 18144 15064 18144 0 _0841_
rlabel metal2 19096 24360 19096 24360 0 _0842_
rlabel metal2 15960 20216 15960 20216 0 _0843_
rlabel metal2 12264 32592 12264 32592 0 _0844_
rlabel metal2 13048 24304 13048 24304 0 _0845_
rlabel metal2 14336 29400 14336 29400 0 _0846_
rlabel metal2 16632 29960 16632 29960 0 _0847_
rlabel metal2 24024 31528 24024 31528 0 _0848_
rlabel metal2 26600 23576 26600 23576 0 _0849_
rlabel metal2 28056 20272 28056 20272 0 _0850_
rlabel metal2 26600 25816 26600 25816 0 _0851_
rlabel metal2 30296 23072 30296 23072 0 _0852_
rlabel metal2 27552 23800 27552 23800 0 _0853_
rlabel metal2 27048 23184 27048 23184 0 _0854_
rlabel metal3 28728 29400 28728 29400 0 _0855_
rlabel metal2 20216 29232 20216 29232 0 _0856_
rlabel metal2 20664 30016 20664 30016 0 _0857_
rlabel metal2 20440 29400 20440 29400 0 _0858_
rlabel metal2 21616 30184 21616 30184 0 _0859_
rlabel metal2 21728 25816 21728 25816 0 _0860_
rlabel metal2 22344 29792 22344 29792 0 _0861_
rlabel metal3 21784 29344 21784 29344 0 _0862_
rlabel metal2 28056 31416 28056 31416 0 _0863_
rlabel metal2 30520 31416 30520 31416 0 _0864_
rlabel metal2 29736 31248 29736 31248 0 _0865_
rlabel metal3 32032 30968 32032 30968 0 _0866_
rlabel metal2 30632 32368 30632 32368 0 _0867_
rlabel metal2 27496 30912 27496 30912 0 _0868_
rlabel metal3 28560 29512 28560 29512 0 _0869_
rlabel metal2 25704 28560 25704 28560 0 _0870_
rlabel metal2 28504 30296 28504 30296 0 _0871_
rlabel metal2 28504 32536 28504 32536 0 _0872_
rlabel metal3 24808 21560 24808 21560 0 _0873_
rlabel metal2 27944 22792 27944 22792 0 _0874_
rlabel metal2 25032 22232 25032 22232 0 _0875_
rlabel metal2 26040 30856 26040 30856 0 _0876_
rlabel metal2 19992 22904 19992 22904 0 _0877_
rlabel metal2 20888 29120 20888 29120 0 _0878_
rlabel metal2 18312 28448 18312 28448 0 _0879_
rlabel metal2 18872 29680 18872 29680 0 _0880_
rlabel metal2 23800 30688 23800 30688 0 _0881_
rlabel metal2 24416 33208 24416 33208 0 _0882_
rlabel metal2 5040 29512 5040 29512 0 _0883_
rlabel metal3 3696 29512 3696 29512 0 _0884_
rlabel metal2 16072 35056 16072 35056 0 _0885_
rlabel metal2 17472 28616 17472 28616 0 _0886_
rlabel metal2 13944 29176 13944 29176 0 _0887_
rlabel metal2 15064 24584 15064 24584 0 _0888_
rlabel metal3 16128 30184 16128 30184 0 _0889_
rlabel metal2 24920 32760 24920 32760 0 _0890_
rlabel metal2 16184 34664 16184 34664 0 _0891_
rlabel metal2 2800 32536 2800 32536 0 _0892_
rlabel metal2 15624 32424 15624 32424 0 _0893_
rlabel metal2 25592 32144 25592 32144 0 _0894_
rlabel metal2 26376 33152 26376 33152 0 _0895_
rlabel metal2 30744 32928 30744 32928 0 _0896_
rlabel metal2 29736 33376 29736 33376 0 _0897_
rlabel metal2 31080 34944 31080 34944 0 _0898_
rlabel metal2 25256 33376 25256 33376 0 _0899_
rlabel metal2 25592 31472 25592 31472 0 _0900_
rlabel metal2 22904 33376 22904 33376 0 _0901_
rlabel metal2 25816 32928 25816 32928 0 _0902_
rlabel metal2 29736 34048 29736 34048 0 _0903_
rlabel metal2 24136 29680 24136 29680 0 _0904_
rlabel metal3 23968 34104 23968 34104 0 _0905_
rlabel metal2 23800 24584 23800 24584 0 _0906_
rlabel metal2 26824 32928 26824 32928 0 _0907_
rlabel metal2 27720 34104 27720 34104 0 _0908_
rlabel metal2 13720 31696 13720 31696 0 _0909_
rlabel metal2 13832 31304 13832 31304 0 _0910_
rlabel metal2 16184 32144 16184 32144 0 _0911_
rlabel metal3 17024 31752 17024 31752 0 _0912_
rlabel metal2 13944 34496 13944 34496 0 _0913_
rlabel metal2 8344 33936 8344 33936 0 _0914_
rlabel metal2 15848 32480 15848 32480 0 _0915_
rlabel metal3 16968 32536 16968 32536 0 _0916_
rlabel metal2 16800 32536 16800 32536 0 _0917_
rlabel metal2 29512 34104 29512 34104 0 _0918_
rlabel metal2 30968 35896 30968 35896 0 _0919_
rlabel metal2 34496 36344 34496 36344 0 _0920_
rlabel metal2 29792 35112 29792 35112 0 _0921_
rlabel metal2 31080 36904 31080 36904 0 _0922_
rlabel metal2 24136 34496 24136 34496 0 _0923_
rlabel metal2 27384 34160 27384 34160 0 _0924_
rlabel metal2 28280 34216 28280 34216 0 _0925_
rlabel metal2 29288 37800 29288 37800 0 _0926_
rlabel metal2 20776 30632 20776 30632 0 _0927_
rlabel metal2 22904 34272 22904 34272 0 _0928_
rlabel metal2 24696 24360 24696 24360 0 _0929_
rlabel metal2 24584 26236 24584 26236 0 _0930_
rlabel metal2 23240 36792 23240 36792 0 _0931_
rlabel metal3 13440 35672 13440 35672 0 _0932_
rlabel metal2 12824 35560 12824 35560 0 _0933_
rlabel metal3 17304 25872 17304 25872 0 _0934_
rlabel metal2 11200 26488 11200 26488 0 _0935_
rlabel metal2 9408 16856 9408 16856 0 _0936_
rlabel metal2 5320 28672 5320 28672 0 _0937_
rlabel metal2 4760 32704 4760 32704 0 _0938_
rlabel metal2 8232 34160 8232 34160 0 _0939_
rlabel metal2 12096 35672 12096 35672 0 _0940_
rlabel metal2 13160 36120 13160 36120 0 _0941_
rlabel metal2 13384 35280 13384 35280 0 _0942_
rlabel metal2 23128 36232 23128 36232 0 _0943_
rlabel metal2 23800 37464 23800 37464 0 _0944_
rlabel metal2 30968 37352 30968 37352 0 _0945_
rlabel metal2 36344 35896 36344 35896 0 _0946_
rlabel metal2 24584 17248 24584 17248 0 _0947_
rlabel metal2 22456 21336 22456 21336 0 _0948_
rlabel metal2 22792 24024 22792 24024 0 _0949_
rlabel metal2 24472 24360 24472 24360 0 _0950_
rlabel metal2 23576 37184 23576 37184 0 _0951_
rlabel metal2 23912 21504 23912 21504 0 _0952_
rlabel metal2 24024 23296 24024 23296 0 _0953_
rlabel metal2 24808 28728 24808 28728 0 _0954_
rlabel metal2 24248 29792 24248 29792 0 _0955_
rlabel metal2 24024 30352 24024 30352 0 _0956_
rlabel metal2 23912 36736 23912 36736 0 _0957_
rlabel metal2 23688 38864 23688 38864 0 _0958_
rlabel metal2 18480 26712 18480 26712 0 _0959_
rlabel metal3 16296 24472 16296 24472 0 _0960_
rlabel metal2 17192 25536 17192 25536 0 _0961_
rlabel metal2 1512 32088 1512 32088 0 _0962_
rlabel metal2 8232 31416 8232 31416 0 _0963_
rlabel metal2 4816 26040 4816 26040 0 _0964_
rlabel metal2 8904 29624 8904 29624 0 _0965_
rlabel metal4 8456 30856 8456 30856 0 _0966_
rlabel metal2 12824 38920 12824 38920 0 _0967_
rlabel metal3 12432 38920 12432 38920 0 _0968_
rlabel metal3 13440 39592 13440 39592 0 _0969_
rlabel metal2 22344 39032 22344 39032 0 _0970_
rlabel metal2 24640 38920 24640 38920 0 _0971_
rlabel metal3 20440 36232 20440 36232 0 _0972_
rlabel metal3 23072 35896 23072 35896 0 _0973_
rlabel metal3 23408 36456 23408 36456 0 _0974_
rlabel metal2 28952 38668 28952 38668 0 _0975_
rlabel metal2 32536 39256 32536 39256 0 _0976_
rlabel metal2 29624 37968 29624 37968 0 _0977_
rlabel metal2 31528 38248 31528 38248 0 _0978_
rlabel metal3 32536 38696 32536 38696 0 _0979_
rlabel metal3 35896 39368 35896 39368 0 _0980_
rlabel metal3 30632 39480 30632 39480 0 _0981_
rlabel metal2 30184 40208 30184 40208 0 _0982_
rlabel metal3 24136 38584 24136 38584 0 _0983_
rlabel metal3 22568 38808 22568 38808 0 _0984_
rlabel metal3 24136 39032 24136 39032 0 _0985_
rlabel metal2 22680 39256 22680 39256 0 _0986_
rlabel metal2 25032 40040 25032 40040 0 _0987_
rlabel metal2 6552 30184 6552 30184 0 _0988_
rlabel metal3 10192 39032 10192 39032 0 _0989_
rlabel metal2 9912 28280 9912 28280 0 _0990_
rlabel metal2 11032 39200 11032 39200 0 _0991_
rlabel metal2 11256 39536 11256 39536 0 _0992_
rlabel metal2 2856 41888 2856 41888 0 _0993_
rlabel metal3 9912 40152 9912 40152 0 _0994_
rlabel metal3 11480 40488 11480 40488 0 _0995_
rlabel metal3 12264 38808 12264 38808 0 _0996_
rlabel metal2 6888 39536 6888 39536 0 _0997_
rlabel metal2 4984 38752 4984 38752 0 _0998_
rlabel metal2 11872 39480 11872 39480 0 _0999_
rlabel metal2 12376 40040 12376 40040 0 _1000_
rlabel metal2 13160 38864 13160 38864 0 _1001_
rlabel metal3 19656 39256 19656 39256 0 _1002_
rlabel metal2 22008 31976 22008 31976 0 _1003_
rlabel metal2 22904 39648 22904 39648 0 _1004_
rlabel metal2 19768 25872 19768 25872 0 _1005_
rlabel metal2 26264 25816 26264 25816 0 _1006_
rlabel metal3 27496 39480 27496 39480 0 _1007_
rlabel metal2 29064 39984 29064 39984 0 _1008_
rlabel metal2 31192 40712 31192 40712 0 _1009_
rlabel metal2 39480 42448 39480 42448 0 _1010_
rlabel via2 31528 42056 31528 42056 0 _1011_
rlabel metal2 30632 40600 30632 40600 0 _1012_
rlabel metal3 32816 41832 32816 41832 0 _1013_
rlabel metal2 23016 40432 23016 40432 0 _1014_
rlabel metal2 26152 42168 26152 42168 0 _1015_
rlabel metal3 26236 40600 26236 40600 0 _1016_
rlabel metal3 29344 42504 29344 42504 0 _1017_
rlabel metal4 23240 29568 23240 29568 0 _1018_
rlabel metal2 22344 42336 22344 42336 0 _1019_
rlabel metal2 21952 42056 21952 42056 0 _1020_
rlabel metal2 22456 42952 22456 42952 0 _1021_
rlabel metal3 18256 41832 18256 41832 0 _1022_
rlabel metal2 22624 42168 22624 42168 0 _1023_
rlabel metal2 23016 43120 23016 43120 0 _1024_
rlabel metal2 10752 40936 10752 40936 0 _1025_
rlabel metal2 8456 44576 8456 44576 0 _1026_
rlabel metal3 8792 40936 8792 40936 0 _1027_
rlabel metal2 6216 36008 6216 36008 0 _1028_
rlabel metal2 8288 36680 8288 36680 0 _1029_
rlabel metal3 9016 36456 9016 36456 0 _1030_
rlabel metal3 12040 35784 12040 35784 0 _1031_
rlabel metal2 10472 39144 10472 39144 0 _1032_
rlabel metal2 9800 35672 9800 35672 0 _1033_
rlabel metal2 11032 40432 11032 40432 0 _1034_
rlabel metal2 11592 40096 11592 40096 0 _1035_
rlabel metal2 11592 40600 11592 40600 0 _1036_
rlabel metal2 22904 42504 22904 42504 0 _1037_
rlabel metal3 29680 42840 29680 42840 0 _1038_
rlabel metal2 35336 42896 35336 42896 0 _1039_
rlabel metal2 36232 43568 36232 43568 0 _1040_
rlabel metal2 29512 42784 29512 42784 0 _1041_
rlabel metal2 32200 41944 32200 41944 0 _1042_
rlabel metal2 32088 43288 32088 43288 0 _1043_
rlabel metal3 25060 41832 25060 41832 0 _1044_
rlabel metal2 24192 39592 24192 39592 0 _1045_
rlabel metal2 24472 39984 24472 39984 0 _1046_
rlabel metal2 24248 41608 24248 41608 0 _1047_
rlabel metal2 1400 31752 1400 31752 0 _1048_
rlabel metal2 11816 41328 11816 41328 0 _1049_
rlabel metal3 12880 42504 12880 42504 0 _1050_
rlabel metal2 14168 42728 14168 42728 0 _1051_
rlabel metal2 12432 43624 12432 43624 0 _1052_
rlabel metal2 13720 43008 13720 43008 0 _1053_
rlabel metal2 13160 42224 13160 42224 0 _1054_
rlabel metal2 10360 40936 10360 40936 0 _1055_
rlabel metal2 10808 40600 10808 40600 0 _1056_
rlabel metal2 11144 40880 11144 40880 0 _1057_
rlabel metal2 12712 41552 12712 41552 0 _1058_
rlabel metal2 23800 41776 23800 41776 0 _1059_
rlabel metal2 29400 42784 29400 42784 0 _1060_
rlabel metal2 31416 43512 31416 43512 0 _1061_
rlabel metal2 39256 40712 39256 40712 0 _1062_
rlabel metal2 24584 44688 24584 44688 0 _1063_
rlabel metal2 24136 40376 24136 40376 0 _1064_
rlabel metal2 25144 41496 25144 41496 0 _1065_
rlabel metal2 25200 42056 25200 42056 0 _1066_
rlabel metal2 25592 41776 25592 41776 0 _1067_
rlabel metal3 12936 41160 12936 41160 0 _1068_
rlabel metal3 21000 40656 21000 40656 0 _1069_
rlabel metal2 33096 41104 33096 41104 0 _1070_
rlabel metal2 30520 41552 30520 41552 0 _1071_
rlabel metal2 31080 43568 31080 43568 0 _1072_
rlabel metal2 43960 42560 43960 42560 0 _1073_
rlabel metal2 33208 42112 33208 42112 0 _1074_
rlabel metal2 40040 43288 40040 43288 0 _1075_
rlabel metal2 43736 33264 43736 33264 0 _1076_
rlabel metal2 43960 30352 43960 30352 0 _1077_
rlabel metal3 44408 31528 44408 31528 0 _1078_
rlabel metal3 45136 39032 45136 39032 0 _1079_
rlabel metal2 15960 7840 15960 7840 0 _1080_
rlabel metal2 23464 16744 23464 16744 0 _1081_
rlabel metal2 26376 17248 26376 17248 0 _1082_
rlabel metal3 20272 16184 20272 16184 0 _1083_
rlabel metal2 18088 18816 18088 18816 0 _1084_
rlabel metal2 11480 17248 11480 17248 0 _1085_
rlabel metal2 22568 18200 22568 18200 0 _1086_
rlabel metal2 17752 9408 17752 9408 0 _1087_
rlabel metal2 16744 7616 16744 7616 0 _1088_
rlabel metal3 18200 8008 18200 8008 0 _1089_
rlabel metal3 17976 8120 17976 8120 0 _1090_
rlabel metal2 29456 17528 29456 17528 0 _1091_
rlabel metal2 23352 18816 23352 18816 0 _1092_
rlabel metal2 26600 14056 26600 14056 0 _1093_
rlabel metal2 20272 9576 20272 9576 0 _1094_
rlabel metal2 6384 16296 6384 16296 0 _1095_
rlabel metal2 15624 5320 15624 5320 0 _1096_
rlabel metal2 22568 25564 22568 25564 0 _1097_
rlabel metal2 23352 7672 23352 7672 0 _1098_
rlabel metal2 23016 7336 23016 7336 0 _1099_
rlabel metal3 16576 5880 16576 5880 0 _1100_
rlabel metal2 12600 15848 12600 15848 0 _1101_
rlabel metal2 18648 6496 18648 6496 0 _1102_
rlabel metal2 16744 6328 16744 6328 0 _1103_
rlabel metal3 16744 1176 16744 1176 0 _1104_
rlabel metal2 17752 7224 17752 7224 0 _1105_
rlabel metal2 17864 7112 17864 7112 0 _1106_
rlabel metal3 29848 8008 29848 8008 0 _1107_
rlabel metal3 27552 16856 27552 16856 0 _1108_
rlabel metal3 34496 15512 34496 15512 0 _1109_
rlabel metal2 26712 15652 26712 15652 0 _1110_
rlabel metal2 26600 7784 26600 7784 0 _1111_
rlabel metal2 27496 8344 27496 8344 0 _1112_
rlabel metal3 28672 7672 28672 7672 0 _1113_
rlabel metal2 27720 5936 27720 5936 0 _1114_
rlabel metal2 31416 8960 31416 8960 0 _1115_
rlabel metal2 29344 5208 29344 5208 0 _1116_
rlabel metal2 27496 6832 27496 6832 0 _1117_
rlabel metal3 32760 11592 32760 11592 0 _1118_
rlabel metal2 23800 13160 23800 13160 0 _1119_
rlabel metal2 27720 16128 27720 16128 0 _1120_
rlabel metal2 30632 9688 30632 9688 0 _1121_
rlabel metal2 32200 15792 32200 15792 0 _1122_
rlabel metal3 31584 12264 31584 12264 0 _1123_
rlabel metal2 30072 9800 30072 9800 0 _1124_
rlabel metal3 31584 9128 31584 9128 0 _1125_
rlabel metal3 18424 34104 18424 34104 0 _1126_
rlabel metal2 18760 34048 18760 34048 0 _1127_
rlabel metal2 32200 15400 32200 15400 0 _1128_
rlabel metal2 33432 26264 33432 26264 0 _1129_
rlabel metal2 42728 23744 42728 23744 0 _1130_
rlabel metal2 39704 24192 39704 24192 0 _1131_
rlabel metal2 23128 12320 23128 12320 0 _1132_
rlabel metal2 33768 25368 33768 25368 0 _1133_
rlabel metal2 33544 25200 33544 25200 0 _1134_
rlabel metal3 34328 24584 34328 24584 0 _1135_
rlabel metal2 34328 24976 34328 24976 0 _1136_
rlabel metal4 26264 28728 26264 28728 0 _1137_
rlabel metal2 26376 28280 26376 28280 0 _1138_
rlabel metal2 26488 27384 26488 27384 0 _1139_
rlabel metal2 41608 24584 41608 24584 0 _1140_
rlabel metal3 18480 2408 18480 2408 0 _1141_
rlabel metal2 21616 39480 21616 39480 0 _1142_
rlabel metal2 25928 30184 25928 30184 0 _1143_
rlabel metal2 25760 29624 25760 29624 0 _1144_
rlabel metal2 22512 32536 22512 32536 0 _1145_
rlabel metal2 21672 33936 21672 33936 0 _1146_
rlabel metal2 22680 32480 22680 32480 0 _1147_
rlabel metal2 21336 33040 21336 33040 0 _1148_
rlabel metal2 21672 31136 21672 31136 0 _1149_
rlabel metal2 19320 32424 19320 32424 0 _1150_
rlabel metal2 19656 33320 19656 33320 0 _1151_
rlabel metal4 17976 30016 17976 30016 0 _1152_
rlabel metal2 19432 35532 19432 35532 0 _1153_
rlabel metal3 19656 34104 19656 34104 0 _1154_
rlabel metal3 19432 36456 19432 36456 0 _1155_
rlabel metal2 19208 35616 19208 35616 0 _1156_
rlabel metal2 18312 40824 18312 40824 0 _1157_
rlabel metal2 18760 35728 18760 35728 0 _1158_
rlabel metal2 21336 36624 21336 36624 0 _1159_
rlabel metal2 20664 36456 20664 36456 0 _1160_
rlabel metal2 21896 38780 21896 38780 0 _1161_
rlabel metal2 21672 37688 21672 37688 0 _1162_
rlabel metal2 21560 38696 21560 38696 0 _1163_
rlabel metal2 21560 38920 21560 38920 0 _1164_
rlabel metal3 21504 40376 21504 40376 0 _1165_
rlabel metal2 21784 40208 21784 40208 0 _1166_
rlabel metal2 20664 40152 20664 40152 0 _1167_
rlabel metal2 21952 39592 21952 39592 0 _1168_
rlabel metal3 19488 41944 19488 41944 0 _1169_
rlabel metal2 21224 42672 21224 42672 0 _1170_
rlabel metal3 15960 38920 15960 38920 0 _1171_
rlabel metal2 19208 41776 19208 41776 0 _1172_
rlabel metal2 17976 42224 17976 42224 0 _1173_
rlabel metal2 19040 41384 19040 41384 0 _1174_
rlabel metal2 18088 41104 18088 41104 0 _1175_
rlabel metal2 15624 39144 15624 39144 0 _1176_
rlabel metal2 17304 40600 17304 40600 0 _1177_
rlabel metal2 17696 39032 17696 39032 0 _1178_
rlabel metal2 8904 32172 8904 32172 0 _1179_
rlabel metal2 9912 30856 9912 30856 0 _1180_
rlabel metal2 11144 34384 11144 34384 0 _1181_
rlabel metal3 11592 32760 11592 32760 0 _1182_
rlabel metal3 10584 33992 10584 33992 0 _1183_
rlabel metal3 9240 34104 9240 34104 0 _1184_
rlabel metal2 15176 34160 15176 34160 0 _1185_
rlabel metal2 14224 36232 14224 36232 0 _1186_
rlabel metal2 14168 36848 14168 36848 0 _1187_
rlabel metal2 14840 34272 14840 34272 0 _1188_
rlabel metal2 15680 34216 15680 34216 0 _1189_
rlabel metal3 16968 34888 16968 34888 0 _1190_
rlabel metal2 15960 36120 15960 36120 0 _1191_
rlabel metal2 16520 37968 16520 37968 0 _1192_
rlabel metal2 16296 37632 16296 37632 0 _1193_
rlabel metal2 14616 38416 14616 38416 0 _1194_
rlabel metal2 15624 38024 15624 38024 0 _1195_
rlabel metal2 10584 38808 10584 38808 0 _1196_
rlabel metal2 11928 37128 11928 37128 0 _1197_
rlabel metal3 12264 36456 12264 36456 0 _1198_
rlabel metal2 10360 38416 10360 38416 0 _1199_
rlabel metal2 10584 37128 10584 37128 0 _1200_
rlabel metal2 6216 37128 6216 37128 0 _1201_
rlabel metal3 4928 37240 4928 37240 0 _1202_
rlabel metal3 2408 31472 2408 31472 0 _1203_
rlabel metal2 6328 37352 6328 37352 0 _1204_
rlabel metal2 4200 36232 4200 36232 0 _1205_
rlabel metal2 3976 38024 3976 38024 0 _1206_
rlabel metal2 3864 39648 3864 39648 0 _1207_
rlabel metal2 2296 40432 2296 40432 0 _1208_
rlabel metal2 2856 40544 2856 40544 0 _1209_
rlabel metal2 40040 24136 40040 24136 0 _1210_
rlabel metal2 15848 40544 15848 40544 0 _1211_
rlabel metal2 4648 39256 4648 39256 0 _1212_
rlabel metal2 4312 39592 4312 39592 0 _1213_
rlabel metal2 3920 41048 3920 41048 0 _1214_
rlabel metal2 4256 41048 4256 41048 0 _1215_
rlabel metal3 3584 42840 3584 42840 0 _1216_
rlabel metal2 4872 42840 4872 42840 0 _1217_
rlabel metal3 3304 44072 3304 44072 0 _1218_
rlabel metal2 5768 44296 5768 44296 0 _1219_
rlabel metal2 3248 44184 3248 44184 0 _1220_
rlabel metal2 3416 44408 3416 44408 0 _1221_
rlabel metal2 5600 42728 5600 42728 0 _1222_
rlabel metal2 6048 42728 6048 42728 0 _1223_
rlabel metal2 15736 43120 15736 43120 0 _1224_
rlabel metal2 16128 41384 16128 41384 0 _1225_
rlabel metal3 15064 43624 15064 43624 0 _1226_
rlabel metal2 20776 5824 20776 5824 0 _1227_
rlabel metal2 3192 16464 3192 16464 0 _1228_
rlabel metal3 15624 43400 15624 43400 0 _1229_
rlabel metal2 2520 30128 2520 30128 0 _1230_
rlabel metal2 2072 29624 2072 29624 0 _1231_
rlabel metal2 3640 29736 3640 29736 0 _1232_
rlabel metal2 3864 29232 3864 29232 0 _1233_
rlabel metal2 3752 29792 3752 29792 0 _1234_
rlabel metal2 2744 29400 2744 29400 0 _1235_
rlabel metal2 2296 32312 2296 32312 0 _1236_
rlabel metal2 3192 31808 3192 31808 0 _1237_
rlabel metal2 8008 36848 8008 36848 0 _1238_
rlabel metal4 2632 31864 2632 31864 0 _1239_
rlabel metal2 3640 32144 3640 32144 0 _1240_
rlabel metal2 3024 31976 3024 31976 0 _1241_
rlabel metal2 4984 32088 4984 32088 0 _1242_
rlabel metal2 5992 31640 5992 31640 0 _1243_
rlabel metal2 5096 32536 5096 32536 0 _1244_
rlabel metal2 5768 33320 5768 33320 0 _1245_
rlabel metal2 3248 33208 3248 33208 0 _1246_
rlabel metal3 5264 34104 5264 34104 0 _1247_
rlabel metal2 2912 33096 2912 33096 0 _1248_
rlabel metal2 3136 33432 3136 33432 0 _1249_
rlabel metal2 6888 34608 6888 34608 0 _1250_
rlabel metal2 6328 34888 6328 34888 0 _1251_
rlabel via2 6552 35896 6552 35896 0 _1252_
rlabel metal3 6720 35784 6720 35784 0 _1253_
rlabel metal2 7560 35952 7560 35952 0 _1254_
rlabel metal2 5880 36960 5880 36960 0 _1255_
rlabel metal2 7336 36904 7336 36904 0 _1256_
rlabel metal3 6776 38472 6776 38472 0 _1257_
rlabel metal2 6328 38808 6328 38808 0 _1258_
rlabel metal2 20104 16912 20104 16912 0 clknet_0_wb_clk_i
rlabel metal2 2856 6832 2856 6832 0 clknet_4_0_0_wb_clk_i
rlabel metal2 40768 17528 40768 17528 0 clknet_4_10_0_wb_clk_i
rlabel metal3 40544 16856 40544 16856 0 clknet_4_11_0_wb_clk_i
rlabel metal3 39368 33432 39368 33432 0 clknet_4_12_0_wb_clk_i
rlabel metal2 29456 41944 29456 41944 0 clknet_4_13_0_wb_clk_i
rlabel metal3 40544 24696 40544 24696 0 clknet_4_14_0_wb_clk_i
rlabel metal2 22904 41328 22904 41328 0 clknet_4_15_0_wb_clk_i
rlabel metal3 2296 18424 2296 18424 0 clknet_4_1_0_wb_clk_i
rlabel metal2 24584 11368 24584 11368 0 clknet_4_2_0_wb_clk_i
rlabel metal2 20776 18368 20776 18368 0 clknet_4_3_0_wb_clk_i
rlabel metal2 1904 39592 1904 39592 0 clknet_4_4_0_wb_clk_i
rlabel metal2 1736 34384 1736 34384 0 clknet_4_5_0_wb_clk_i
rlabel metal2 19432 38920 19432 38920 0 clknet_4_6_0_wb_clk_i
rlabel metal2 22344 40880 22344 40880 0 clknet_4_7_0_wb_clk_i
rlabel metal3 35784 16856 35784 16856 0 clknet_4_8_0_wb_clk_i
rlabel metal2 38472 16912 38472 16912 0 clknet_4_9_0_wb_clk_i
rlabel metal3 47208 42112 47208 42112 0 custom_settings[0]
rlabel metal3 44408 42616 44408 42616 0 custom_settings[1]
rlabel metal3 48762 2744 48762 2744 0 io_in_1[0]
rlabel metal2 48216 7616 48216 7616 0 io_in_1[1]
rlabel metal2 48216 12656 48216 12656 0 io_in_1[2]
rlabel metal3 46592 18424 46592 18424 0 io_in_1[3]
rlabel metal2 48104 21224 48104 21224 0 io_in_1[4]
rlabel metal2 48216 27608 48216 27608 0 io_in_1[5]
rlabel metal2 48104 32032 48104 32032 0 io_in_1[6]
rlabel metal2 43904 25592 43904 25592 0 io_in_1[7]
rlabel metal2 1848 42112 1848 42112 0 io_in_2
rlabel metal2 19320 47698 19320 47698 0 io_out[10]
rlabel metal2 20888 47698 20888 47698 0 io_out[11]
rlabel metal3 23856 46088 23856 46088 0 io_out[12]
rlabel metal2 30296 47642 30296 47642 0 io_out[17]
rlabel metal2 31864 46914 31864 46914 0 io_out[18]
rlabel metal2 33432 47698 33432 47698 0 io_out[19]
rlabel metal2 35000 46354 35000 46354 0 io_out[20]
rlabel metal3 36904 44520 36904 44520 0 io_out[21]
rlabel metal2 40376 46032 40376 46032 0 io_out[22]
rlabel metal2 39704 47810 39704 47810 0 io_out[23]
rlabel metal2 41272 47698 41272 47698 0 io_out[24]
rlabel metal2 42840 48034 42840 48034 0 io_out[25]
rlabel metal2 44408 47642 44408 47642 0 io_out[26]
rlabel metal2 45976 46466 45976 46466 0 io_out[27]
rlabel metal3 15792 44520 15792 44520 0 io_out[8]
rlabel metal2 17752 47642 17752 47642 0 io_out[9]
rlabel metal3 45472 23128 45472 23128 0 net1
rlabel metal3 24360 15568 24360 15568 0 net10
rlabel metal2 2240 42728 2240 42728 0 net11
rlabel metal3 2296 16968 2296 16968 0 net12
rlabel metal2 19656 45136 19656 45136 0 net13
rlabel metal2 20776 45416 20776 45416 0 net14
rlabel metal2 45304 45136 45304 45136 0 net15
rlabel metal3 23016 44016 23016 44016 0 net16
rlabel metal2 32424 44352 32424 44352 0 net17
rlabel metal2 35112 45920 35112 45920 0 net18
rlabel metal2 35224 37800 35224 37800 0 net19
rlabel metal2 47992 24360 47992 24360 0 net2
rlabel metal2 39032 39928 39032 39928 0 net20
rlabel metal2 41608 39760 41608 39760 0 net21
rlabel metal2 43232 42056 43232 42056 0 net22
rlabel metal2 43960 44800 43960 44800 0 net23
rlabel metal2 40040 44576 40040 44576 0 net24
rlabel metal2 42840 40376 42840 40376 0 net25
rlabel metal2 45640 39984 45640 39984 0 net26
rlabel metal2 16072 45136 16072 45136 0 net27
rlabel metal2 16856 44744 16856 44744 0 net28
rlabel metal2 3752 45752 3752 45752 0 net29
rlabel metal2 18648 7896 18648 7896 0 net3
rlabel metal2 5544 46592 5544 46592 0 net30
rlabel metal2 6888 45752 6888 45752 0 net31
rlabel metal2 8568 46368 8568 46368 0 net32
rlabel metal2 10024 45752 10024 45752 0 net33
rlabel metal2 11592 45752 11592 45752 0 net34
rlabel metal2 12600 46648 12600 46648 0 net35
rlabel metal2 14616 47530 14616 47530 0 net36
rlabel metal2 23464 44184 23464 44184 0 net37
rlabel metal2 26712 47320 26712 47320 0 net38
rlabel metal2 27496 46592 27496 46592 0 net39
rlabel metal2 47936 7672 47936 7672 0 net4
rlabel metal2 28728 47530 28728 47530 0 net40
rlabel metal3 19544 24920 19544 24920 0 net41
rlabel metal2 47768 44632 47768 44632 0 net42
rlabel metal2 33544 42280 33544 42280 0 net43
rlabel metal2 20216 23856 20216 23856 0 net44
rlabel metal2 11872 20104 11872 20104 0 net45
rlabel metal2 12040 27384 12040 27384 0 net46
rlabel metal2 33656 29680 33656 29680 0 net47
rlabel metal2 10248 28784 10248 28784 0 net48
rlabel metal2 26712 31584 26712 31584 0 net49
rlabel metal3 45472 12824 45472 12824 0 net5
rlabel metal2 16464 32312 16464 32312 0 net50
rlabel metal2 10248 25872 10248 25872 0 net51
rlabel metal2 15792 35784 15792 35784 0 net52
rlabel metal2 34216 36064 34216 36064 0 net53
rlabel metal3 41160 37408 41160 37408 0 net54
rlabel metal2 31976 43456 31976 43456 0 net55
rlabel metal3 39704 36568 39704 36568 0 net56
rlabel metal3 33320 36456 33320 36456 0 net57
rlabel metal2 14504 31024 14504 31024 0 net58
rlabel metal3 10192 29512 10192 29512 0 net59
rlabel metal2 47880 18144 47880 18144 0 net6
rlabel metal2 15400 21056 15400 21056 0 net60
rlabel metal2 10024 18256 10024 18256 0 net61
rlabel metal2 26712 16912 26712 16912 0 net7
rlabel metal2 26040 17416 26040 17416 0 net8
rlabel metal2 23968 15512 23968 15512 0 net9
rlabel metal2 1680 17080 1680 17080 0 rst_n
rlabel metal2 11256 19656 11256 19656 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[0\]
rlabel metal3 17976 20216 17976 20216 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[1\]
rlabel metal2 15792 21560 15792 21560 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[2\]
rlabel metal2 2184 25032 2184 25032 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\]
rlabel metal2 8624 18424 8624 18424 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.in
rlabel metal3 2128 21448 2128 21448 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[0\]
rlabel metal2 6552 17528 6552 17528 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[1\]
rlabel metal2 8232 21616 8232 21616 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\]
rlabel metal3 2352 19320 2352 19320 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[3\]
rlabel metal2 2408 22848 2408 22848 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.in
rlabel metal2 19768 22400 19768 22400 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[0\]
rlabel metal3 19544 22344 19544 22344 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[1\]
rlabel metal2 21448 18704 21448 18704 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[2\]
rlabel metal2 15680 20888 15680 20888 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[3\]
rlabel metal2 23072 24696 23072 24696 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.in
rlabel metal2 28224 18312 28224 18312 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[0\]
rlabel metal3 22400 20776 22400 20776 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[1\]
rlabel metal2 25424 20776 25424 20776 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[2\]
rlabel metal2 23576 20020 23576 20020 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\]
rlabel metal2 40264 19600 40264 19600 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.in
rlabel metal2 45640 25928 45640 25928 0 tt_um_rejunity_sn76489.clk_counter\[0\]
rlabel metal2 46200 26320 46200 26320 0 tt_um_rejunity_sn76489.clk_counter\[1\]
rlabel metal2 46872 25928 46872 25928 0 tt_um_rejunity_sn76489.clk_counter\[2\]
rlabel metal2 47544 25480 47544 25480 0 tt_um_rejunity_sn76489.clk_counter\[3\]
rlabel metal2 45192 24640 45192 24640 0 tt_um_rejunity_sn76489.clk_counter\[4\]
rlabel metal2 45528 21896 45528 21896 0 tt_um_rejunity_sn76489.clk_counter\[5\]
rlabel metal2 43848 22904 43848 22904 0 tt_um_rejunity_sn76489.clk_counter\[6\]
rlabel metal2 32984 18144 32984 18144 0 tt_um_rejunity_sn76489.control_noise\[0\]\[0\]
rlabel metal2 31864 20216 31864 20216 0 tt_um_rejunity_sn76489.control_noise\[0\]\[1\]
rlabel metal2 36680 18704 36680 18704 0 tt_um_rejunity_sn76489.control_noise\[0\]\[2\]
rlabel metal2 13496 7952 13496 7952 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[0\]
rlabel metal2 17752 5824 17752 5824 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[1\]
rlabel metal2 16632 5544 16632 5544 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[2\]
rlabel metal3 16436 6440 16436 6440 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[3\]
rlabel metal2 6720 10472 6720 10472 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[4\]
rlabel metal4 7000 9296 7000 9296 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[5\]
rlabel metal2 6328 13552 6328 13552 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[6\]
rlabel metal2 5992 11984 5992 11984 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[7\]
rlabel metal2 9912 13104 9912 13104 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[8\]
rlabel metal2 9016 16744 9016 16744 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[9\]
rlabel metal2 30968 7504 30968 7504 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[0\]
rlabel metal3 29512 6104 29512 6104 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[1\]
rlabel metal3 30520 4984 30520 4984 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[2\]
rlabel metal2 27048 6384 27048 6384 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[3\]
rlabel metal2 16576 10584 16576 10584 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[4\]
rlabel metal2 18536 9352 18536 9352 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[5\]
rlabel metal2 20552 11200 20552 11200 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[6\]
rlabel metal3 18928 11704 18928 11704 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[7\]
rlabel metal3 19768 13048 19768 13048 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[8\]
rlabel metal2 20776 14280 20776 14280 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[9\]
rlabel metal2 41048 10976 41048 10976 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[0\]
rlabel metal2 32088 10248 32088 10248 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[1\]
rlabel metal2 40152 9520 40152 9520 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[2\]
rlabel metal2 38920 9240 38920 9240 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[3\]
rlabel metal2 31416 15148 31416 15148 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[4\]
rlabel metal2 27832 9968 27832 9968 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[5\]
rlabel metal2 30184 10416 30184 10416 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[6\]
rlabel metal2 32088 12768 32088 12768 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[7\]
rlabel metal2 26600 12824 26600 12824 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[8\]
rlabel metal2 26488 14672 26488 14672 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[9\]
rlabel metal2 2184 26236 2184 26236 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[0\]
rlabel metal2 1848 31416 1848 31416 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[1\]
rlabel metal4 3416 31416 3416 31416 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[2\]
rlabel metal2 5880 32704 5880 32704 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[3\]
rlabel metal2 4368 33432 4368 33432 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[4\]
rlabel metal3 5376 36344 5376 36344 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[5\]
rlabel metal2 7000 39648 7000 39648 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[6\]
rlabel metal2 7168 42504 7168 42504 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[7\]
rlabel metal2 7448 44576 7448 44576 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[8\]
rlabel metal2 12600 43792 12600 43792 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[9\]
rlabel metal3 10360 33320 10360 33320 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[0\]
rlabel metal2 10024 33656 10024 33656 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[1\]
rlabel metal2 15400 34104 15400 34104 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[2\]
rlabel metal2 14728 37408 14728 37408 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[3\]
rlabel metal3 15176 38752 15176 38752 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[4\]
rlabel metal2 4536 37128 4536 37128 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[5\]
rlabel metal2 4872 38864 4872 38864 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[6\]
rlabel metal2 3136 42616 3136 42616 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[7\]
rlabel metal3 5488 44408 5488 44408 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[8\]
rlabel metal2 15512 43120 15512 43120 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[9\]
rlabel metal2 33432 27888 33432 27888 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[0\]
rlabel metal2 33096 24696 33096 24696 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[1\]
rlabel metal2 26264 28280 26264 28280 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[2\]
rlabel metal2 23128 34328 23128 34328 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[3\]
rlabel metal2 20776 31528 20776 31528 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[4\]
rlabel metal2 20440 36512 20440 36512 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[5\]
rlabel metal2 20328 37744 20328 37744 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[6\]
rlabel metal2 22232 39648 22232 39648 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[7\]
rlabel via2 20328 42728 20328 42728 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[8\]
rlabel metal2 16856 39704 16856 39704 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[9\]
rlabel metal2 37016 24360 37016 24360 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[0\]
rlabel metal2 39592 26628 39592 26628 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[1\]
rlabel metal2 34776 29792 34776 29792 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[2\]
rlabel metal2 33544 31808 33544 31808 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[3\]
rlabel metal2 34888 34104 34888 34104 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[4\]
rlabel metal2 26264 36120 26264 36120 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[5\]
rlabel metal2 26040 38248 26040 38248 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[6\]
rlabel metal2 26712 41944 26712 41944 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[7\]
rlabel metal2 26712 43680 26712 43680 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[8\]
rlabel metal2 24304 44296 24304 44296 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[9\]
rlabel metal2 10976 16744 10976 16744 0 tt_um_rejunity_sn76489.latch_control_reg\[0\]
rlabel metal3 14784 15512 14784 15512 0 tt_um_rejunity_sn76489.latch_control_reg\[1\]
rlabel metal2 16968 19936 16968 19936 0 tt_um_rejunity_sn76489.latch_control_reg\[2\]
rlabel metal2 41160 13048 41160 13048 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[0\]
rlabel metal2 39816 13384 39816 13384 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[1\]
rlabel metal2 39368 16408 39368 16408 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[2\]
rlabel metal2 38080 18648 38080 18648 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[3\]
rlabel metal3 36680 20776 36680 20776 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[4\]
rlabel metal2 37912 20608 37912 20608 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[5\]
rlabel metal2 39256 21224 39256 21224 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[6\]
rlabel metal2 48160 15512 48160 15512 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[10\]
rlabel metal2 47880 20132 47880 20132 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[11\]
rlabel metal2 46760 19824 46760 19824 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[12\]
rlabel metal2 46424 17080 46424 17080 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[13\]
rlabel metal2 43736 16352 43736 16352 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[14\]
rlabel metal2 39032 18480 39032 18480 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[1\]
rlabel metal2 44016 7672 44016 7672 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[2\]
rlabel metal3 46088 4984 46088 4984 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[3\]
rlabel metal3 46928 6440 46928 6440 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[4\]
rlabel metal2 47432 8008 47432 8008 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[5\]
rlabel metal2 47432 9296 47432 9296 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[6\]
rlabel metal3 45696 11256 45696 11256 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[7\]
rlabel metal3 47096 12040 47096 12040 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[8\]
rlabel metal2 47824 13944 47824 13944 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[9\]
rlabel metal2 41832 15456 41832 15456 0 tt_um_rejunity_sn76489.noise\[0\].gen.restart_noise
rlabel metal2 44632 19600 44632 19600 0 tt_um_rejunity_sn76489.noise\[0\].gen.signal_edge.previous_signal_state_0
rlabel metal2 39872 30296 39872 30296 0 tt_um_rejunity_sn76489.pwm.accumulator\[0\]
rlabel metal2 43848 41552 43848 41552 0 tt_um_rejunity_sn76489.pwm.accumulator\[10\]
rlabel metal2 45304 43120 45304 43120 0 tt_um_rejunity_sn76489.pwm.accumulator\[11\]
rlabel metal2 41384 29120 41384 29120 0 tt_um_rejunity_sn76489.pwm.accumulator\[1\]
rlabel metal3 39032 31864 39032 31864 0 tt_um_rejunity_sn76489.pwm.accumulator\[2\]
rlabel metal2 38696 33768 38696 33768 0 tt_um_rejunity_sn76489.pwm.accumulator\[3\]
rlabel metal2 35672 36176 35672 36176 0 tt_um_rejunity_sn76489.pwm.accumulator\[4\]
rlabel metal2 36008 37240 36008 37240 0 tt_um_rejunity_sn76489.pwm.accumulator\[5\]
rlabel metal2 37464 39704 37464 39704 0 tt_um_rejunity_sn76489.pwm.accumulator\[6\]
rlabel metal2 36512 39592 36512 39592 0 tt_um_rejunity_sn76489.pwm.accumulator\[7\]
rlabel metal2 34720 43624 34720 43624 0 tt_um_rejunity_sn76489.pwm.accumulator\[8\]
rlabel metal2 39368 44856 39368 44856 0 tt_um_rejunity_sn76489.pwm.accumulator\[9\]
rlabel metal2 44072 35168 44072 35168 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[0\]
rlabel metal3 45304 30184 45304 30184 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[1\]
rlabel metal2 47320 29288 47320 29288 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[2\]
rlabel metal2 47208 34552 47208 34552 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[3\]
rlabel metal2 46816 33544 46816 33544 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[4\]
rlabel metal2 41384 34048 41384 34048 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[0\]
rlabel metal2 45304 38612 45304 38612 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[10\]
rlabel metal2 45752 35616 45752 35616 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[11\]
rlabel metal2 41496 35504 41496 35504 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[1\]
rlabel metal2 42728 34776 42728 34776 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[2\]
rlabel metal2 41944 37184 41944 37184 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[3\]
rlabel metal3 43792 38136 43792 38136 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[4\]
rlabel metal2 44184 39032 44184 39032 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[5\]
rlabel metal2 42728 40824 42728 40824 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[6\]
rlabel metal2 39928 42000 39928 42000 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[7\]
rlabel metal2 41496 40656 41496 40656 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[8\]
rlabel metal2 43904 39592 43904 39592 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[9\]
rlabel metal2 12040 8288 12040 8288 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[0\]
rlabel metal2 11312 6888 11312 6888 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[1\]
rlabel metal2 11480 6328 11480 6328 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[2\]
rlabel metal2 9016 5040 9016 5040 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[3\]
rlabel metal2 6776 6720 6776 6720 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[4\]
rlabel metal3 8680 8232 8680 8232 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[5\]
rlabel metal2 8008 8848 8008 8848 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[6\]
rlabel metal2 9800 10248 9800 10248 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[7\]
rlabel metal3 13216 12152 13216 12152 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[8\]
rlabel metal2 8288 16184 8288 16184 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[9\]
rlabel metal2 32200 7392 32200 7392 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[0\]
rlabel metal3 30632 5936 30632 5936 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[1\]
rlabel metal2 33432 5264 33432 5264 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[2\]
rlabel metal2 25536 5096 25536 5096 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[3\]
rlabel metal2 23128 4648 23128 4648 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[4\]
rlabel metal3 20944 6664 20944 6664 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[5\]
rlabel metal2 21448 8960 21448 8960 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[6\]
rlabel metal2 22120 10416 22120 10416 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[7\]
rlabel metal2 24696 11928 24696 11928 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[8\]
rlabel metal2 22288 13832 22288 13832 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[9\]
rlabel metal2 41776 10584 41776 10584 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[0\]
rlabel metal2 42000 8232 42000 8232 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[1\]
rlabel metal2 40880 7448 40880 7448 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[2\]
rlabel metal2 39144 9184 39144 9184 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[3\]
rlabel metal2 39032 5992 39032 5992 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[4\]
rlabel metal2 38864 3640 38864 3640 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[5\]
rlabel metal4 36344 5432 36344 5432 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[6\]
rlabel metal2 35784 11704 35784 11704 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[7\]
rlabel metal2 39704 12712 39704 12712 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[8\]
rlabel metal2 39480 13328 39480 13328 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[9\]
rlabel metal3 14672 3304 14672 3304 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
