magic
tech gf180mcuD
magscale 1 10
timestamp 1702458819
<< nwell >>
rect 1258 41120 44662 41984
rect 1258 40391 3773 40416
rect 1258 39577 44662 40391
rect 1258 39552 18221 39577
rect 1258 38823 2653 38848
rect 1258 38009 44662 38823
rect 1258 37984 10300 38009
rect 1258 37255 20909 37280
rect 1258 36416 44662 37255
rect 1258 35687 2653 35712
rect 1258 34873 44662 35687
rect 1258 34848 30989 34873
rect 1258 34119 5005 34144
rect 1258 33280 44662 34119
rect 1258 32551 20797 32576
rect 1258 31737 44662 32551
rect 1258 31712 2989 31737
rect 1258 30983 6909 31008
rect 1258 30169 44662 30983
rect 1258 30144 11432 30169
rect 1258 29415 2653 29440
rect 1258 28576 44662 29415
rect 1258 27847 21624 27872
rect 1258 27033 44662 27847
rect 1258 27008 41853 27033
rect 1258 25465 44662 26304
rect 1258 25440 39566 25465
rect 1258 24711 36253 24736
rect 1258 23897 44662 24711
rect 1258 23872 18351 23897
rect 1258 23143 13182 23168
rect 1258 22329 44662 23143
rect 1258 22304 2653 22329
rect 1258 21575 14030 21600
rect 1258 20736 44662 21575
rect 1258 20007 3213 20032
rect 1258 19193 44662 20007
rect 1258 19168 23709 19193
rect 1258 18439 20616 18464
rect 1258 17625 44662 18439
rect 1258 17600 41741 17625
rect 1258 16871 4445 16896
rect 1258 16057 44662 16871
rect 1258 16032 2653 16057
rect 1258 15303 27784 15328
rect 1258 14464 44662 15303
rect 1258 13735 41853 13760
rect 1258 12896 44662 13735
rect 1258 12167 4221 12192
rect 1258 11353 44662 12167
rect 1258 11328 2653 11353
rect 1258 10599 30429 10624
rect 1258 9785 44662 10599
rect 1258 9760 26509 9785
rect 1258 9031 35805 9056
rect 1258 8217 44662 9031
rect 1258 8192 7512 8217
rect 1258 6649 44662 7488
rect 1258 6624 11544 6649
rect 1258 5895 26061 5920
rect 1258 5081 44662 5895
rect 1258 5056 16541 5081
rect 1258 4327 14301 4352
rect 1258 3488 44662 4327
<< pwell >>
rect 1258 41984 44662 42422
rect 1258 40416 44662 41120
rect 1258 38848 44662 39552
rect 1258 37280 44662 37984
rect 1258 35712 44662 36416
rect 1258 34144 44662 34848
rect 1258 32576 44662 33280
rect 1258 31008 44662 31712
rect 1258 29440 44662 30144
rect 1258 27872 44662 28576
rect 1258 26304 44662 27008
rect 1258 24736 44662 25440
rect 1258 23168 44662 23872
rect 1258 21600 44662 22304
rect 1258 20032 44662 20736
rect 1258 18464 44662 19168
rect 1258 16896 44662 17600
rect 1258 15328 44662 16032
rect 1258 13760 44662 14464
rect 1258 12192 44662 12896
rect 1258 10624 44662 11328
rect 1258 9056 44662 9760
rect 1258 7488 44662 8192
rect 1258 5920 44662 6624
rect 1258 4352 44662 5056
rect 1258 3050 44662 3488
<< obsm1 >>
rect 1344 3076 44576 42396
<< metal2 >>
rect 1792 45200 1904 46000
rect 5600 45200 5712 46000
rect 9408 45200 9520 46000
rect 13216 45200 13328 46000
rect 17024 45200 17136 46000
rect 20832 45200 20944 46000
rect 24640 45200 24752 46000
rect 28448 45200 28560 46000
rect 32256 45200 32368 46000
rect 36064 45200 36176 46000
rect 39872 45200 39984 46000
rect 43680 45200 43792 46000
<< obsm2 >>
rect 1964 45140 5540 45332
rect 5772 45140 9348 45332
rect 9580 45140 13156 45332
rect 13388 45140 16964 45332
rect 17196 45140 20772 45332
rect 21004 45140 24580 45332
rect 24812 45140 28388 45332
rect 28620 45140 32196 45332
rect 32428 45140 36004 45332
rect 36236 45140 39812 45332
rect 40044 45140 43620 45332
rect 43852 45140 44100 45332
rect 1820 3098 44100 45140
<< obsm3 >>
rect 1922 3108 44110 42364
<< metal4 >>
rect 4448 3076 4768 42396
rect 19808 3076 20128 42396
rect 35168 3076 35488 42396
<< obsm4 >>
rect 15372 8978 15876 10846
<< labels >>
rlabel metal2 s 9408 45200 9520 46000 6 io_in
port 1 nsew signal input
rlabel metal2 s 13216 45200 13328 46000 6 io_out[0]
port 2 nsew signal output
rlabel metal2 s 17024 45200 17136 46000 6 io_out[1]
port 3 nsew signal output
rlabel metal2 s 20832 45200 20944 46000 6 io_out[2]
port 4 nsew signal output
rlabel metal2 s 24640 45200 24752 46000 6 io_out[3]
port 5 nsew signal output
rlabel metal2 s 28448 45200 28560 46000 6 io_out[4]
port 6 nsew signal output
rlabel metal2 s 32256 45200 32368 46000 6 io_out[5]
port 7 nsew signal output
rlabel metal2 s 36064 45200 36176 46000 6 io_out[6]
port 8 nsew signal output
rlabel metal2 s 39872 45200 39984 46000 6 io_out[7]
port 9 nsew signal output
rlabel metal2 s 43680 45200 43792 46000 6 io_out[8]
port 10 nsew signal output
rlabel metal2 s 5600 45200 5712 46000 6 rst_n
port 11 nsew signal input
rlabel metal4 s 4448 3076 4768 42396 6 vdd
port 12 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 42396 6 vdd
port 12 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 42396 6 vss
port 13 nsew ground bidirectional
rlabel metal2 s 1792 45200 1904 46000 6 wb_clk_i
port 14 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 46000 46000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1002460
string GDS_FILE /media/lucah/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1-multi/openlane/diceroll/runs/23_12_13_10_10/results/signoff/diceroll.magic.gds
string GDS_START 240128
<< end >>

