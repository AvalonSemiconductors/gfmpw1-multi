* NGSPICE file created from wrapped_qcpu.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
.ends

.subckt wrapped_qcpu custom_settings[0] custom_settings[10] custom_settings[11] custom_settings[12]
+ custom_settings[13] custom_settings[14] custom_settings[15] custom_settings[16]
+ custom_settings[17] custom_settings[18] custom_settings[19] custom_settings[1] custom_settings[20]
+ custom_settings[21] custom_settings[22] custom_settings[23] custom_settings[24]
+ custom_settings[25] custom_settings[26] custom_settings[27] custom_settings[28]
+ custom_settings[29] custom_settings[2] custom_settings[30] custom_settings[31] custom_settings[3]
+ custom_settings[4] custom_settings[5] custom_settings[6] custom_settings[7] custom_settings[8]
+ custom_settings[9] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15]
+ io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23]
+ io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31]
+ io_in[32] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0]
+ io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17]
+ io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0]
+ io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17]
+ io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[24] io_out[25]
+ io_out[27] io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] rst_n sram_addr[0] sram_addr[1]
+ sram_addr[2] sram_addr[3] sram_addr[4] sram_addr[5] sram_gwe sram_in[0] sram_in[1]
+ sram_in[2] sram_in[3] sram_in[4] sram_in[5] sram_in[6] sram_in[7] sram_out[0] sram_out[1]
+ sram_out[2] sram_out[3] sram_out[4] sram_out[5] sram_out[6] sram_out[7] vdd vss
+ wb_clk_i io_oeb[22] io_out[26] io_out[23]
XFILLER_0_94_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05903_ cpu.timer_div\[1\] _01407_ _01182_ _01408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09671_ _04686_ _04681_ _04698_ _04699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06883_ cpu.PC\[4\] _02381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07534__A1 cpu.regs\[11\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08622_ _02772_ _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06888__A3 _02385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05834_ _01339_ _01340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08553_ _03727_ _03735_ _00336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05765_ _01269_ _01270_ _01271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_77_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08484_ _03672_ _00330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07504_ _02916_ _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07435_ _02867_ _02868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05696_ _01201_ _01202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_81_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07366_ _02791_ _02804_ _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09105_ _04150_ _04160_ _04161_ _00462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06317_ cpu.timer_div\[5\] _01184_ _01818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07297_ _02748_ _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_102_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09036_ _00591_ _02561_ _04102_ _04109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06248_ _01657_ _01659_ _01749_ _01750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_79_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09062__I1 _03090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06179_ _01161_ net92 _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_92_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09938_ cpu.PORTA_DDR\[7\] _04899_ _04908_ _04904_ _04909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_5_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09869_ _04846_ _04858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07525__A1 cpu.regs\[12\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09278__A1 _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output37_I net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_104_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10575_ _00513_ clknet_leaf_70_wb_clk_i cpu.ROM_spi_cycle\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06264__B2 _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06264__A1 _01465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10060__A2 _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05311__I0 cpu.regs\[8\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08005__A2 _03288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06016__A1 _01054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07764__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_60_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_60_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10009_ _04718_ _02040_ _02043_ _04973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_64_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05550_ cpu.IO_addr_buff\[4\] _01056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05451__I _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05481_ _00769_ _00989_ _00990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_46_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07220_ cpu.timer_capture\[1\] _02674_ _02686_ _02687_ _02688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_73_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07151_ _02613_ _02622_ _02627_ _02628_ _00041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08244__A2 _03451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09441__A1 _02418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06255__A1 _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06102_ cpu.br_rel_dest\[3\] _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_89_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07082_ _02569_ _00031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09807__B net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06033_ _01498_ _01173_ _01535_ _01536_ _01259_ _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_2_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07984_ _03280_ _00222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09723_ _00662_ _04740_ _04722_ _04741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06935_ _02363_ _02365_ _02421_ _02431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05081__I2 cpu.regs\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09654_ _04685_ _00487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06866_ _02090_ _02095_ _02364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_38_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08605_ _03768_ _03770_ _00353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05817_ _00950_ _01323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_96_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09585_ _04596_ _04618_ _00690_ _00485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06797_ _02288_ _00994_ _02295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05748_ _01253_ _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08536_ _03695_ _03696_ _03714_ _03721_ _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_38_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05679_ _01184_ _01185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08467_ _02772_ _03660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07418_ _02840_ cpu.uart.receive_div_counter\[15\] _02846_ _02847_ _02850_ _02851_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_08398_ _03609_ _03610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08672__I _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06494__A1 _00646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07349_ _02786_ _02327_ _02789_ _02790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_115_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10360_ _00299_ clknet_leaf_55_wb_clk_i cpu.orig_IO_addr_buff\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10291_ _00230_ clknet_leaf_44_wb_clk_i cpu.uart.dout\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09019_ _04095_ _00802_ _04096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09499__A1 _04209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05221__A2 _00756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07349__I1 _02327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06485__A1 cpu.toggle_top\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07198__I _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09423__A1 _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10627_ _00565_ clknet_leaf_0_wb_clk_i cpu.regs\[15\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10558_ _00496_ clknet_leaf_74_wb_clk_i cpu.startup_cycle\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10489_ _00427_ clknet_leaf_49_wb_clk_i cpu.uart.divisor\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_59_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06004__A4 _01243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05446__I _00955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06720_ _02216_ _02217_ _02179_ _02218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_06651_ _02145_ _02146_ _02149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_91_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05602_ _01107_ _01105_ _01108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_115_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09370_ _02562_ _04409_ _04410_ _04411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06582_ _00637_ _00955_ _02080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08321_ _03548_ _03549_ _03550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05533_ _01036_ _01037_ _01038_ _01039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08252_ cpu.uart.receive_buff\[1\] _03494_ _03498_ cpu.uart.receive_buff\[0\] _03499_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05464_ _00973_ _00974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07203_ _02672_ _00049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_55_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08183_ _03343_ _03439_ _03442_ _03443_ _03444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_54_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05395_ _00007_ _00907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07134_ _02615_ _02601_ _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10024__A2 _02721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07065_ _02547_ _02549_ _02553_ _02542_ _02554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_112_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06016_ _01054_ _01199_ _01518_ _01519_ _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_76_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09178__B1 _02721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07967_ _03229_ _03223_ _00788_ _03269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09706_ _02450_ _04727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06918_ _02169_ _02357_ _02415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07898_ _03195_ cpu.spi.div_counter\[4\] _03210_ _03214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_97_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09637_ cpu.last_addr\[0\] cpu.ROM_addr_buff\[0\] _04669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_69_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06849_ _02204_ _02233_ _02347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_87_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09568_ _02375_ _00925_ _04601_ _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08519_ _03702_ _03703_ _03704_ _03705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06467__A1 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08456__A2 _03574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09499_ _04209_ _04524_ _04535_ _04326_ _04536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_41_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10412_ _00351_ clknet_leaf_104_wb_clk_i cpu.pwm_counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10343_ _00282_ clknet_leaf_36_wb_clk_i cpu.uart.receive_div_counter\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07746__I cpu.PC\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09169__B1 _02109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10274_ _00213_ clknet_leaf_60_wb_clk_i cpu.spi.data_out_buff\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09182__B _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_14_Left_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_83_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08998__A3 _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_104_Right_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_83_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05180_ cpu.base_address\[3\] _00717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05969__B1 _01466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_23_Left_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08870_ _03354_ _03975_ _00413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07821_ cpu.timer\[11\] _03142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07752_ _03081_ _03082_ _02074_ _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07683_ cpu.regs\[4\]\[1\] _03029_ _03031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06703_ _02177_ _02199_ _02200_ _02201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_32_Left_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_94_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09422_ _02380_ _02783_ _02560_ _04461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06634_ _02126_ _02127_ _02132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_35_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09353_ _00763_ _04394_ _04395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08304_ _03535_ _03536_ _00286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_4_5_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06449__A1 _01910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06565_ _01365_ _01156_ _01349_ _02063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_118_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09284_ _04324_ _04297_ _04325_ _04327_ _04328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05516_ _01022_ _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_06496_ _01994_ _01995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08235_ cpu.uart.data_buff\[8\] _03458_ _03486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05447_ _00956_ _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08166_ _03378_ _03430_ _03431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05378_ cpu.regs\[8\]\[0\] cpu.regs\[9\]\[0\] cpu.regs\[10\]\[0\] cpu.regs\[11\]\[0\]
+ _00888_ _00889_ _00890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_43_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_41_Left_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07117_ _02601_ _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08097_ _03372_ _03374_ cpu.uart.div_counter\[1\] _03375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07048_ _02049_ _02051_ _02537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_100_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05188__A1 _00723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08999_ cpu.IO_addr_buff\[7\] _04066_ _04080_ _04069_ _04081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08397__I _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05035__S1 _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06688__B2 _00891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08346__B _03570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10326_ _00265_ clknet_leaf_53_wb_clk_i cpu.uart.data_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06612__A1 _02109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10257_ _00196_ clknet_leaf_48_wb_clk_i cpu.spi.dout\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10188_ _00127_ clknet_leaf_121_wb_clk_i cpu.regs\[10\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09865__A1 _04014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06350_ _01739_ _00987_ _01851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06281_ _01326_ _01773_ _01777_ _01332_ _01782_ _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_05301_ _00832_ net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08020_ cpu.uart.receive_buff\[7\] _03307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08770__I _03121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05232_ _00764_ _00767_ _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05163_ _00700_ _00701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08199__A4 _03456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09971_ _04933_ _04922_ _04937_ _03347_ _00552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_110_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05094_ _00618_ _00634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08922_ _04000_ _04015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08853_ cpu.spi.divisor\[3\] _03960_ _03964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06906__A2 _02401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05996_ cpu.spi.busy _01100_ _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07804_ cpu.timer_div_counter\[1\] _03125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08784_ cpu.timer\[14\] _03908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05634__I _01127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05590__A1 _00675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07735_ _02551_ _02348_ _03067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09550__B _00776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09405_ _02571_ _04317_ _04445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07666_ _02990_ _03016_ _03020_ _00164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06617_ _00588_ _00984_ _02115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07597_ cpu.regs\[8\]\[3\] _02969_ _02975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06548_ _00666_ _00667_ _02046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_75_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09336_ _02530_ _04352_ _04377_ _04378_ _04195_ _04379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_23_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09267_ _04299_ _04296_ _04308_ _04310_ _04311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_08218_ _00947_ _03455_ _03472_ _03473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06479_ cpu.timer_capture\[7\] _01182_ _01975_ _01977_ _01242_ _01978_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_50_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09198_ _00707_ _01133_ _04210_ _04244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_31_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08149_ cpu.uart.div_counter\[10\] _03370_ _03416_ _03417_ _03418_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07296__I _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10111_ _00054_ clknet_leaf_29_wb_clk_i cpu.timer_capture\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output67_I net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10042_ _05003_ _05004_ _05005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08898__A2 _03995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_10_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08855__I _03958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_85_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_85_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_54_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_14_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_14_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_112_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10309_ _00248_ clknet_leaf_38_wb_clk_i cpu.uart.div_counter\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05850_ _01355_ _01356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_89_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07520_ _01875_ cpu.regs\[12\]\[5\] _02916_ _02928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05781_ cpu.regs\[4\]\[7\] cpu.regs\[5\]\[7\] cpu.regs\[6\]\[7\] cpu.regs\[7\]\[7\]
+ _00961_ _01286_ _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_clkbuf_leaf_99_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07451_ _02870_ _02881_ _02882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_88_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06402_ _01171_ _01900_ _01901_ _01902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_45_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07382_ _02819_ _02108_ _02789_ _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09121_ _04166_ _04171_ _04172_ _00467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_45_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06333_ _01769_ _01772_ _01834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09052_ _02378_ _04095_ _04120_ _04121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06264_ _01465_ _01759_ _01765_ _01461_ _01766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_114_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08003_ cpu.uart.dout\[2\] _03294_ _03295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05215_ cpu.uart.busy cpu.spi.busy _00723_ _00751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_13_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06195_ net29 _01697_ _01599_ _01698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05146_ _00684_ _00012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06052__A2 _00944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09954_ _04921_ _04922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05077_ _00576_ _00618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09885_ _04846_ _04870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08905_ _04000_ _04002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_57_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05792__C _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08836_ cpu.timer_capture\[14\] _03941_ _03951_ _03939_ _03952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_79_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08767_ cpu.timer\[11\] _03894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_56_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05979_ _01331_ _01484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07718_ _00787_ _02596_ _00692_ _03050_ _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
X_08698_ _03835_ _03836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_0_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07649_ _01873_ _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_94_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05866__A2 _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09319_ _04358_ _04351_ _00776_ _04362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10591_ _00529_ clknet_leaf_66_wb_clk_i net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_106_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_97_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05618__A2 _01087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput42 net42 io_oeb[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput64 net64 io_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput75 net75 io_out[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05475__S _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput53 net53 io_oeb[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput97 net97 sram_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput86 net86 sram_addr[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_37_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10025_ _01469_ _04987_ _04988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_106_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06282__A2 _01548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06951_ _02440_ _02445_ _02446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09670_ _04695_ _04697_ _04698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05902_ _01406_ _01407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08621_ _03658_ _03779_ _03782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06882_ cpu.PC\[6\] _02380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_6_Left_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05833_ _01324_ _01338_ _01339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08552_ _03707_ _03733_ _03735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05764_ _01040_ _01270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07298__A1 _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08483_ cpu.toggle_top\[5\] _03666_ _03670_ _03671_ _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07503_ _02889_ _02915_ _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07434_ _02845_ _02864_ _02866_ _02867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05695_ _01200_ _01201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_81_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07365_ _02333_ _02329_ _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_94_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06316_ _01803_ _01610_ _01815_ _01816_ _01184_ _01817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_09104_ cpu.last_addr\[6\] _04157_ _04161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07296_ _02748_ _02749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09035_ _04108_ _00445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06247_ _01656_ _01749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06178_ _01574_ _01577_ _01681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05129_ _00666_ _00667_ _00668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_92_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09937_ _04837_ _04900_ _04908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_5_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09868_ _04018_ _04854_ _04857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07525__A2 _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08819_ _03142_ _03928_ _03929_ _03937_ _03938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09799_ _04796_ _03758_ _03763_ _04801_ _04802_ _04803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_68_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10574_ _00512_ clknet_leaf_73_wb_clk_i cpu.ROM_spi_cycle\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07461__A1 _02071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06016__A2 _01199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07213__A1 cpu.timer_capture\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_79_Left_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05775__A1 _01279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07516__A2 _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10008_ _04930_ _02481_ _04971_ _04972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_19_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05480_ _00988_ _00989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_104_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07150_ _02617_ _02628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_54_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06255__A2 net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07081_ _02361_ _02568_ _02544_ _02569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06101_ _01167_ _01603_ _01604_ _00015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06032_ cpu.pwm_top\[2\] _01254_ _01172_ _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06007__A2 _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09722_ _02451_ _02462_ _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07983_ cpu.spi.data_in_buff\[5\] _03277_ _03278_ cpu.spi.data_in_buff\[4\] _03280_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07327__C _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08704__A1 cpu.timer_capture\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06934_ _02414_ _02420_ _02430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09653_ _04640_ _04643_ _04682_ _04684_ _04685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06865_ _02360_ _02362_ _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_38_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09584_ _04346_ _04613_ _04617_ _04618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08604_ _03769_ _03767_ _03770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05816_ _01315_ _01319_ _01321_ _01322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_118_Right_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08535_ _03688_ _03692_ _03716_ _03720_ _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__06191__A1 _01484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06796_ _02273_ _02293_ _02294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__05642__I _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05747_ _01252_ _01253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07997__C _02628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05678_ _01183_ _01184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_64_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08953__I _04032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08466_ _03658_ _03655_ _03659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07417_ cpu.uart.receive_div_counter\[5\] _01804_ _02848_ _02849_ _02850_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_92_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08397_ _00688_ _03609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06494__A2 _01294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07348_ _02788_ _02789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09432__A2 _04028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07279_ _02644_ _02729_ _02734_ _02737_ _00060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_5_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10290_ _00229_ clknet_4_13_0_wb_clk_i cpu.uart.dout\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09018_ _00702_ _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_60_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08943__A1 _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06182__B2 _01462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06182__A1 _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05368__S0 _00878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10626_ _00564_ clknet_leaf_118_wb_clk_i cpu.regs\[15\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07434__A1 _02845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10557_ _00495_ clknet_leaf_74_wb_clk_i cpu.startup_cycle\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05296__I0 cpu.regs\[8\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10488_ _00426_ clknet_leaf_41_wb_clk_i cpu.uart.divisor\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05996__A1 cpu.spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_87_Left_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07737__A2 _03065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08103__I _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_12_0_wb_clk_i clknet_0_wb_clk_i clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_06650_ _00821_ _01955_ _02148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05601_ _01044_ _01047_ _01107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_86_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06581_ _02078_ _01996_ _02079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08320_ _03543_ _03544_ _02862_ _03549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_96_Left_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05532_ _01028_ _00759_ _01038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_24_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08251_ _03497_ _03498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05463_ _00972_ _00973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_117_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07202_ cpu.uart.divisor\[7\] _02651_ _02671_ _02662_ _02672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_74_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08182_ _03339_ _03368_ _03443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_55_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05394_ cpu.regs\[4\]\[1\] cpu.regs\[5\]\[1\] cpu.regs\[6\]\[1\] cpu.regs\[7\]\[1\]
+ _00899_ _00902_ _00906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_07133_ _02614_ _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_70_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07064_ _02534_ _02337_ _02550_ _02552_ _02553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06015_ net8 _01517_ _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09178__A1 _01022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07728__A2 _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05739__A1 cpu.timer_capture\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07966_ _03268_ _00216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09705_ _04726_ _00497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input29_I sram_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06917_ _02413_ _02414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07897_ _03195_ _03210_ cpu.spi.div_counter\[4\] _03213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09636_ cpu.last_addr\[3\] cpu.ROM_addr_buff\[3\] _04667_ _04668_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_65_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06848_ _02284_ _02344_ _02345_ _02346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_87_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05911__A1 cpu.timer_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09567_ _04600_ _04582_ _04576_ _04601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06779_ _02269_ _02270_ _02277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09498_ cpu.orig_PC\[9\] _04033_ _04535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08683__I _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08518_ cpu.toggle_ctr\[3\] _01608_ _01498_ cpu.toggle_ctr\[2\] _03704_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_108_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08449_ _02393_ _03633_ _03647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10411_ _00350_ clknet_leaf_105_wb_clk_i cpu.pwm_counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10342_ _00281_ clknet_leaf_38_wb_clk_i cpu.uart.receive_div_counter\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output97_I net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07967__A2 _03223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09169__A1 _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10273_ _00212_ clknet_leaf_60_wb_clk_i cpu.spi.data_out_buff\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07719__A2 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_39_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_39_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_49_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09644__A2 cpu.ROM_addr_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10609_ _00547_ clknet_leaf_60_wb_clk_i cpu.PORTA_DDR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_40_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07937__I _02660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05969__A1 _01462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07820_ cpu.timer\[12\] _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__05197__A2 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07751_ net19 _03064_ _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06702_ _02197_ _02198_ _02200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05192__I _00728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07682_ _02980_ _03028_ _03030_ _00170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09421_ _04459_ _04460_ _04381_ _00479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06633_ _02081_ _02130_ _02131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06564_ _00687_ _02047_ _02061_ _02062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_09352_ _01704_ _04314_ _04393_ _04321_ _04394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_47_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08303_ cpu.uart.receive_div_counter\[6\] _03531_ _03529_ _03536_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06449__A2 _01948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05515_ _01021_ _01022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09283_ _04326_ _04327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06495_ _01292_ _01289_ _00913_ _01994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08234_ _03485_ _00267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05446_ _00955_ _00956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_27_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08165_ cpu.uart.div_counter\[14\] _03426_ _03427_ _03430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09548__B _04440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05377_ _00873_ _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08071__A1 _03347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07116_ _02596_ _02599_ _02600_ _02511_ _02601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_15_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08096_ _03369_ _03374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05504__S0 _00871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07047_ cpu.rom_data_dist _02536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_100_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09571__A1 _00771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06385__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08998_ _01953_ _04029_ _04040_ _04079_ _04059_ _04080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__07582__I _02965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07949_ _03233_ _03255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_46_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06198__I _01700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09619_ _04162_ _04650_ _04651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_66_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_26_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10325_ _00264_ clknet_leaf_54_wb_clk_i cpu.uart.data_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06612__A2 _01294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10256_ _00195_ clknet_leaf_49_wb_clk_i cpu.spi.dout\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07693__S _03026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09562__A1 _02393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08365__A2 _03581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10187_ _00126_ clknet_leaf_125_wb_clk_i cpu.regs\[10\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_89_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06280_ _01780_ _01781_ _01782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05300_ _00831_ _00832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_115_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05231_ _00766_ _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05162_ net71 _00700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09970_ _02460_ _04936_ _04922_ _04937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_73_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05093_ _00617_ _00633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_110_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08921_ _01005_ _04014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10026__C _04196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08852_ _02644_ _03959_ _03963_ _00407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07803_ cpu.timer_div\[3\] cpu.timer_div_counter\[3\] _03124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06367__B2 _01331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08783_ _03843_ _03906_ _03907_ _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05995_ cpu.timer_capture\[10\] _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_07734_ _02259_ _02346_ _02347_ _03066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07665_ cpu.regs\[5\]\[2\] _03017_ _03020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09404_ _04313_ _04444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06616_ _02098_ _02113_ _02114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_109_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07596_ _02923_ _02970_ _02974_ _00140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06547_ _02044_ _02045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09335_ _04338_ _04378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_23_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06478_ _01976_ _01407_ _01633_ _01977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08961__I _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09266_ _04309_ _04310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08217_ cpu.uart.data_buff\[4\] _03464_ _03472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05429_ _00870_ _00939_ _00940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_90_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10275__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09197_ _04233_ _04238_ _04242_ _00759_ _04243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_7_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07577__I _02965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08148_ _03318_ _03411_ _03417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08079_ _03354_ _03359_ _00237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10110_ _00053_ clknet_leaf_22_wb_clk_i cpu.timer_capture\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09544__A1 cpu.PC\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_123_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10041_ _01675_ _04987_ _05004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_59_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_6_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06530__A1 net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08871__I _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_54_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_54_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10308_ _00247_ clknet_leaf_38_wb_clk_i cpu.uart.div_counter\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_60_Left_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09207__I _04252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10239_ _00178_ clknet_leaf_107_wb_clk_i cpu.regs\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_83_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05780_ _00874_ _01286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07450_ _02823_ cpu.uart.receive_counter\[1\] _02876_ _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__06521__A1 _01466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06521__B2 _01484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06401_ cpu.pwm_top\[6\] _01178_ _01901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07381_ _01699_ _02780_ _02818_ _02819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09120_ cpu.last_addr\[11\] _04142_ _04172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06332_ _01306_ _01832_ _01833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09051_ _00702_ cpu.regs\[3\]\[0\] _04120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08002_ _03286_ _03294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_103_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06263_ _01762_ _01764_ _01765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08026__B2 _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08026__A1 _02853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05214_ _00749_ _00722_ _00660_ _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_4_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06194_ _01549_ _01654_ _01696_ _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_114_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05145_ _00683_ _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08730__B _03529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09953_ _02499_ _00696_ _02489_ _02505_ _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_05076_ _00572_ _00617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09884_ _04819_ _04866_ _04869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08904_ _04000_ _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_99_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08835_ _03920_ _03950_ _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08766_ _01499_ _03841_ _03893_ _03616_ _00391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09561__B _00690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input11_I io_in[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07717_ _02055_ _02470_ _02597_ _03050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_79_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05978_ _01310_ _01319_ _01318_ _01483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08697_ _03366_ _01058_ _02727_ _03835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_0_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07648_ _03008_ _00158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07579_ _01495_ _02966_ _00131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07068__A2 _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09318_ _02811_ _02614_ _04360_ _04361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_36_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10590_ _00528_ clknet_leaf_67_wb_clk_i net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_63_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09249_ _04292_ _04293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09065__I0 cpu.regs\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput43 net43 io_oeb[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput65 net65 io_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput54 net54 io_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput76 net76 io_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput87 net87 sram_addr[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_37_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10024_ _04986_ _02721_ _02011_ _04987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08866__I _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_101_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_101_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_85_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05490__A1 _00992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09508__A1 _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06950_ _02031_ _02073_ _02443_ _02444_ _02070_ _02445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA_input3_I io_in[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05901_ _01077_ _00650_ _01115_ _01079_ _01406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__05465__I _00974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06881_ cpu.PC\[7\] _02379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08620_ _03781_ _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05832_ _00718_ _00950_ _01338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07680__I _03026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08551_ _03732_ _03733_ _03734_ _00335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_11_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05763_ cpu.C _01269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05694_ _01196_ _01199_ _01200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08482_ _02772_ _03671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07502_ _01130_ _01135_ _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_07433_ cpu.uart.receiving _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_81_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_77_Right_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09103_ _04114_ _04159_ _04160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_61_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07364_ _02802_ _02796_ _02803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06315_ cpu.spi.divisor\[5\] _01097_ _01610_ _01816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_60_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07295_ _01204_ _02747_ _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_45_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09034_ _04107_ cpu.ROM_addr_buff\[3\] _04104_ _04108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06246_ _01741_ _01747_ _01748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_107_Left_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_103_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05481__A1 _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06177_ _01663_ _01680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05128_ cpu.ROM_spi_cycle\[4\] cpu.ROM_spi_cycle\[0\] _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_92_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_86_Right_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09936_ _04907_ _00547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_5_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05059_ _00575_ _00601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07076__B _02563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05375__I _00877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09867_ _04856_ _00529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_116_Left_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09798_ cpu.pwm_top\[6\] cpu.pwm_counter\[6\] _04802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08818_ _00998_ _03930_ _03937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07590__I _02968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08749_ _02720_ _03871_ _03879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08486__A1 cpu.toggle_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_95_Right_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_83_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_101_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09310__I _04033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10573_ _00511_ clknet_leaf_69_wb_clk_i cpu.ROM_spi_cycle\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10045__A1 _01299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07461__A2 _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05311__I2 cpu.regs\[10\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09185__C _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10007_ _04929_ _04969_ _04970_ _04971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05378__I2 cpu.regs\[10\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_67_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07080_ _01874_ _02566_ _02567_ _02568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06100_ cpu.regs\[9\]\[2\] _01375_ _01604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06031_ cpu.timer_top\[10\] _01175_ _01532_ _01534_ _01179_ _01535_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_112_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_78_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07982_ _03279_ _00221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05215__A1 cpu.uart.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09721_ _04738_ _04716_ _04739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05195__I _00700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06933_ _02428_ _02421_ _02422_ _02410_ _02429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_09652_ _04683_ _04684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_38_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06864_ _02361_ _01997_ _02359_ _02362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06715__A1 _00820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09583_ _04333_ _04599_ _04616_ _04541_ _04403_ _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08603_ cpu.pwm_counter\[4\] _03769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06795_ _00801_ _02083_ _02293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05815_ _01315_ _01320_ _01321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05746_ _01124_ _01252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08534_ _03682_ _03678_ _03719_ _03686_ _03720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_49_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05677_ _01073_ _01098_ _01045_ _01080_ _01183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__08455__B _03646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08465_ _00921_ _03658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07416_ cpu.uart.receive_div_counter\[2\] _02849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_92_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08396_ cpu.orig_flags\[2\] _03607_ _03608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07347_ _02037_ _02077_ _02541_ _02787_ _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__10027__A1 _04292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07278_ _02736_ _02737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09017_ _04094_ _00441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_33_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06229_ _01643_ _01729_ _01730_ _01731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_41_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09919_ _04823_ _04889_ _04895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output42_I net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05065__S0 _00600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08459__A1 _01052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05368__S1 _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10018__A1 _01269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10018__B2 _02721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10625_ _00563_ clknet_leaf_121_wb_clk_i cpu.regs\[15\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07434__A2 _02864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10556_ _00494_ clknet_leaf_72_wb_clk_i cpu.startup_cycle\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10487_ _00425_ clknet_leaf_50_wb_clk_i cpu.uart.divisor\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_75_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06945__A1 cpu.regs\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05600_ _01104_ _01105_ _01106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06173__A2 _00956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06580_ _00836_ _02078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_86_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05531_ _00754_ _01037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08250_ _02872_ _03496_ _03497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08870__A1 _03354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05462_ _00960_ _00966_ _00971_ _00972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_07201_ _02670_ _02654_ _02671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08181_ _03345_ _03440_ _03442_ _00257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_62_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_9_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_9_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_54_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05393_ _00006_ _00905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_07132_ _01139_ _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07063_ net1 _02037_ _02551_ _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06014_ _01506_ _01053_ _01513_ _01516_ _01517_ _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_100_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07728__A3 _02401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07965_ cpu.spi.data_out_buff\[7\] _03255_ _03267_ _03258_ _03268_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09704_ _02456_ _04722_ _04725_ _04684_ _04726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06916_ _02355_ _02358_ _02360_ _02413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07896_ _03203_ _03212_ _00202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09635_ cpu.last_addr\[2\] _04647_ _04667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06847_ _02235_ _02258_ _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05911__A2 _01175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09566_ _04577_ _04600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06778_ _02269_ _02270_ _02276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05729_ _01081_ _01235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08517_ cpu.toggle_ctr\[2\] _01498_ _01419_ cpu.toggle_ctr\[1\] _03703_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_09497_ _04370_ _04533_ _04534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08861__A1 cpu.spi.divisor\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08448_ _03644_ _03645_ _03646_ _00320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_13_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08379_ _03595_ _03596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10410_ _00349_ clknet_leaf_16_wb_clk_i cpu.pwm_counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10341_ _00280_ clknet_leaf_37_wb_clk_i cpu.uart.receive_div_counter\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10272_ _00211_ clknet_leaf_62_wb_clk_i cpu.spi.data_out_buff\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09169__A2 _02261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07719__A3 _02072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_79_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_79_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_79_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_69_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08852__A1 _02644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10608_ _00546_ clknet_leaf_60_wb_clk_i cpu.PORTA_DDR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_51_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10539_ _00477_ clknet_leaf_93_wb_clk_i cpu.PC\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07750_ _03075_ _03080_ _03064_ _03081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06701_ _02197_ _02198_ _02199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07681_ cpu.regs\[4\]\[0\] _03029_ _03030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09420_ _02586_ _04262_ _04460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06632_ _00638_ _00996_ _02129_ _02130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_35_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09096__A1 cpu.ROM_addr_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06563_ cpu.rom_data_dist _02060_ _02061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09351_ _04316_ _04383_ _04392_ _04319_ _04393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_19_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08302_ cpu.uart.receive_div_counter\[6\] _03525_ _03534_ _03520_ _03535_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09282_ _00761_ _04326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05514_ _00895_ _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08233_ cpu.uart.data_buff\[6\] _03475_ _03484_ _03462_ _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06494_ _00646_ _01294_ _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_35_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05445_ _00954_ _00955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08164_ _03425_ _03429_ _00253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05376_ _00887_ _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_08095_ _00793_ _03373_ _00240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07115_ _00696_ _02599_ _02600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_30_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07046_ _00787_ _02535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_42_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05504__S1 _00900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_113_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09020__A1 _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08997_ cpu.orig_IO_addr_buff\[7\] _04056_ _04057_ _02722_ _04079_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07948_ _03254_ _00212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07709__I0 _03007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05383__I _00894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07879_ _03191_ _03194_ _03198_ _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__07885__A2 _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09618_ cpu.last_addr\[6\] cpu.last_addr\[5\] _04649_ _04650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__09087__A1 cpu.ROM_addr_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09549_ _04578_ _04582_ _04583_ _04584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_126_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_126_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_33_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10324_ _00263_ clknet_leaf_52_wb_clk_i cpu.uart.data_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10255_ _00194_ clknet_leaf_49_wb_clk_i cpu.spi.dout\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10186_ _00125_ clknet_leaf_126_wb_clk_i cpu.regs\[10\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07573__A1 _01114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05887__A1 net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05230_ _00765_ _00766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05161_ _00698_ _00699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05092_ _00632_ net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_110_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08920_ _04000_ _04013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08851_ cpu.spi.divisor\[2\] _03960_ _03963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09553__A2 _04178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07802_ cpu.timer_div\[4\] cpu.timer_div_counter\[4\] _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08782_ cpu.timer_capture\[13\] _03836_ _03761_ _03907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05994_ cpu.toggle_top\[2\] _01498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__06299__I _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07316__A1 cpu.toggle_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07733_ _02376_ _02388_ _03065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07664_ _02988_ _03016_ _03019_ _00163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_84_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09403_ _04299_ _04432_ _04442_ _04310_ _04443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06615_ _02107_ _02112_ _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07595_ cpu.regs\[8\]\[2\] _02971_ _02974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06546_ _02041_ _02043_ _02044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09334_ _02108_ _04334_ _04376_ _04377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_23_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06477_ cpu.timer_div\[7\] _01976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_51_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09265_ _04233_ _04309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08216_ _03471_ _00263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_62_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09196_ _04239_ _04240_ _04241_ _04232_ _04242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_05428_ cpu.regs\[8\]\[2\] cpu.regs\[9\]\[2\] cpu.regs\[10\]\[2\] cpu.regs\[11\]\[2\]
+ _00872_ _00889_ _00939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_15_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08147_ _03404_ _03415_ _03416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05359_ _00004_ _00871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_30_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08078_ _03098_ _03349_ _03358_ _03348_ _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_101_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07029_ _02521_ _02522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10040_ _02022_ _05002_ _01480_ _05003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07555__A1 cpu.regs\[10\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08035__A2 cpu.uart.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05288__I cpu.regs\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07094__I0 _02416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10307_ _00246_ clknet_leaf_40_wb_clk_i cpu.uart.div_counter\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10238_ _00177_ clknet_leaf_116_wb_clk_i cpu.regs\[4\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_23_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_23_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10169_ _00108_ clknet_leaf_3_wb_clk_i cpu.regs\[12\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09299__A1 _02810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06400_ cpu.timer_top\[14\] _01640_ _01252_ _01899_ _01900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_57_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07380_ _02546_ _02817_ _02818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06331_ _00749_ _01148_ _01831_ _01832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09050_ _04119_ _00449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06262_ net94 _01763_ _01764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07678__I _03026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06285__B2 _01786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08001_ cpu.uart.receive_buff\[2\] _03293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05213_ _00748_ _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06193_ _01552_ _01669_ _01686_ _01695_ _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_114_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05144_ _00650_ _00682_ _00683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06037__B2 _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10037__C _04196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09952_ _04713_ _04920_ _00550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05075_ _00616_ net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08903_ _01070_ _01186_ _02632_ _04000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__05260__A2 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09883_ _04868_ _00533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08834_ _03908_ _03922_ _03949_ _03950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08765_ _03148_ _03800_ _03833_ _03892_ _03840_ _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_68_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07716_ _02032_ _03041_ _03049_ _00185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05977_ _01480_ _01481_ _01482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08696_ _03833_ _03834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_0_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07647_ _03007_ cpu.regs\[6\]\[4\] _03000_ _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10242__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07578_ _01374_ _02966_ _00130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_91_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06529_ _01031_ _02027_ _02028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09317_ _04304_ _04359_ _04360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07588__I _02968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09248_ _04249_ _04292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_8_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09065__I1 _02393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09179_ cpu.Z _01120_ _04207_ _04225_ _04226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_50_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06028__A1 _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput66 net66 io_out[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_output72_I net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput55 net55 io_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput44 net44 io_oeb[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput77 net77 io_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput88 net88 sram_addr[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07256__C _02712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07528__A1 _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10023_ _01990_ _04986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_106_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09205__A1 _03456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05490__A2 _00998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05900_ _01383_ _01402_ _01404_ _01185_ _01405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_06880_ _02377_ _02378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05831_ _01299_ _01320_ _01336_ _01337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08550_ cpu.toggle_ctr\[2\] _03730_ _03734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05762_ _01267_ _01268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06577__I _02062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05693_ _01069_ _01067_ _01051_ _01199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_49_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08481_ _02766_ _03667_ _03670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08495__A2 _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07501_ _01373_ _02914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07432_ _00787_ cpu.uart.receiving _02845_ _02864_ _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_81_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09102_ _04137_ _04159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_61_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09444__A1 _02588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07363_ _02383_ _02802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06314_ cpu.uart.dout\[5\] _01194_ _01812_ _01814_ _01101_ _01815_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_73_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07294_ _01056_ _01055_ _02746_ _02747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_09033_ _03623_ _04095_ _04106_ _04107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06245_ _01341_ _01742_ _01746_ _01452_ _01747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_103_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05481__A2 _00989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06176_ _01675_ _01677_ _01678_ _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05127_ cpu.ROM_spi_cycle\[3\] cpu.ROM_spi_cycle\[2\] cpu.ROM_spi_cycle\[1\] _00666_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_40_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09935_ cpu.PORTA_DDR\[6\] _04899_ _04906_ _04904_ _04907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_5_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05058_ _00571_ _00600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09866_ net55 _04853_ _04855_ _04847_ _04856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08817_ _03936_ _00399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07930__A1 _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09797_ cpu.pwm_top\[2\] _04801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08748_ _03878_ _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_95_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08679_ _02644_ _03817_ _03822_ _03820_ _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_83_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10572_ _00510_ clknet_leaf_69_wb_clk_i cpu.ROM_spi_cycle\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08207__I _03450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05311__I3 cpu.regs\[11\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10006_ _04738_ _04707_ _04951_ _04970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07781__I _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05378__I3 cpu.regs\[11\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07021__I _02513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06030_ _01174_ _01533_ _01534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_10_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07981_ cpu.spi.data_in_buff\[4\] _03277_ _03278_ cpu.spi.data_in_buff\[3\] _03279_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05215__A2 cpu.spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06412__A1 _00630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09720_ _02451_ _02453_ _04738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06932_ _02353_ _02366_ _02428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_38_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09651_ _02771_ _04683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_38_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06863_ _00605_ _02361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_89_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08602_ _03552_ _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09582_ _00591_ _04614_ _04615_ _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06794_ _00918_ _02287_ _02291_ _02292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05814_ _00817_ _00894_ _01320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_05745_ cpu.timer_top\[8\] _01175_ _01179_ _01250_ _01251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_08533_ _03717_ cpu.toggle_top\[10\] cpu.toggle_top\[9\] _03718_ _03719_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06479__A1 cpu.timer_capture\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05676_ _01181_ _01182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_77_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08464_ _03657_ _00325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07415_ cpu.uart.divisor\[2\] _02848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08395_ _03595_ _03607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09417__A1 _02416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07346_ _02535_ _02536_ _00693_ _02599_ _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_73_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07277_ _02735_ _02736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09016_ _00992_ _04084_ _04093_ _04089_ _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_5_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06228_ cpu.pwm_top\[4\] _01179_ _01730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_79_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06159_ _01138_ _00860_ _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06403__A1 cpu.toggle_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05386__I _00878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09918_ _04894_ _00542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_69_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09849_ _04815_ _04842_ _04843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05065__S1 _00601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07754__I1 _00837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06010__I _01088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output35_I net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06890__A1 _02378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10624_ _00562_ clknet_leaf_123_wb_clk_i cpu.regs\[15\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10555_ _00493_ clknet_leaf_74_wb_clk_i cpu.startup_cycle\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08381__B _03570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10486_ _00424_ clknet_leaf_40_wb_clk_i cpu.uart.divisor\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06642__A1 _00972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05296__I2 cpu.regs\[10\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_14_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08400__I _03586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05530_ cpu.br_rel_dest\[7\] _01036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__05133__A1 net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05461_ _00967_ _00970_ _00971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08180_ _03441_ _03323_ _03338_ _03442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07200_ _02669_ _02670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_74_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05392_ _00897_ _00903_ _00904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07131_ _02531_ _02613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07062_ _02063_ _02551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_113_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06013_ _01205_ _01517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_103_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10045__C _04904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07964_ _02669_ _03241_ _03266_ _03267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09703_ _04703_ _04711_ _04723_ _04724_ _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_07895_ _03211_ _03210_ _03212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06915_ _02353_ _02366_ _02411_ _02412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09634_ cpu.last_addr\[6\] _04665_ _04666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_65_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06846_ _02302_ _02342_ _02343_ _02344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09638__A1 _04140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09565_ _04598_ _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06777_ _02246_ _02247_ _02275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05372__A1 _00006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05728_ _01233_ _01234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_65_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08516_ cpu.toggle_ctr\[1\] _01419_ _01170_ cpu.toggle_ctr\[0\] _03702_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09496_ _00865_ _04444_ _04532_ _04448_ _04533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08185__C _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08447_ _03609_ _03646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_65_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05659_ _01145_ _01164_ _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_37_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08378_ _03594_ _03577_ _03595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07329_ _02668_ _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_33_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10340_ _00279_ clknet_leaf_43_wb_clk_i cpu.uart.receive_buff\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05278__I2 cpu.regs\[10\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10271_ _00210_ clknet_leaf_63_wb_clk_i cpu.spi.data_out_buff\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06927__A2 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07719__A4 _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_48_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_48_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_83_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10607_ _00545_ clknet_leaf_60_wb_clk_i cpu.PORTA_DDR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_64_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10538_ _00476_ clknet_leaf_99_wb_clk_i cpu.PC\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10469_ _00408_ clknet_leaf_30_wb_clk_i cpu.spi.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_75_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09868__A1 _04018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06700_ _02156_ _02157_ _02144_ _02198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_07680_ _03026_ _03029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07343__A2 _02168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06631_ _02079_ _02080_ _02129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06562_ _02049_ _02051_ _02055_ _02059_ _02060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_87_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_86_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09350_ _02548_ _04317_ _04392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08301_ cpu.uart.receive_div_counter\[6\] _03531_ _03534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09281_ cpu.orig_PC\[2\] _04178_ _04325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05513_ _00868_ _01020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08232_ _02657_ _03476_ _03483_ _03484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06493_ _01770_ _01992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05657__A2 _01158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05444_ _00953_ _00954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_27_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08163_ _03426_ _03374_ _03428_ _03379_ _03429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_55_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05375_ _00877_ _00887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_27_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08094_ _03365_ _03370_ _03372_ _03373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07114_ _02597_ _02598_ _02599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_70_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06606__A1 _00850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07045_ _02036_ _02534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08996_ _04074_ _04078_ _00436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07947_ cpu.spi.data_out_buff\[3\] _03234_ _03253_ _03247_ _03254_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_89_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07709__I1 cpu.regs\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07878_ _03195_ _03187_ _03196_ cpu.spi.divisor\[6\] _03197_ _03198_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_97_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09617_ _04153_ _04648_ _04649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06829_ _02167_ _02327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09548_ _04578_ _04582_ _04440_ _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09479_ _04514_ _04492_ _04516_ _04292_ _04517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_54_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08047__B1 cpu.uart.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08598__A1 _03573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10323_ _00262_ clknet_leaf_52_wb_clk_i cpu.uart.data_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07270__A1 cpu.timer_top\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10254_ _00193_ clknet_leaf_52_wb_clk_i cpu.spi.dout\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10185_ _00124_ clknet_leaf_3_wb_clk_i cpu.regs\[10\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_70_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_109_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09078__A2 _04140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07089__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06836__A1 _02168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05160_ _00693_ _00697_ _00698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_52_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05091_ _00631_ _00632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_0_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08850_ _02732_ _03959_ _03962_ _00406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07801_ _03121_ _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08781_ _03904_ _03811_ _03834_ _03905_ _03906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05993_ _01161_ _01378_ _01380_ _01497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_34_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07732_ _02535_ _02596_ _00692_ _03050_ _03064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_07663_ cpu.regs\[5\]\[1\] _03017_ _03019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05327__A1 _00581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09402_ _04436_ _04439_ _04441_ _04442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06614_ _02110_ _02111_ _02112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09333_ _04375_ _04352_ _04376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07594_ _02921_ _02970_ _02973_ _00139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06545_ _00663_ _02042_ _02043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06476_ _01961_ _01611_ _01973_ _01974_ _01185_ _01975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_75_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09264_ _04302_ _04305_ _04307_ _04308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_118_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08215_ cpu.uart.data_buff\[2\] _03460_ _03470_ _03467_ _03471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_62_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08463__C _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09195_ _01131_ _04239_ _04241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05427_ _00935_ _00937_ _00938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08146_ _03318_ _03411_ _03415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07627__I0 _02943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05358_ _00869_ _00870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08077_ _03098_ _03357_ _03358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05289_ _00820_ _00821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07028_ _02520_ _02521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08979_ _00676_ _04038_ _04064_ _04050_ _04065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_59_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09469__C _04313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10306_ _00245_ clknet_leaf_42_wb_clk_i cpu.uart.div_counter\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_72_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10237_ _00176_ clknet_leaf_114_wb_clk_i cpu.regs\[4\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08743__A1 cpu.timer_capture\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09932__C _04904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10168_ _00107_ clknet_leaf_4_wb_clk_i cpu.regs\[12\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10099_ _00042_ clknet_leaf_40_wb_clk_i cpu.uart.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_63_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_63_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_88_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06330_ _00988_ _01542_ _01791_ _01830_ _01831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06863__I _00605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06809__A1 _00850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06261_ _01760_ _01761_ _01763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06285__A2 _01738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08000_ _03291_ _03288_ _03292_ _02628_ _00226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05212_ _00652_ _00748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05479__I _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09223__A2 _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06192_ _01689_ _01690_ _01692_ _01694_ _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_05143_ _00675_ _00681_ _00682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07234__A1 cpu.timer_capture\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09951_ net75 _04914_ _04919_ _04910_ _04920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08982__B2 _00989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05074_ _00615_ _00616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08902_ _00732_ _03998_ _03999_ _00421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09882_ cpu.PORTB_DDR\[0\] _04865_ _04867_ _04858_ _04868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08833_ _03923_ _02715_ _03949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08764_ _03890_ _03891_ _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05976_ _01442_ _01477_ _01481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_56_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07715_ cpu.regs\[3\]\[7\] _03039_ _03049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08695_ _03832_ _03833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07646_ _01787_ _03007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07577_ _02965_ _02966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_36_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06528_ _01990_ _01549_ _02026_ _02027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_09316_ _04302_ _04303_ _04359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09247_ _04291_ _00474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10537__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06459_ _01038_ _01280_ _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05389__I _00900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09178_ _01022_ _04223_ _01272_ _02721_ _04224_ _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_08129_ _03332_ cpu.uart.div_counter\[6\] _03394_ _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__08973__A1 _01161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput34 net34 io_oeb[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput56 net56 io_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput67 net67 io_out[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_101_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput45 net45 io_oeb[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput78 net78 io_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_output65_I net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput89 net89 sram_gwe vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07528__A2 _02932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06013__I _01205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10022_ _01299_ _00760_ _04984_ _04985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__06200__A2 _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09150__A1 _04196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_113_Right_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08964__B2 _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_9_0_wb_clk_i clknet_0_wb_clk_i clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__05778__B2 _00920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05830_ _01269_ _01320_ _01335_ _01336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_118_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05761_ _01266_ _01267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07500_ _02033_ _02905_ _02913_ _00105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05692_ _01197_ _01198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08480_ _03669_ _00329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07431_ _02855_ _02859_ _02861_ _02863_ _02864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_57_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07362_ _02801_ _00079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_33_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06313_ _00684_ _01813_ _01814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09101_ _04150_ _04156_ _04158_ _00461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_61_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07293_ _01091_ _00766_ _02746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_5_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09032_ _00702_ _00851_ _04106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06244_ _01745_ _01746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06175_ _01658_ _01676_ _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05126_ _00662_ _00663_ _00664_ _00665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__10062__I0 _01788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08313__I cpu.uart.receive_div_counter\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05769__A1 _00658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09934_ _02664_ _04900_ _04906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05057_ _00567_ _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_09865_ _04014_ _04854_ _04855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_5_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08183__A2 _03439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08816_ cpu.timer_capture\[10\] _03919_ _03935_ _03916_ _03936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07930__A2 _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09796_ _04794_ _04795_ _04798_ _04799_ _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_08747_ cpu.timer_capture\[7\] _03843_ _03877_ _03795_ _03878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05959_ _01316_ _01463_ _01464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_95_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08678_ cpu.timer_top\[10\] _03818_ _03822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07629_ _02945_ cpu.regs\[7\]\[6\] _02983_ _02996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_82_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10571_ _00509_ clknet_leaf_70_wb_clk_i cpu.ROM_spi_cycle\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07997__A2 _03288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08946__A1 _04033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_2_Left_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_39_Left_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_112_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10005_ _00663_ _04968_ _04969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_48_Left_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_57_Left_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_78_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07980_ _03271_ _03278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05215__A3 _00723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06412__A2 _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06931_ net19 _02404_ _02427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09650_ _04642_ _04646_ _04681_ _04682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09362__B2 _04378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_66_Left_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08601_ _03573_ _03766_ _03767_ _00352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06862_ _00605_ _01996_ _02359_ _02360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__06176__A1 _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09581_ _04614_ _04599_ _04615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_38_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06793_ _02288_ _00996_ _02290_ _02291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05813_ _01316_ _01318_ _01319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05744_ _01238_ _01245_ _01249_ _01174_ _01250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_54_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08532_ _03680_ _03718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08463_ cpu.toggle_top\[0\] _03654_ _03656_ _02773_ _03657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_49_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07414_ cpu.uart.divisor\[14\] _02847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05675_ _01180_ _01181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_77_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08394_ _00794_ _03598_ _03606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05782__S0 _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07428__A1 _02847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07345_ _01372_ _02780_ _02785_ _02786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07276_ _02535_ _02735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_75_Left_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06227_ cpu.timer_top\[12\] _01414_ _01252_ _01728_ _01729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_61_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09015_ _02531_ _04085_ _04093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06158_ _01605_ _01654_ _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05109_ cpu.IO_addr_buff\[0\] _00648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06089_ _01481_ _01581_ _01593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09917_ cpu.PORTA_DDR\[1\] _04888_ _04892_ _04893_ _04894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09848_ _04840_ _04842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06498__I _01996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09779_ cpu.ROM_spi_cycle\[2\] _04785_ _04787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_96_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10623_ _00561_ clknet_leaf_0_wb_clk_i cpu.regs\[15\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10554_ _00492_ clknet_leaf_71_wb_clk_i cpu.mem_cycle\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10485_ _00423_ clknet_leaf_41_wb_clk_i cpu.uart.divisor\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05296__I3 cpu.regs\[11\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07792__I _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05526__B _01031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08128__I _00792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05460_ _00968_ _00969_ _00897_ _00970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06330__A1 _00988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05391_ cpu.regs\[0\]\[1\] cpu.regs\[1\]\[1\] cpu.regs\[2\]\[1\] cpu.regs\[3\]\[1\]
+ _00899_ _00902_ _00903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_70_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07130_ _02610_ _02603_ _02612_ _02606_ _00036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_27_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07061_ _02335_ _02336_ _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06012_ net61 _01515_ _01053_ _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08798__I _03918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06397__A1 cpu.timer_capture\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07963_ cpu.spi.data_out_buff\[6\] _03231_ _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09702_ _04703_ _02459_ _04716_ _04724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_07894_ _03195_ _03211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06914_ _02363_ _02365_ _02411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06149__A1 _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09633_ cpu.last_addr\[5\] _04649_ _04665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07207__I _01082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06845_ _02260_ _02283_ _02343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09564_ _04597_ _04569_ _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08515_ cpu.toggle_ctr\[5\] _03701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06776_ _02167_ _00987_ _02273_ _02274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05372__A2 _00882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05727_ _01232_ _01233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09495_ _04364_ _04523_ _04531_ _04446_ _04532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_78_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06321__A1 _01802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08446_ cpu.orig_PC\[11\] _03642_ _03645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05658_ _01148_ _01153_ _01163_ _01164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XPHY_EDGE_ROW_83_Left_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08377_ _00673_ _03594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05589_ _01090_ _01094_ _01095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_46_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07328_ _02774_ _00072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09297__C _04340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07259_ _01997_ _02721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05278__I3 cpu.regs\[11\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10270_ _00209_ clknet_leaf_63_wb_clk_i cpu.spi.data_out_buff\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09574__A1 _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_92_Left_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09326__A1 _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07117__I _02601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09332__I _04252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06312__A1 cpu.uart.divisor\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_12_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10606_ _00544_ clknet_leaf_61_wb_clk_i cpu.PORTA_DDR\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xclkbuf_leaf_88_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_88_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_37_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_17_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_17_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10537_ _00475_ clknet_4_8_0_wb_clk_i cpu.PC\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10468_ _00407_ clknet_leaf_30_wb_clk_i cpu.spi.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09935__C _04904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10399_ _00338_ clknet_leaf_8_wb_clk_i cpu.toggle_ctr\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08411__I _03586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06630_ _02126_ _02127_ _02128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06561_ _02057_ _02058_ _02059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XTAP_TAPCELL_ROW_86_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08300_ _02860_ _03527_ _03533_ _03414_ _00285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_87_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05512_ _01019_ net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09280_ _04042_ _04324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06492_ _01848_ _01920_ _01991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08231_ cpu.uart.data_buff\[7\] _03458_ _03483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05443_ _00935_ _00937_ _00942_ _00940_ _00953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_117_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08162_ _03426_ _03427_ _03428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05374_ _00885_ _00886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08093_ _03365_ _03371_ _03372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07113_ _02052_ _02483_ _02475_ _02598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__07803__A1 cpu.timer_div\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07044_ _02533_ _00029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08995_ cpu.IO_addr_buff\[6\] _04066_ _04077_ _04069_ _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07946_ _00975_ _03242_ _03252_ _03253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input27_I sram_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07877_ cpu.spi.div_counter\[1\] cpu.spi.divisor\[1\] _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09616_ cpu.last_addr\[3\] cpu.last_addr\[2\] _04647_ _04648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06828_ _02186_ _02263_ _02326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_66_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09547_ _04579_ _04580_ _04581_ _04582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06759_ _02255_ _02256_ _02257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08991__I _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09478_ _00802_ _04515_ _04516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07601__S _02968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_11_0_wb_clk_i clknet_0_wb_clk_i clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08429_ _03631_ _03632_ _03630_ _00315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_65_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output95_I net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10322_ _00261_ clknet_leaf_52_wb_clk_i cpu.uart.data_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10253_ _00192_ clknet_leaf_49_wb_clk_i cpu.spi.dout\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10184_ _00123_ clknet_leaf_4_wb_clk_i cpu.regs\[10\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_70_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05423__I3 cpu.regs\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08522__A2 cpu.toggle_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09665__C _04684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07261__A2 _02722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05090_ _00630_ _00631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_110_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07800_ _02520_ _03121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08780_ _03904_ _03899_ _03905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06772__A1 _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07731_ _00823_ _03052_ _03063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05992_ _01167_ _01495_ _01496_ _00014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07662_ _02980_ _03016_ _03018_ _00162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09401_ _04436_ _04439_ _04440_ _04441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06613_ _02105_ _02106_ _02111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07593_ cpu.regs\[8\]\[1\] _02971_ _02973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06544_ _00664_ _02042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_87_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09332_ _04252_ _04375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06475_ cpu.spi.divisor\[7\] _01628_ _01611_ _01974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09263_ _04302_ _04305_ _04306_ _04307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08029__A1 _02853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08029__B2 cpu.uart.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08214_ _00922_ _03455_ _03469_ _03470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09194_ _03613_ _00770_ _04240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_7_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05426_ _00905_ _00936_ _00907_ _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_08145_ _03310_ _03410_ _03412_ _03414_ _00249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_71_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05357_ _00006_ _00869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_101_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08076_ _03221_ cpu.spi.counter\[1\] _03099_ _03357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_05288_ cpu.regs\[1\]\[1\] _00820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07027_ _02519_ _02520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08978_ _04047_ _04062_ _04063_ _04064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07929_ _03230_ _03239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_59_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06515__A1 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_3_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09068__I0 cpu.regs\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07491__A2 _02903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_20_Left_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10305_ _00244_ clknet_leaf_40_wb_clk_i cpu.uart.div_counter\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_72_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10236_ _00175_ clknet_leaf_113_wb_clk_i cpu.regs\[4\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10167_ _00106_ clknet_leaf_4_wb_clk_i cpu.regs\[12\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10098_ _00041_ clknet_leaf_104_wb_clk_i cpu.br_rel_dest\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06506__A1 _01992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07305__I _02661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_32_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_32_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_72_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06809__A2 _00894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06260_ _00597_ _01760_ _01761_ _01762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_115_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05211_ _00731_ _00744_ _00747_ _00010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07040__I _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06191_ _01484_ _01693_ _01694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05142_ cpu.IO_addr_buff\[2\] _00680_ _00681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08431__A1 _02588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09950_ _04644_ _04915_ _04917_ _04918_ _04919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_05073_ _00614_ _00615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_94_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_49_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08901_ _02536_ _03998_ _03999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09881_ _04815_ _04866_ _04867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08832_ _03948_ _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06745__A1 _02108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08763_ _03885_ _03886_ _03148_ _03891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05975_ _01479_ _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_56_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07714_ _03048_ _00184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08694_ _03831_ _03179_ _03832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_0_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07170__A1 _02644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07645_ _02992_ _03001_ _03006_ _00157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07576_ _01145_ _01163_ _02964_ _02915_ _02965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_36_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09315_ _04274_ _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06527_ _01552_ _02006_ _02021_ _02025_ _02026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__10057__A1 _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09246_ _02797_ _04177_ _04290_ _04089_ _04291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06458_ _01956_ _01957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_105_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08670__A1 _01111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05409_ _00920_ _00921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06389_ _01881_ _01201_ _01887_ _01888_ _01502_ _01889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA_clkbuf_leaf_88_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09177_ _01271_ _01280_ _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08128_ _00792_ _03400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08422__A1 _02563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08059_ _02735_ _03344_ _03345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput57 net57 io_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput46 net46 io_oeb[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput35 net35 io_oeb[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput68 net68 io_out[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput79 net79 io_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10021_ _04980_ _04983_ _00760_ _04984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_8_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09922__A1 _00975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08489__A1 cpu.toggle_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07161__A1 _02636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08665__B _03811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_94_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09913__A1 cpu.PORTA_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07744__B _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10219_ _00158_ clknet_leaf_116_wb_clk_i cpu.regs\[6\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05760_ _00706_ _01038_ _01265_ _01266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_27_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05950__A2 _00929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05691_ _01196_ _01070_ _01176_ _01197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_43_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07430_ _02857_ _02862_ cpu.uart.receive_div_counter\[3\] _01612_ _02863_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_76_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_122_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07361_ _02800_ _02792_ _02789_ _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06312_ cpu.uart.divisor\[13\] _01502_ _01813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09100_ cpu.last_addr\[5\] _04157_ _04158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_61_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_33_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09031_ _04105_ _00444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07292_ _02670_ _02739_ _02745_ _02744_ _00065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05466__A1 _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06243_ _01744_ _01745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06174_ _01670_ _01676_ _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05125_ cpu.startup_cycle\[3\] cpu.startup_cycle\[2\] _00664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_clkbuf_leaf_5_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05769__A2 _01030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09933_ _04905_ _00546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05056_ _00598_ net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_09864_ _04840_ _04854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06718__A1 _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08815_ _03170_ _03928_ _03929_ _03934_ _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09795_ cpu.pwm_top\[5\] cpu.pwm_counter\[5\] _04799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08746_ _02720_ _03837_ _03832_ _03876_ _03845_ _03877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_05958_ _01438_ _01463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05889_ net7 _01206_ _01391_ _01393_ _01394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_67_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08677_ _02732_ _03817_ _03821_ _03820_ _00374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08891__A1 cpu.timer_div\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07628_ _02995_ _00151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07559_ cpu.regs\[10\]\[2\] _02951_ _02954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10570_ _00508_ clknet_leaf_75_wb_clk_i cpu.ROM_spi_dat_out\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_101_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09229_ _04236_ _04274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08504__I cpu.toggle_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10004_ _02464_ _04967_ _04968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_73_Right_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_103_Left_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07134__A1 _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08882__A1 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_82_Right_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09938__C _04904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_30_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07739__B _02072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_112_Left_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_91_Right_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05620__A1 _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06930_ _02403_ _02426_ _00022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_38_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I io_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08600_ cpu.pwm_counter\[3\] _03765_ _03767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06861_ _02355_ _02358_ _02359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09580_ _04513_ _04614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_38_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06792_ _00917_ _02289_ _02287_ _02290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05812_ _01317_ _00818_ _01318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05743_ cpu.timer_top\[0\] _01248_ _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08531_ cpu.toggle_ctr\[10\] _03717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07125__A1 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05674_ _01115_ _01082_ _01180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08462_ _02636_ _03655_ _03656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07413_ cpu.uart.receive_div_counter\[14\] _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08873__A1 cpu.timer_div\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07676__A2 _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08393_ _03604_ _03589_ _03605_ _03591_ _00306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_57_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08625__A1 _02754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07344_ _02783_ _02547_ _02567_ _02784_ _02785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_73_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07275_ cpu.timer_top\[2\] _02730_ _02734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08324__I _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06226_ _01708_ _01248_ _01726_ _01727_ _01640_ _01728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_60_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09014_ _04092_ _00440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07368__C _02567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06157_ _01658_ _01659_ _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05108_ cpu.IO_addr_buff\[1\] _00647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06088_ _01332_ _01591_ _01592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09916_ _03236_ _04893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05039_ _00577_ _00578_ _00581_ _00582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09847_ _04840_ _04841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09778_ _04784_ _04785_ _04786_ _00510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08729_ cpu.timer\[4\] _03811_ _03834_ _03862_ _03856_ _03863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_68_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05470__S0 _00871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08864__A1 _02670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09758__C _04765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10622_ _00560_ clknet_leaf_3_wb_clk_i cpu.regs\[15\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10553_ _00491_ clknet_leaf_72_wb_clk_i cpu.mem_cycle\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_64_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10484_ _00422_ clknet_leaf_40_wb_clk_i cpu.uart.divisor\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09592__A2 _00772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07107__A1 _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07313__I _01005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05390_ _00901_ _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_82_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07060_ _02548_ _02385_ _02549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06011_ _01514_ _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_70_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09583__A2 _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09701_ _04710_ _04708_ _04723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07962_ _03265_ _00215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07893_ _03206_ _03209_ _03210_ _00201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06913_ _02367_ _02369_ _02372_ _02410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09632_ cpu.last_addr\[7\] cpu.ROM_addr_buff\[7\] _04650_ _04664_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_65_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06844_ _02322_ _02340_ _02341_ _02302_ _02342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__08747__C _03795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09563_ cpu.PC\[12\] _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08514_ _03699_ cpu.toggle_top\[6\] _03700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06775_ _02265_ _02262_ _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_81_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05726_ _01045_ _01081_ _01186_ _01232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09494_ _03637_ _04028_ _04531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08445_ _03090_ _03633_ _03644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05657_ _01155_ _01158_ _01162_ _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_37_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08376_ cpu.IO_addr_buff\[5\] _03592_ _03593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05588_ _00721_ _01092_ _01093_ _01094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_45_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07327_ cpu.toggle_top\[14\] _02761_ _02770_ _02773_ _02774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_34_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07258_ cpu.timer\[7\] _02720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06209_ cpu.PORTA_DDR\[4\] _01613_ _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07189_ _02660_ _02661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07585__A1 _01910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output40_I net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09769__B _00790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10605_ _00543_ clknet_leaf_61_wb_clk_i cpu.PORTA_DDR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_64_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10536_ _00474_ clknet_4_8_0_wb_clk_i cpu.PC\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_108_Right_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10467_ _00406_ clknet_leaf_30_wb_clk_i cpu.spi.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05823__A1 _01311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_57_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_57_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10398_ _00337_ clknet_leaf_7_wb_clk_i cpu.toggle_ctr\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07308__I _02647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05256__C _00791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08525__B1 cpu.toggle_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06000__A1 cpu.uart.divisor\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06560_ cpu.mem_cycle\[2\] _02058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_87_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08828__A1 _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05511_ _00773_ _01007_ _01018_ _01019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_59_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06491_ _00646_ _01990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08230_ _03482_ _00266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05442_ _00951_ _00952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08161_ _03422_ _03427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05373_ _00869_ _00885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08092_ _03323_ _03338_ _03344_ _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_07112_ _02048_ _02466_ _02597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_43_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09005__A1 _02517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07043_ _02530_ _02514_ _02532_ _02522_ _02533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08602__I _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08994_ _04047_ _04075_ _04076_ _04077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07945_ cpu.spi.data_out_buff\[2\] _03243_ _03252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07319__A1 _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09615_ cpu.last_addr\[1\] cpu.last_addr\[0\] _04647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07876_ cpu.spi.div_counter\[6\] _03196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__05961__I _01465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05425__S0 _00872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06827_ _02316_ _02324_ _02325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09546_ cpu.PC\[10\] _01323_ _04581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06758_ _02253_ _02254_ _02256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05709_ _01107_ _01177_ _01215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_65_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09477_ _04513_ _04515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08428_ cpu.orig_PC\[6\] _03628_ _03632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06689_ cpu.regs\[1\]\[7\] _01994_ _02186_ _02187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_80_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08047__A2 _01962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08359_ _03578_ _03581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10321_ _00260_ clknet_leaf_50_wb_clk_i cpu.uart.counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10252_ _00191_ clknet_leaf_50_wb_clk_i cpu.spi.dout\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10183_ _00122_ clknet_leaf_126_wb_clk_i cpu.regs\[10\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06230__A1 cpu.toggle_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_104_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_104_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_57_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_53_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10519_ _00457_ clknet_leaf_77_wb_clk_i cpu.last_addr\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_39_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07549__A1 cpu.regs\[11\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07730_ _03053_ _03060_ _03061_ _03062_ _00186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_34_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05991_ cpu.regs\[9\]\[1\] _01375_ _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_88_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07661_ cpu.regs\[5\]\[0\] _03017_ _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09400_ _04274_ _04440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06612_ _02109_ _01294_ _02110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07592_ _02914_ _02970_ _02972_ _00138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06543_ _02038_ _02040_ _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09331_ _04347_ _04352_ _04372_ _04373_ _04374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_48_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06474_ cpu.uart.dout\[7\] _01195_ _01970_ _01972_ _01102_ _01973_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_09262_ _04274_ _04306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07501__I _01373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_78_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08213_ cpu.uart.data_buff\[3\] _03464_ _03469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09193_ _00738_ _00780_ _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_05425_ cpu.regs\[4\]\[2\] cpu.regs\[5\]\[2\] cpu.regs\[6\]\[2\] cpu.regs\[7\]\[2\]
+ _00872_ _00874_ _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XTAP_TAPCELL_ROW_99_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08144_ _03413_ _03414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_43_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05356_ _00867_ _00868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_43_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08075_ _03354_ _03356_ _00236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05287_ cpu.regs\[4\]\[1\] cpu.regs\[5\]\[1\] cpu.regs\[6\]\[1\] cpu.regs\[7\]\[1\]
+ _00803_ _00573_ _00819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07026_ _00685_ _02519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06212__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07960__A1 _02664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08977_ _02615_ _04030_ _04063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_2_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_2_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07928_ _03229_ _03238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07859_ _03137_ _03179_ _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_3_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08000__C _02628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09529_ _04455_ _04547_ _04564_ _04541_ _04565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08507__I cpu.toggle_top\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09217__A1 _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09766__C _04765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09338__I _00689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10304_ _00243_ clknet_leaf_39_wb_clk_i cpu.uart.div_counter\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09782__B _00790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10235_ _00174_ clknet_leaf_112_wb_clk_i cpu.regs\[4\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07951__A1 _02652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10166_ _00105_ clknet_leaf_124_wb_clk_i cpu.regs\[13\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10097_ _00040_ clknet_leaf_104_wb_clk_i cpu.br_rel_dest\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09006__C _04020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07703__A1 cpu.regs\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07522__S _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_112_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09208__A1 _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05210_ _00746_ _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06190_ _01680_ _01691_ _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_4_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_72_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_72_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09676__C _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05141_ _00676_ _00679_ _00680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05245__A2 _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05072_ _00599_ _00608_ _00613_ _00614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__06442__A1 _01471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09880_ _04864_ _04866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_94_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08900_ _03997_ _03998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08195__A1 _03439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08831_ cpu.timer_capture\[13\] _03941_ _03947_ _03939_ _03948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_0_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07942__A1 _00947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08762_ _03148_ _03885_ _03886_ _03890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_05974_ _00991_ _01323_ _00657_ _01479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_79_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08693_ _03136_ _03831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07713_ _03011_ cpu.regs\[3\]\[6\] _03038_ _03048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07644_ cpu.regs\[6\]\[3\] _03000_ _03006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07575_ _02961_ _02963_ _01153_ _02964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_TAPCELL_ROW_36_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09314_ _04353_ _04352_ _04355_ _04356_ _04357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06526_ _01449_ _02001_ _02022_ _02024_ _02025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_09245_ _00729_ _00784_ _03594_ _04289_ _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_8_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06457_ _01955_ _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08771__B _03897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05408_ _00919_ _00920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06388_ net13 _01517_ _01207_ _01888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_90_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09176_ _00708_ _01265_ _04223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08127_ _03398_ _03399_ _00246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05339_ cpu.PORTA_DDR\[6\] net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_102_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08058_ _03342_ _03343_ _03344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08062__I _02735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06433__B2 _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput58 net58 io_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_07009_ cpu.ROM_addr_buff\[3\] _02501_ _02502_ cpu.ROM_addr_buff\[7\] _02477_ _02503_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
Xoutput47 net47 io_oeb[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput36 net36 io_oeb[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput69 net69 io_out[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10020_ _01021_ _04180_ _04982_ _04983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_8_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06292__S0 _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05635__B _00992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08665__C _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06672__B2 _00801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10218_ _00157_ clknet_leaf_109_wb_clk_i cpu.regs\[6\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10149_ _00088_ clknet_leaf_43_wb_clk_i cpu.uart.receive_counter\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05690_ _01044_ _01196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_85_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10039__A2 _02722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07360_ _01493_ _02780_ _02799_ _02800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06311_ _01804_ _01207_ _01810_ _01811_ _01502_ _01812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_61_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_33_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09030_ _04103_ cpu.ROM_addr_buff\[2\] _04104_ _04105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07291_ cpu.timer_top\[7\] _02740_ _02745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05466__A2 _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06242_ _01743_ _01742_ _01744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09601__A1 _00751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06173_ _01551_ _00956_ _01584_ _01676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05124_ cpu.startup_cycle\[6\] cpu.startup_cycle\[5\] cpu.startup_cycle\[4\] _00663_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_41_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09932_ cpu.PORTA_DDR\[5\] _04899_ _04903_ _04904_ _04905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_40_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05055_ _00597_ _00598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_1_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09863_ _04840_ _04853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_5_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08814_ _02692_ _03930_ _03934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09794_ _04796_ _03758_ _04797_ cpu.pwm_top\[1\] _04798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_08745_ cpu.timer\[7\] _03871_ _03876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_108_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05957_ _01461_ _01462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05888_ _01392_ _01393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08676_ cpu.timer_top\[9\] _03818_ _03821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07627_ _02943_ cpu.regs\[7\]\[5\] _02983_ _02995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07558_ _02921_ _02950_ _02953_ _00123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06509_ net96 _01800_ _02008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09840__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07489_ cpu.regs\[13\]\[2\] _02905_ _02908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09228_ _04269_ _04271_ _04272_ _04273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09159_ _00997_ _00988_ _01018_ _04206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_44_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output70_I net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10003_ _02042_ _04706_ _04966_ _02453_ _04967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07136__I _02617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07134__A2 _02601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05448__A2 _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09300__B _03853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07070__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08430__I _03586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05620__A2 _01106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06860_ _02356_ _02357_ _02358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07046__I _00787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05811_ cpu.br_rel_dest\[0\] _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__05384__A1 _00868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06791_ _00849_ _00926_ _02289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05742_ _01247_ _01248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08530_ _03715_ _01261_ _03694_ _03696_ _03716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05673_ _01178_ _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08461_ _03653_ _03655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07412_ _02828_ _02831_ _02837_ _02844_ _02845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_18_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08392_ cpu.orig_flags\[1\] _03587_ _03605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07343_ _02406_ _02168_ _02552_ _02784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07274_ _02732_ _02729_ _02733_ _00791_ _00059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_72_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06225_ cpu.timer_capture\[12\] _01233_ _01639_ _01727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09013_ _00952_ _04084_ _04091_ _04089_ _04092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_14_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08389__A1 cpu.orig_flags\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06156_ _01556_ _01561_ _01555_ _01659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_111_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06087_ _01574_ _01589_ _01591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05107_ _00646_ net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_0_111_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09915_ _04819_ _04889_ _04892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05038_ _00580_ _00581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09846_ _01063_ _04812_ _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09777_ cpu.ROM_spi_cycle\[1\] _04781_ _04786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06989_ _02467_ _02483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08728_ _03860_ _03861_ _03862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05470__S1 _00977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08659_ _03801_ _03807_ _03808_ _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_95_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10621_ _00559_ clknet_leaf_2_wb_clk_i cpu.regs\[15\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10552_ _00490_ clknet_leaf_62_wb_clk_i cpu.mem_cycle\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10483_ _00012_ clknet_leaf_44_wb_clk_i cpu.uart.clr_hb vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_114_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07052__A1 _01137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05874__I _01158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06866__A1 _02090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05133__A4 _00671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06618__A1 cpu.regs\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06010_ _01088_ _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_70_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09032__A2 _00851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07961_ cpu.spi.data_out_buff\[6\] _03255_ _03264_ _03258_ _03265_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09700_ _02459_ _04716_ _04722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06912_ _02063_ _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07892_ cpu.spi.div_counter\[2\] _03208_ _03210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09631_ cpu.last_addr\[8\] cpu.ROM_addr_buff\[8\] _04651_ _04663_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_06843_ _02286_ _02301_ _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09562_ _02393_ _04520_ _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06774_ _02266_ _02271_ _02272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05725_ _01185_ _01229_ _01230_ _01231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08513_ _03698_ _03699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07504__I _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09493_ _04299_ _04523_ _04529_ _04310_ _04530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_08444_ _03640_ _03596_ _03643_ _00319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06857__A1 _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05024__I _00566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05656_ _01161_ _01147_ _01158_ _00924_ _01162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_105_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08375_ _03579_ _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05587_ _00659_ _01037_ _00652_ _01093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_116_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07326_ _02772_ _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07257_ _02719_ _00056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06208_ cpu.uart.divisor\[4\] _01710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_103_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07188_ _02519_ _02660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_60_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06139_ _01609_ _01414_ _01638_ _01641_ _01252_ _01642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__08782__A1 cpu.timer_capture\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07585__A2 _01948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09829_ _04827_ _00520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05348__A1 net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07414__I cpu.uart.divisor\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10604_ _00542_ clknet_leaf_61_wb_clk_i cpu.PORTA_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_40_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07273__A1 cpu.timer_top\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10535_ _00473_ clknet_leaf_89_wb_clk_i cpu.PC\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10466_ _00405_ clknet_leaf_30_wb_clk_i cpu.spi.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_29_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10397_ _00336_ clknet_leaf_6_wb_clk_i cpu.toggle_ctr\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07576__A2 _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_97_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_97_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_19_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_26_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_26_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_48_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06490_ _01953_ _01305_ _01987_ _01988_ _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_19_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05510_ _01017_ _01018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_118_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07500__A2 _02905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05441_ _00950_ _00951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_68_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08160_ cpu.uart.div_counter\[13\] _03426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07111_ cpu.rom_data_dist _02596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_7_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05372_ _00006_ _00882_ _00883_ _00884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_27_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08091_ _03369_ _03370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_70_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07042_ _02515_ _02531_ _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05814__A2 _00894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07016__A1 _00793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05370__S0 _00878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08104__B _03381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05578__A1 _01054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08993_ _01877_ _04030_ _04076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07944_ _03251_ _00211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07875_ cpu.spi.div_counter\[3\] _03195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09614_ _02051_ _04645_ _04646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06826_ _02312_ _02313_ _02308_ _02324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05425__S1 _00874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09545_ _04550_ _04580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06757_ _02253_ _02254_ _02255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05708_ _01113_ _01212_ _01213_ _01090_ _01214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_93_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09476_ _04513_ _04514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_38_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06688_ _00876_ _00881_ _00884_ _00891_ _02185_ _02186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_93_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08427_ _02586_ _03619_ _03631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05639_ _01144_ _01145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_08358_ _03579_ _03580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08289_ _03522_ _03524_ _00283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_61_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07309_ _02758_ _02750_ _02759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10320_ _00259_ clknet_leaf_51_wb_clk_i cpu.uart.counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10251_ _00190_ clknet_leaf_65_wb_clk_i cpu.spi.dout\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10182_ _00121_ clknet_leaf_125_wb_clk_i cpu.regs\[11\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_70_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_102_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07080__S _02567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10518_ _00456_ clknet_leaf_78_wb_clk_i cpu.last_addr\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08703__I _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10449_ _00388_ clknet_leaf_25_wb_clk_i cpu.timer\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07763__B _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05990_ _01494_ _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_88_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07660_ _03014_ _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_27_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06611_ _02108_ _02109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_07591_ cpu.regs\[8\]\[0\] _02971_ _02972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06542_ _02039_ _02040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09330_ _04330_ _04373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09261_ _04303_ _04304_ _04305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06473_ _01522_ _01971_ _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08212_ _03468_ _00262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09226__A2 _00771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09192_ _02781_ _04237_ _04238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_16_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05424_ _00870_ _00934_ _00935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_28_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08143_ _00779_ _03413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05355_ _00866_ _00867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08074_ _03099_ _03349_ _03355_ _03348_ _03356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_102_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07025_ _02515_ _02517_ _02518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05286_ _00818_ net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_30_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08737__A1 cpu.timer_capture\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input32_I sram_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08976_ cpu.orig_IO_addr_buff\[3\] _04044_ _04045_ _00998_ _04062_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07927_ _03236_ _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07858_ _03178_ _03179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_07789_ _03112_ _03114_ _00747_ _00193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05723__A1 cpu.spi.dout\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06809_ _00850_ _00894_ _02307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09528_ _00837_ _04515_ _04564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_104_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09459_ _04465_ _04495_ _04496_ _04497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_81_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07228__A1 cpu.timer_capture\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08976__B2 _00998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10303_ _00242_ clknet_leaf_42_wb_clk_i cpu.uart.div_counter\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10234_ _00173_ clknet_leaf_109_wb_clk_i cpu.regs\[4\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10165_ _00104_ clknet_leaf_121_wb_clk_i cpu.regs\[13\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06203__A2 _01010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10096_ _00039_ clknet_leaf_104_wb_clk_i cpu.br_rel_dest\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05962__A1 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05714__A1 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07703__A2 _03041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05323__S _00581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05140_ _00677_ _00678_ _00679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_53_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05071_ _00567_ _00610_ _00612_ _00613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
Xclkbuf_leaf_41_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_41_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_94_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08195__A2 _03450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08830_ _03920_ _03946_ _03947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08761_ _03888_ _03889_ _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05953__A1 _01454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05973_ _01442_ _01477_ _01478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08692_ _02670_ _03824_ _03830_ _03827_ _00380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07712_ _03047_ _00183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07713__S _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07643_ _02990_ _03001_ _03005_ _00156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09313_ _04326_ _04356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07574_ _01175_ _01215_ _01263_ _02962_ _02963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_48_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07512__I _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06525_ _02007_ _02023_ _01480_ _02024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_36_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09244_ _00729_ _04288_ _04289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06456_ _01954_ _01955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_90_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09175_ _01093_ _04221_ _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05407_ _00918_ _00919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05032__I _00574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06387_ net4 _01389_ _01884_ _01886_ _01109_ _01887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_08126_ _03331_ _03394_ _03237_ _03399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05338_ cpu.PORTB_DDR\[6\] net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_0_113_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08057_ cpu.uart.counter\[3\] cpu.uart.counter\[2\] _03343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05269_ cpu.regs\[2\]\[0\] _00802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07008_ _02479_ _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xoutput48 net48 io_oeb[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_12_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput37 net37 io_oeb[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput59 net59 io_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08959_ _01317_ _04039_ _04041_ _04046_ _04047_ _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__06292__S1 _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06466__C _01215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06121__A1 _01612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05307__S0 _00570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06424__A2 _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10217_ _00156_ clknet_leaf_108_wb_clk_i cpu.regs\[6\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10148_ _00087_ clknet_leaf_39_wb_clk_i cpu.uart.receive_counter\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10079_ _00022_ clknet_leaf_111_wb_clk_i cpu.regs\[2\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09812__I _04813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06310_ net11 _01205_ _01200_ _01811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07290_ _02665_ _02739_ _02743_ _02744_ _00064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_33_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06241_ _01740_ _01743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_96_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07860__A1 _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05466__A3 _00975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06172_ _01471_ _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05123_ cpu.startup_cycle\[1\] cpu.startup_cycle\[0\] _00662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_111_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09931_ _03236_ _04904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05054_ _00596_ _00597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09365__A1 _02563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09862_ _04852_ _00528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_110_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06179__A1 _01161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08813_ _03933_ _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09793_ cpu.pwm_counter\[1\] _04797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05926__A1 _00721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08744_ _03874_ _03875_ _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05956_ _01460_ _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_84_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08766__C _03616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05887_ net22 _01218_ _01109_ _01392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08675_ _02726_ _03817_ _03819_ _03820_ _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_95_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07626_ _02994_ _00150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07557_ cpu.regs\[10\]\[1\] _02951_ _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08782__B _03761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06508_ _01993_ _01998_ _02007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07488_ _01495_ _02904_ _02907_ _00099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07851__A1 cpu.timer_top\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07851__B2 cpu.timer_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09227_ _02608_ _04269_ _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06439_ _01360_ _01918_ _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_91_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09158_ _01468_ _04198_ _04201_ _04204_ _02027_ _04205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_0_32_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08109_ _03311_ _03382_ _03385_ _03306_ _00242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09089_ _03360_ _04148_ _04149_ _00458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_31_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08801__I _03921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output63_I net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10002_ _04718_ _02040_ _04966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05917__A1 _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_80_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08095__A1 _00793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_17_Left_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07842__B2 cpu.timer_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_26_Left_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05810_ _01131_ _00816_ _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_89_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06581__A1 _02078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06790_ _00822_ _02288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05384__A2 _00895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05741_ _01246_ _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05672_ _01104_ _01177_ _01178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08460_ _03653_ _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07411_ _02838_ _02839_ _02843_ _02844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_77_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08391_ cpu.Z _03604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_18_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07062__I _02063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_35_Left_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_70_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07342_ _02782_ _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07273_ cpu.timer_top\[1\] _02730_ _02733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06097__B1 _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06224_ cpu.timer_capture\[4\] _01633_ _01723_ _01725_ _01241_ _01726_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_61_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09012_ _02527_ _04085_ _04091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06155_ _01656_ _01657_ _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_1_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_44_Left_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05106_ _00599_ _00640_ _00645_ _00646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_06086_ _01574_ _01589_ _01590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09914_ _04891_ _00541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05037_ _00579_ _00580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09845_ _04839_ _00524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_95_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08777__B _03897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09776_ cpu.ROM_spi_cycle\[1\] _04781_ _04785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06988_ _02044_ _02481_ _02482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08727_ cpu.timer\[3\] _03849_ cpu.timer\[4\] _03861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05939_ _01315_ _01443_ _01444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08658_ cpu.timer_div_counter\[3\] _03804_ cpu.timer_div_counter\[4\] _03808_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_53_Left_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_4_8_0_wb_clk_i clknet_0_wb_clk_i clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07609_ _02981_ _02982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_08589_ _03758_ _03759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09401__B _04440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07700__I _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10620_ _00558_ clknet_leaf_2_wb_clk_i cpu.regs\[15\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10551_ _00489_ clknet_leaf_61_wb_clk_i cpu.mem_cycle\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10482_ _00421_ clknet_leaf_87_wb_clk_i cpu.rom_data_dist vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_19_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_62_Left_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_71_Left_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06315__A1 cpu.spi.divisor\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_58_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08706__I _03835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09568__A1 _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07960_ _02664_ _03241_ _03263_ _03264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07057__I _02541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06911_ cpu.PC\[13\] _02394_ _02408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07891_ cpu.spi.div_counter\[2\] _03208_ _03209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09630_ cpu.last_addr\[9\] cpu.ROM_addr_buff\[9\] _04661_ _04662_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_4_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06842_ _02339_ _02338_ _02340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_09561_ _04567_ _04595_ _00690_ _00484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_97_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05506__S _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06773_ _02269_ _02270_ _02271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05724_ cpu.timer_div\[0\] _01185_ _01230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08512_ cpu.toggle_ctr\[6\] _03698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06306__A1 net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09492_ _04526_ _04527_ _04528_ _04529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_93_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08443_ _03641_ _03642_ _03116_ _03643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_65_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06857__A2 _02092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05655_ _01160_ _01161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_86_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08059__A1 _02735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08374_ _00677_ _03589_ _03590_ _03591_ _00301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05586_ _00651_ _00655_ _01091_ _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_46_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07325_ _02771_ _02772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_90_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07256_ cpu.timer_capture\[6\] _02701_ _02718_ _02712_ _02719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_46_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06207_ cpu.spi.dout\[4\] _01709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__09559__A1 _04256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05040__I _00581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07187_ _02658_ _02654_ _02659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05975__I _01479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06138_ cpu.timer_top\[3\] _01639_ _01640_ _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06069_ _01350_ _01556_ _01559_ _01452_ _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09828_ net62 _04814_ _04826_ _04821_ _04827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05348__A2 cpu.ROM_spi_mode vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09759_ _04772_ _00505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08298__A1 _03495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06474__C _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10603_ _00541_ clknet_leaf_62_wb_clk_i cpu.PORTA_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_64_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10534_ _00472_ clknet_leaf_91_wb_clk_i cpu.Z vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08470__A1 _02754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06046__I _00845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10465_ _00404_ clknet_leaf_23_wb_clk_i cpu.timer_capture\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07025__A2 _02517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10396_ _00335_ clknet_leaf_7_wb_clk_i cpu.toggle_ctr\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07576__A3 _02964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08525__A2 cpu.toggle_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09820__I _04683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_66_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_66_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_35_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05440_ cpu.base_address\[2\] _00950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07340__I cpu.PC\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05371_ _00007_ _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_83_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07110_ _02517_ _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08090_ _03344_ _03368_ _03369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_43_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07041_ net20 _02516_ _02531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_2_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05370__S1 _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10020__A1 _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08992_ cpu.orig_IO_addr_buff\[6\] _04044_ _04045_ _01957_ _04075_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07943_ cpu.spi.data_out_buff\[2\] _03234_ _03250_ _03247_ _03251_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07874_ _03188_ cpu.spi.divisor\[4\] cpu.spi.div_counter\[6\] _03192_ _03193_ _03194_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__08516__A2 _01419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09613_ _04644_ _02598_ _04645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06825_ _02317_ _02319_ _02323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07515__I _01700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09544_ cpu.PC\[10\] _01323_ _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06756_ _02222_ _02223_ _02226_ _02254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_05707_ net39 _01113_ _01213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06687_ _00800_ _02185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_09475_ _01366_ _01324_ _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_93_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08426_ _03627_ _03629_ _03630_ _00314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_65_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05638_ _01033_ _01141_ _01143_ _01144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_05569_ _01073_ _01074_ _01075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08357_ _03578_ _03579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08288_ cpu.uart.receive_div_counter\[3\] _03511_ _03523_ _02869_ _03524_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_104_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07308_ _02647_ _02758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07239_ _00989_ _02697_ _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10250_ _00189_ clknet_leaf_101_wb_clk_i cpu.regs\[2\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09952__A1 _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05569__A2 _01074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10181_ _00120_ clknet_leaf_119_wb_clk_i cpu.regs\[11\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06518__A1 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07160__I _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08443__A1 _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10517_ _00455_ clknet_leaf_79_wb_clk_i cpu.ROM_addr_buff\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_113_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_113_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_110_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10448_ _00387_ clknet_leaf_25_wb_clk_i cpu.timer\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09943__A1 cpu.ROM_spi_mode vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10379_ _00318_ clknet_leaf_85_wb_clk_i cpu.orig_PC\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06509__A1 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07182__A1 _02653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_9_Left_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06610_ _00850_ _02108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07590_ _02968_ _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06541_ cpu.startup_cycle\[0\] _02039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_87_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10069__A1 _02032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06472_ cpu.uart.divisor\[15\] _01503_ _01971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09260_ _02383_ _01159_ _04304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08211_ cpu.uart.data_buff\[1\] _03460_ _03466_ _03467_ _03468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05423_ cpu.regs\[0\]\[2\] cpu.regs\[1\]\[2\] cpu.regs\[2\]\[2\] cpu.regs\[3\]\[2\]
+ _00872_ _00874_ _00934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__07485__A2 _02905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09191_ _01317_ _04236_ _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08142_ cpu.uart.div_counter\[9\] _03383_ _03411_ _03378_ _03412_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_99_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05354_ _00716_ _00866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08073_ _03099_ _03352_ _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_102_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05099__I1 _00638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05285_ _00817_ _00818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06996__A1 _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07024_ net1 _02516_ _02517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_11_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09934__A1 _02664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08975_ _04055_ _04061_ _00432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07926_ _02520_ _03236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input25_I rst_n vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05971__A2 _01345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07857_ _01607_ _03177_ _03178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07788_ cpu.spi.dout\[3\] _03113_ _03114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06920__A1 _02416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06808_ _00822_ _00955_ _02306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09527_ _04514_ _04547_ _04563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06739_ _00849_ _00953_ _02237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09458_ _02379_ _01036_ _04496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08409_ cpu.orig_PC\[1\] _03607_ _03618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09389_ _04333_ _04412_ _04429_ _04378_ _04403_ _04430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_50_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10302_ _00241_ clknet_leaf_42_wb_clk_i cpu.uart.div_counter\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output93_I net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10233_ _00172_ clknet_leaf_107_wb_clk_i cpu.regs\[4\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10164_ _00103_ clknet_leaf_122_wb_clk_i cpu.regs\[13\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05411__A1 _00865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10095_ _00038_ clknet_leaf_104_wb_clk_i cpu.br_rel_dest\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05962__A2 _01354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05714__A2 _01053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06911__A1 cpu.PC\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07104__B _02407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05070_ _00583_ _00611_ _00612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_6_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_10_0_wb_clk_i clknet_0_wb_clk_i clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_57_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_81_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_81_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08760_ cpu.timer_capture\[9\] _03883_ _03869_ _03889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05972_ _01310_ _01362_ _01476_ _01477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08691_ cpu.timer_top\[15\] _03825_ _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_10_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_10_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07711_ _03009_ cpu.regs\[3\]\[5\] _03038_ _03047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07642_ cpu.regs\[6\]\[2\] _03002_ _03005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06902__A1 _00591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09312_ cpu.orig_PC\[3\] _04354_ _04355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07573_ _01114_ _01173_ _01254_ _02962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_48_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06524_ _01926_ _02008_ _02023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_36_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09243_ _04265_ _04267_ _04287_ _04256_ _04288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06455_ _01797_ _01794_ _00913_ _01954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10078__D _00021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06386_ _01217_ _01885_ _01886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08407__A1 _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09174_ _01270_ _04210_ _04179_ _04221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05406_ _00917_ _00918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08125_ _03331_ _03374_ _03397_ _03390_ _03398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05337_ cpu.PORTA_DDR\[5\] net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_44_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08056_ cpu.uart.counter\[0\] cpu.uart.counter\[1\] _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_05268_ _00800_ _00801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09907__A1 cpu.PORTB_DDR\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07007_ _02474_ _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05199_ _00671_ _00734_ _00735_ _00692_ _00736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_3_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput49 net49 io_oeb[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_12_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput38 net38 io_oeb[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08958_ _04031_ _04047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07909_ cpu.spi.counter\[0\] _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08889_ _03989_ _00418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07146__A1 _01877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07697__A2 _02932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05307__S1 _00574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07621__A2 _02985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09374__A2 _00756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10216_ _00155_ clknet_leaf_12_wb_clk_i cpu.regs\[6\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10147_ _00086_ clknet_leaf_39_wb_clk_i cpu.uart.receive_counter\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06003__B cpu.PORTA_DDR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10078_ _00021_ clknet_leaf_111_wb_clk_i cpu.regs\[2\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05699__A1 _01196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08885__A1 _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07613__I _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_99_Left_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06240_ _00597_ _01004_ _01742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07860__A2 _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06171_ _01452_ _01671_ _01666_ _01466_ _01673_ _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_13_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05122_ _00652_ _00655_ _00658_ _00660_ _00661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_4_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09930_ _02657_ _04900_ _04903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05053_ _00567_ _00582_ _00595_ _00596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09861_ net82 _04841_ _04851_ _04847_ _04852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_111_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06179__A2 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08812_ cpu.timer_capture\[9\] _03919_ _03932_ _03916_ _03933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_09792_ cpu.pwm_top\[0\] _04796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05926__A2 _01156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08743_ cpu.timer_capture\[6\] _03858_ _03869_ _03875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05955_ _01347_ _00867_ _01330_ _01460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_108_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05886_ _01090_ _01387_ _01388_ _01390_ _01391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_08674_ _02736_ _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07625_ _02941_ cpu.regs\[7\]\[4\] _02984_ _02994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07556_ _02914_ _02950_ _02952_ _00122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05043__I _00002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06507_ _01991_ _02005_ _02006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_90_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07300__A1 _02732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09226_ _02796_ _00771_ _04270_ _04271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07487_ cpu.regs\[13\]\[1\] _02905_ _02907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06438_ _01484_ _01930_ _01932_ _01461_ _01937_ _01938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_90_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10536__D _00474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06369_ net95 _01365_ _01869_ _01870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09157_ _01870_ _01946_ _04203_ _04204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08108_ cpu.uart.div_counter\[2\] _03383_ _03384_ _03378_ _03385_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09088_ cpu.last_addr\[2\] _04143_ _04149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08039_ cpu.uart.div_counter\[14\] _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_31_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08303__B _03529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09118__C _03980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10001_ _02497_ _04964_ _04965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08022__C _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output56_I net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05473__S0 _00877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_48_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_80_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07358__A1 _02797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09823__I _00946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07544__S _02933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_87_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_38_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06581__A2 _01996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08858__A1 _02653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05740_ _01063_ _01116_ _01246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_54_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05671_ _00676_ _01077_ _01176_ _01177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_07410_ _02827_ cpu.uart.receive_div_counter\[8\] _02832_ cpu.uart.divisor\[7\] _02842_
+ _02843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_08390_ _01311_ _03589_ _03603_ _03591_ _00305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_58_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07341_ _02781_ _02782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05798__I _01131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07272_ _00922_ _02732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_45_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06223_ _01633_ _01724_ _01725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09011_ _04090_ _00439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09586__A2 _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06154_ net93 _00997_ _01657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_103_Right_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05105_ _00599_ _00642_ _00644_ _00645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06085_ _01575_ _01485_ _01589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09913_ cpu.PORTA_DDR\[0\] _04888_ _04890_ _04881_ _04891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05036_ _00002_ _00579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09844_ net67 _04828_ _04838_ _04833_ _04839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09733__I _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09775_ _03812_ _04783_ _04784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06987_ _02472_ _02051_ _00694_ _02481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__08849__A1 cpu.spi.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08726_ _02702_ _02696_ _03854_ _03860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_05938_ _01346_ _01442_ _01443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_96_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08657_ cpu.timer_div_counter\[3\] cpu.timer_div_counter\[4\] _03804_ _03807_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_05869_ _01166_ _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07608_ _01144_ _01163_ _02888_ _02981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_83_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08588_ cpu.pwm_counter\[0\] _03758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06088__A1 _01332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07539_ _02925_ _02935_ _02940_ _00117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_37_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10550_ _00488_ clknet_leaf_72_wb_clk_i cpu.mem_cycle\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10481_ _00420_ clknet_leaf_51_wb_clk_i cpu.timer_div\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09209_ _02327_ _04253_ _04254_ _04249_ _04255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__09577__A2 _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07629__S _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_121_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06012__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_4_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09818__I _00921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09568__A2 _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08240__A2 _03451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06910_ _02374_ _02407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07890_ _03206_ _03207_ _03208_ _00200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__06003__A1 _01196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09040__I1 cpu.ROM_addr_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06841_ _02304_ _02321_ _02339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07751__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09560_ _04487_ _04591_ _04592_ _04594_ _04049_ _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06772_ _00836_ _00994_ _02270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05723_ cpu.spi.dout\[0\] _01189_ _01192_ _01228_ _01229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10540__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08511_ cpu.toggle_ctr\[7\] _03697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09491_ _04526_ _04527_ _04440_ _04528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08442_ _03595_ _03642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07503__A1 _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07801__I _03121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05654_ _01159_ _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_105_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08373_ _03413_ _03591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05585_ _01027_ _01091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_116_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07324_ _02519_ _02771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_46_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07255_ _02678_ _02717_ _02718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09008__A1 _02524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05321__I cpu.regs\[2\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06206_ cpu.timer_top\[4\] _01708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_6_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06490__A1 _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07186_ _02657_ _02658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06137_ _01123_ _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07248__I _02661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06068_ _00945_ _01353_ _01555_ _01341_ _01356_ _01572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_111_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08788__B _03897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05428__S0 _00872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09827_ _04010_ _04816_ _04826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09758_ cpu.ROM_spi_dat_out\[4\] _04760_ _04771_ _04765_ _04772_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08300__C _03414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08709_ _03180_ _03844_ _03845_ _03846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09689_ _02038_ _04709_ _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_69_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08807__I _03921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10602_ _00540_ clknet_leaf_62_wb_clk_i cpu.PORTB_DDR\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_40_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10533_ _00471_ clknet_leaf_88_wb_clk_i cpu.IE vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06481__A1 _01960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10464_ _00403_ clknet_leaf_23_wb_clk_i cpu.timer_capture\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_20_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10395_ _00334_ clknet_leaf_8_wb_clk_i cpu.toggle_ctr\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_75_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07158__I _01429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07576__A4 _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07094__S _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05406__I _00917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05511__A3 _01018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05370_ cpu.regs\[12\]\[0\] cpu.regs\[13\]\[0\] cpu.regs\[14\]\[0\] cpu.regs\[15\]\[0\]
+ _00878_ _00879_ _00882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
Xclkbuf_leaf_35_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_35_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_83_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08452__I cpu.PC\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07040_ _00740_ _02530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06224__A1 cpu.timer_capture\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10020__A2 _04180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08991_ _03552_ _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07942_ _00947_ _03242_ _03249_ _03250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07873_ cpu.spi.div_counter\[2\] cpu.spi.divisor\[2\] _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09612_ _02473_ _04644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06824_ _02304_ _02321_ _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07724__A1 _02378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09543_ _04576_ _04577_ _04578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05316__I _00570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06755_ _02250_ _02251_ _02252_ _02253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05706_ cpu.PORTA_DDR\[0\] net79 _01211_ _01212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_93_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09474_ _04488_ _04492_ _04510_ _04511_ _04512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06686_ _02147_ _02148_ _02181_ _02184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__07531__I _02933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08425_ _03609_ _03630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05637_ _01142_ _01128_ _01143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_108_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08356_ _00673_ _03577_ _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_46_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05568_ _01060_ _01074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07307_ _02757_ _00068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08287_ _02841_ _03519_ _03523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05499_ _00654_ _01005_ _01006_ _01007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07238_ _02676_ _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05266__A2 cpu.ROM_spi_mode vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07169_ _00947_ _02644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10180_ _00119_ clknet_leaf_122_wb_clk_i cpu.regs\[11\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06610__I _00850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09165__B1 _02109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07715__A1 cpu.regs\[3\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08272__I _03510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10516_ _00454_ clknet_leaf_87_wb_clk_i cpu.ROM_addr_buff\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10447_ _00386_ clknet_leaf_25_wb_clk_i cpu.timer\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07403__B1 _02629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10378_ _00317_ clknet_leaf_89_wb_clk_i cpu.orig_PC\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07616__I _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07706__A1 _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09831__I _04813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06540_ cpu.startup_cycle\[1\] _02038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_88_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06471_ _01962_ _01202_ _01968_ _01969_ _01503_ _01970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_87_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08210_ _03246_ _03467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05422_ _00896_ _00931_ _00932_ _00933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_117_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09190_ _00949_ _04235_ _04236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08141_ cpu.uart.div_counter\[9\] _03407_ _03401_ _03411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_99_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05353_ _00864_ _00865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08072_ _03122_ _03354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05099__I2 cpu.regs\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05284_ _00816_ _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07023_ _00733_ _02516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_12_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08974_ _01077_ _04038_ _04060_ _04050_ _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07925_ cpu.spi.data_out_buff\[0\] _03234_ _03235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_89_Right_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05420__A2 _00930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07856_ _03157_ _03158_ _03169_ _03176_ _03177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input18_I io_in[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07787_ _03106_ _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06807_ _02294_ _02290_ _02295_ _02305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_94_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09526_ _04488_ _04547_ _04561_ _04511_ _04562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05490__B _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06920__A2 _01997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06738_ cpu.regs\[1\]\[5\] _00892_ _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09457_ cpu.PC\[7\] _01036_ _04495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_38_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09870__A1 net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_98_Right_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08408_ _02797_ _03598_ _03617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06669_ _00801_ _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09388_ _02361_ _04334_ _04428_ _04429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_50_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08339_ _03553_ _03564_ _00293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06436__A1 _01465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10301_ _00240_ clknet_leaf_42_wb_clk_i cpu.uart.div_counter\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09916__I _03236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07936__A1 _00922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10232_ _00171_ clknet_leaf_107_wb_clk_i cpu.regs\[4\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06295__S0 _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10163_ _00102_ clknet_leaf_123_wb_clk_i cpu.regs\[13\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05411__A2 _00896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06340__I _00614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10094_ _00037_ clknet_leaf_106_wb_clk_i cpu.br_rel_dest\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09651__I _02771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07711__I1 cpu.regs\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_94_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07547__S _02933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07710_ _03046_ _00182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05971_ _00818_ _01345_ _01476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08690_ _02665_ _03824_ _03829_ _03827_ _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_79_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07641_ _02988_ _03001_ _03004_ _00155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07572_ _01102_ _01297_ _01390_ _02960_ _02961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_TAPCELL_ROW_0_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_50_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_50_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_76_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09311_ _04042_ _04354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06523_ _01926_ _02008_ _01999_ _02022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09852__A1 _04819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08905__I _04000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09242_ _00768_ _04284_ _04286_ _04249_ _04287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06454_ _00659_ _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_29_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06385_ net66 _01089_ _01885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09604__A1 _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09173_ cpu.orig_flags\[1\] _04209_ _04180_ _01540_ _04219_ _04220_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_8_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05405_ _00909_ _00916_ _00917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08124_ _03331_ _03394_ _03397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08126__B _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05336_ cpu.PORTB_DDR\[5\] net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_0_71_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08055_ cpu.uart.data_buff\[0\] _03340_ _03341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05267_ cpu.regs\[1\]\[0\] _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07006_ cpu.ROM_addr_buff\[11\] _02481_ _02480_ _02500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05198_ cpu.IE cpu.needs_interrupt _00704_ _00735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput39 net39 io_oeb[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07918__A1 _03227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08957_ cpu.orig_IO_addr_buff\[0\] _04044_ _04045_ _01022_ _04046_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07908_ net70 _03220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08888_ cpu.timer_div\[5\] _03972_ _03986_ _03988_ _03989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07839_ cpu.timer_top\[2\] _02690_ _02683_ cpu.timer_top\[1\] _03160_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_55_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07146__A2 _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_38_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09843__A1 _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09509_ _03077_ _04349_ _04545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_117_Right_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_117_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10215_ _00154_ clknet_leaf_13_wb_clk_i cpu.regs\[6\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07166__I _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10146_ _00085_ clknet_leaf_105_wb_clk_i _00003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_77_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10077_ _00020_ clknet_leaf_118_wb_clk_i cpu.regs\[9\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06896__A1 _02393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05414__I _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06648__A1 _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_96_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06170_ _01454_ _01657_ _01672_ _01673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05121_ _00659_ cpu.br_rel_dest\[6\] cpu.br_rel_dest\[4\] _00660_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_41_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08460__I _03653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05052_ _00585_ _00594_ _00595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05623__A2 _01127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09860_ _04010_ _04842_ _04851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08811_ _03171_ _03928_ _03929_ _03931_ _03932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_09791_ cpu.pwm_top\[7\] cpu.pwm_counter\[7\] _04795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08742_ _02714_ _03865_ _03871_ _03873_ _03856_ _03874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05954_ _01450_ _01452_ _01458_ _01459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_108_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08673_ cpu.timer_top\[8\] _03818_ _03819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09291__I _04252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05885_ _01389_ _01390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_07624_ _02992_ _02985_ _02993_ _00149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09825__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07555_ cpu.regs\[10\]\[0\] _02951_ _02952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06506_ _01992_ _02001_ _02004_ _02005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07486_ _01374_ _02904_ _02906_ _00098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09225_ _00770_ _04264_ _04270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06437_ _01935_ _01936_ _01937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_60_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06368_ _01847_ _01849_ _01868_ _01869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09156_ _01598_ _01697_ _01784_ _04202_ _04203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_31_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08107_ cpu.uart.div_counter\[2\] cpu.uart.div_counter\[1\] cpu.uart.div_counter\[0\]
+ _03384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09087_ cpu.ROM_addr_buff\[2\] _04145_ _04148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06299_ _01799_ _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05319_ cpu.regs\[1\]\[3\] _00849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_101_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08038_ cpu.uart.div_counter\[12\] _03324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05614__A2 _00754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06811__A1 _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_111_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10000_ _00697_ _04963_ _02499_ _04964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09989_ _02454_ _04911_ _04954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05473__S1 _00977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06327__B1 _01266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07650__S _02999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09816__A1 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09150__B _00714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05409__I _00920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07358__A2 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05369__A1 _00006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10129_ _00072_ clknet_leaf_12_wb_clk_i cpu.toggle_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05670_ _00647_ _00648_ _01176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_9_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07340_ cpu.PC\[0\] _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07669__I0 _03007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07271_ _02726_ _02729_ _02731_ _00791_ _00058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09010_ _00865_ _04084_ _04088_ _04089_ _04090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_5_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06097__A2 _01547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06222_ cpu.timer_div\[4\] _01631_ _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06153_ _01654_ _00972_ _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08794__A1 cpu.timer_capture\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05104_ _00623_ _00643_ _00644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08123__C _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06084_ _01572_ _01573_ _01587_ _01588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09912_ _04815_ _04889_ _04890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05035_ cpu.regs\[8\]\[4\] cpu.regs\[9\]\[4\] cpu.regs\[10\]\[4\] cpu.regs\[11\]\[4\]
+ _00572_ _00576_ _00578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05319__I cpu.regs\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09843_ _04837_ _04829_ _04838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09774_ cpu.ROM_spi_cycle\[4\] _00666_ _04781_ _04783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06986_ _02474_ _02479_ _02480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06309__B1 _01807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08725_ _03857_ _03859_ _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05937_ _01441_ _01442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08656_ _03802_ _03806_ _00368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05054__I _00596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05868_ _01373_ _01374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08587_ _03729_ _03757_ _00348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07607_ _01372_ _02980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07538_ cpu.regs\[11\]\[3\] _02934_ _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05799_ _01148_ _01305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__05989__I _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07285__A1 _02653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07469_ cpu.regs\[14\]\[2\] _02893_ _02896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10480_ _00419_ clknet_leaf_20_wb_clk_i cpu.timer_div\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09208_ _02783_ _04253_ _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09139_ _02647_ _04186_ _04187_ _04188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_114_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_107_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_107_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08275__I _03495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06009__B _01215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07619__I _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06840_ _02332_ _02337_ _02338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07751__A2 _03064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06771_ _02266_ _02268_ _02269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05722_ _01193_ _01226_ _01227_ _01228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08510_ cpu.toggle_ctr\[15\] _03693_ _03696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09490_ _03076_ _00864_ _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_81_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08441_ _03077_ _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07503__A2 _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05653_ cpu.br_rel_dest\[2\] _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05584_ _01089_ _01090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08372_ cpu.orig_IO_addr_buff\[4\] _03587_ _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_58_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07267__A1 _01243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07323_ _02769_ _02763_ _02770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07254_ _02714_ _02703_ _02716_ _02717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06205_ _01706_ _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_103_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07185_ _01707_ _02657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_76_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07529__I _02933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06136_ _01246_ _01639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06067_ _01446_ _01570_ _01571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09744__I _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09826_ _04825_ _00519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05428__S1 _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09757_ _04755_ _04770_ _04771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06969_ _00662_ _02463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_100_Left_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_5_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_5_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_96_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08708_ _03835_ _03845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09688_ _04709_ _04712_ _04713_ _00493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_69_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08639_ cpu.pwm_top\[5\] _03787_ _03793_ _03795_ _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05512__I _01019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10601_ _00539_ clknet_leaf_62_wb_clk_i cpu.PORTB_DDR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10532_ _00470_ clknet_leaf_88_wb_clk_i cpu.TIE vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08823__I _03918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10463_ _00402_ clknet_leaf_22_wb_clk_i cpu.timer_capture\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10394_ _00333_ clknet_leaf_7_wb_clk_i cpu.toggle_ctr\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07430__B2 _01612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09183__A1 _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07174__I _02647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06792__I0 _00917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09238__A2 _04281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07249__A1 cpu.timer_capture\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08997__B2 _02722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_75_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_75_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_70_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07421__A1 _02853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07793__B _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08990_ _04055_ _04073_ _00435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07941_ cpu.spi.data_out_buff\[1\] _03243_ _03249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07872_ cpu.spi.divisor\[6\] _03192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09611_ _04642_ _04643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06823_ _02315_ _02320_ _02321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09542_ cpu.PC\[11\] _00951_ _04577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06754_ _02248_ _02249_ _02252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05705_ _01210_ _01211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_78_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09473_ _04330_ _04511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06685_ _02181_ _02182_ _02183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08424_ cpu.orig_PC\[5\] _03628_ _03629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05636_ _01036_ _01142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08355_ _00727_ _03576_ _03577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05567_ _00647_ _01073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_116_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08988__A1 _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07306_ cpu.toggle_top\[10\] _02749_ _02755_ _02756_ _02757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_34_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08286_ _00792_ _03522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05498_ _00990_ _01000_ _01006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07237_ cpu.timer\[4\] _02702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_14_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07168_ _02641_ _02634_ _02643_ _00791_ _00043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07259__I _01997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06119_ net9 _01517_ _01207_ _01622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07099_ _02379_ _02380_ _02386_ _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__05974__A1 _00991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09165__B2 _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09809_ _04810_ _04811_ _00516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_70_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05041__I3 cpu.regs\[7\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09640__A2 cpu.ROM_addr_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10515_ _00453_ clknet_leaf_80_wb_clk_i cpu.ROM_addr_buff\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07169__I _00947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10446_ _00385_ clknet_leaf_26_wb_clk_i cpu.timer\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10377_ _00316_ clknet_leaf_86_wb_clk_i cpu.orig_PC\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_122_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_122_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06390__A1 cpu.uart.divisor\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06470_ net14 _01206_ _01208_ _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__06142__A1 _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05152__I _00689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05421_ _00864_ _00930_ _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08140_ _03407_ _03401_ _03410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05352_ _00863_ _00864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08071_ _03347_ _03351_ _03353_ _00235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05099__I3 cpu.regs\[3\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05283_ _00810_ _00815_ _00816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_113_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07022_ _02513_ _02515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07079__I _02541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08973_ _01161_ _04039_ _04041_ _04058_ _04059_ _04060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__05500__S0 _00887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07924_ _03233_ _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09147__A1 _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07855_ _03140_ _03153_ _03173_ _03175_ _03176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_TAPCELL_ROW_108_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07786_ cpu.spi.data_in_buff\[3\] _03102_ _03112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06806_ _02292_ _02303_ _02304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09525_ _04558_ _04560_ _04561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06737_ _02212_ _02231_ _02235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_94_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06133__A1 cpu.timer_capture\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09456_ _04353_ _04492_ _04493_ _04397_ _04494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06668_ _02137_ _02165_ _02166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08407_ _03614_ _03592_ _03615_ _03616_ _00309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05619_ _01121_ _01123_ _01124_ _01125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_108_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09387_ _04335_ _04412_ _04428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06599_ _02096_ _02097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_22_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08338_ cpu.uart.receive_div_counter\[13\] _03547_ _03561_ _03563_ _03564_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08269_ _03307_ _03507_ _03508_ _00279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10300_ _00239_ clknet_leaf_53_wb_clk_i cpu.uart.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_61_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10231_ _00170_ clknet_leaf_107_wb_clk_i cpu.regs\[4\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06295__S1 _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10162_ _00101_ clknet_leaf_0_wb_clk_i cpu.regs\[13\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_67_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05411__A3 _00922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10093_ _00036_ clknet_leaf_102_wb_clk_i cpu.br_rel_dest\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07653__S _02999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06372__A1 _01833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05700__I _01205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_94_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10429_ _00368_ clknet_leaf_27_wb_clk_i cpu.timer_div_counter\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05970_ _01449_ _01443_ _01459_ _01474_ _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__09842__I _02668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08352__A2 _03574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07640_ cpu.regs\[6\]\[1\] _03002_ _03004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06363__A1 _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07571_ _01084_ _01169_ _01431_ _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_0_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09310_ _04033_ _04353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06522_ _02010_ _02012_ _02020_ _02021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__06115__A1 net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09241_ _04253_ _04265_ _04285_ _04286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06453_ _01952_ _00019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06384_ net46 _01616_ _01882_ _01883_ _01514_ _01884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_103_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_90_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_90_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09289__I _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05404_ _00911_ _00915_ _00916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09172_ _04211_ _04212_ _04214_ _04218_ _04219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_08123_ _03393_ _03389_ _03396_ _03306_ _00245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05335_ cpu.PORTA_DDR\[4\] net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__07030__C _02522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08054_ _03339_ _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07005_ _02045_ _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08921__I _01005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05266_ _00799_ cpu.ROM_spi_mode net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__07091__A2 _02572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_101_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05197_ _00701_ net18 _00734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_3_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08040__B2 cpu.uart.divisor\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input30_I sram_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08956_ _04034_ _04045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07473__S _02891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08887_ _03987_ _03988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07907_ _03203_ _03219_ _00206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_98_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07838_ cpu.timer_top\[1\] _02684_ _02675_ cpu.timer_top\[0\] _03159_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08368__I _03586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09540__A1 _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07272__I _00922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07769_ cpu.spi.counter\[3\] _03098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09508_ _03641_ _04520_ _04544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09439_ _04294_ _04463_ _04477_ _04331_ _04478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_54_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10214_ _00153_ clknet_leaf_116_wb_clk_i cpu.regs\[7\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10145_ _00084_ clknet_leaf_105_wb_clk_i _00002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10076_ _00019_ clknet_leaf_120_wb_clk_i cpu.regs\[9\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_4_10_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05699__A3 _01204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06896__A2 _02391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07845__A1 _01879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05120_ cpu.br_rel_dest\[7\] _00659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_4_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05051_ _00587_ _00592_ _00593_ _00594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08810_ _02642_ _03930_ _03931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09790_ cpu.pwm_top\[4\] cpu.pwm_counter\[4\] _04794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06584__A1 _00590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08741_ _03832_ _03872_ _03873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05953_ _01454_ _01455_ _01457_ _01458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05884_ _01216_ _01389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08672_ _03816_ _03818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07623_ cpu.regs\[7\]\[3\] _02984_ _02993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_105_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08916__I _02647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08089__A1 _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07554_ _02948_ _02951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06505_ _01992_ _02003_ _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07485_ cpu.regs\[13\]\[0\] _02905_ _02906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09224_ _04268_ _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06436_ _01465_ _01911_ _01936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05340__I cpu.PORTB_DDR\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06367_ _01853_ _01856_ _01857_ _01331_ _01867_ _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_16_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09155_ _01367_ _01489_ _04199_ _04202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_32_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08106_ _03369_ _03383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09086_ _03360_ _04146_ _04147_ _00457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06298_ _00960_ _01794_ _01798_ _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05318_ cpu.regs\[4\]\[3\] cpu.regs\[5\]\[3\] cpu.regs\[6\]\[3\] cpu.regs\[7\]\[3\]
+ _00846_ _00847_ _00848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08037_ _03315_ _03317_ _03319_ _03322_ _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
X_05249_ _00730_ _00783_ _00784_ cpu.instr_cycle\[3\] _00785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_3_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09988_ _02449_ _04704_ _02461_ _04952_ _04953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08939_ _04027_ _04028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_99_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06327__B2 _01004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06327__A1 _01121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05515__I _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06566__A1 _02062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10128_ _00071_ clknet_leaf_12_wb_clk_i cpu.toggle_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10059_ _01602_ _05013_ _05017_ _00560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_38_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_29_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_29_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08736__I _03121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07270_ cpu.timer_top\[0\] _02730_ _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06221_ _01709_ _01611_ _01721_ _01722_ _01631_ _01723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_72_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06152_ _01446_ _01570_ _01655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_111_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05103_ cpu.regs\[8\]\[7\] cpu.regs\[9\]\[7\] cpu.regs\[10\]\[7\] cpu.regs\[11\]\[7\]
+ _00633_ _00634_ _00643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06083_ _01152_ _01562_ _01578_ _01462_ _01586_ _01587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10050__A1 _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09911_ _04887_ _04889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05034_ cpu.regs\[12\]\[4\] cpu.regs\[13\]\[4\] cpu.regs\[14\]\[4\] cpu.regs\[15\]\[4\]
+ _00572_ _00576_ _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_111_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09842_ _02668_ _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_13_Left_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_111_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09773_ _04781_ _04782_ _00509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06985_ _02472_ _02466_ _02468_ _02059_ _02479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_08724_ cpu.timer_capture\[3\] _03858_ _03529_ _03859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06309__A1 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05335__I cpu.PORTA_DDR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05936_ _00831_ _00918_ _01441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08655_ cpu.timer_div_counter\[3\] _03804_ _03806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05867_ _01372_ _01373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08586_ cpu.toggle_ctr\[14\] _03755_ cpu.toggle_ctr\[15\] _03757_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07606_ _02930_ _02971_ _02979_ _00145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07809__A1 cpu.timer_div\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05798_ _01131_ _01304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07537_ _02923_ _02935_ _02939_ _00116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Left_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07468_ _01495_ _02892_ _02895_ _00091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07399_ cpu.uart.receive_div_counter\[7\] _02832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_106_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09207_ _04252_ _04253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06419_ _01437_ _01918_ _01919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09138_ cpu.orig_flags\[3\] _04186_ _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09477__I _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07037__A2 _02527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06096__I0 net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10041__A1 _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09069_ _04132_ cpu.ROM_addr_buff\[13\] _04126_ _04133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_31_Left_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output61_I net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09940__I _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_43_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08473__A1 _02758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09973__A1 cpu.ROM_addr_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08776__A2 _03811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08528__A2 cpu.toggle_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06003__A3 _01063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07635__I _02999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06770_ _02264_ _00917_ _02267_ _02268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05721_ cpu.uart.busy _01100_ _01191_ _01227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08440_ cpu.orig_PC\[10\] _03640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05652_ _00720_ _01156_ _01157_ _01158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_86_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05583_ _01088_ _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08371_ _03579_ _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_85_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07322_ _02715_ _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07253_ _02697_ _02715_ _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07184_ _02656_ _00046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_83_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06204_ _00960_ _01013_ _01705_ _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_5_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09964__A1 net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06135_ cpu.timer_capture\[11\] _01242_ _01635_ _01637_ _01244_ _01638_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_60_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09964__B2 _04931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06066_ _01554_ _01562_ _01569_ _01570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_111_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09825_ net61 _04814_ _04824_ _04821_ _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09756_ cpu.ROM_spi_dat_out\[3\] _04715_ _04762_ _04770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06968_ cpu.startup_cycle\[2\] _02462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__06950__A1 _02031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09687_ _00790_ _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08707_ cpu.timer\[1\] _03838_ _03844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05919_ _01421_ _01422_ _01423_ _01424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08638_ _03794_ _03795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06899_ net1 _02075_ _02396_ _02397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08569_ _03727_ _03746_ _00341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_37_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10600_ _00538_ clknet_leaf_62_wb_clk_i cpu.PORTB_DDR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10531_ _00469_ clknet_leaf_78_wb_clk_i cpu.last_addr\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_40_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10462_ _00401_ clknet_leaf_8_wb_clk_i cpu.timer_capture\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10393_ _00332_ clknet_leaf_13_wb_clk_i cpu.toggle_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_20_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05292__I1 _00822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09183__A2 _04205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08286__I _00792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07190__I _02661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06534__I _02032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07421__A2 cpu.uart.receive_div_counter\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_7_0_wb_clk_i clknet_0_wb_clk_i clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_50_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07940_ _03248_ _00210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_44_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_44_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07871_ _03185_ _03186_ _03189_ _03190_ _03191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_09610_ _04641_ _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06822_ _02317_ _02319_ _02320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09580__I _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09541_ _03089_ _00951_ _04576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06753_ _02242_ _02243_ _02251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05704_ _01043_ _01046_ _01062_ _01210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_09472_ _04494_ _04509_ _04510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06684_ _02147_ _02148_ _02182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08423_ _03595_ _03628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05635_ _01139_ _01140_ _00992_ _01141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08354_ cpu.instr_cycle\[3\] cpu.instr_cycle\[1\] _03576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05566_ _00680_ _01067_ _01068_ _01070_ _01071_ _01072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__08437__A1 _03637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07305_ _02661_ _02756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08285_ _03517_ _03518_ _03521_ _03414_ _00282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05497_ _01004_ _01005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_27_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07236_ _02673_ _02701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07167_ _02642_ _02637_ _02643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09937__A1 _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06118_ net24 _01389_ _01618_ _01620_ _01109_ _01621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_42_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07098_ _02534_ _02344_ _02582_ _02583_ _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06049_ _01324_ _01314_ _01553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_100_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09165__A2 _02185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09808_ _03738_ _00744_ _04811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_70_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09739_ _04755_ _04756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06923__A1 _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_15_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08676__A1 cpu.timer_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07479__A2 _02891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05034__S0 _00572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10514_ _00452_ clknet_leaf_80_wb_clk_i cpu.ROM_addr_buff\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09928__A1 cpu.PORTA_DDR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10445_ _00384_ clknet_leaf_26_wb_clk_i cpu.timer\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07403__A2 _02641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10376_ _00315_ clknet_leaf_86_wb_clk_i cpu.orig_PC\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07185__I _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07167__A1 _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05273__S0 _00803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08419__A1 _02561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05420_ _00864_ _00930_ _00931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05351_ _00862_ _00863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_114_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08070_ _03100_ _03352_ _03348_ _03353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05282_ _00812_ _00814_ _00815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07642__A2 _03002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09919__A1 _04823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07021_ _02513_ _02514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09395__A2 cpu.br_rel_dest\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08972_ _04031_ _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05500__S1 _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07095__I _02581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07923_ _03229_ _03231_ _03232_ _03233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07854_ _03145_ _03174_ _03156_ _03158_ _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07823__I cpu.timer_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06805_ _02297_ _02298_ _02303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07785_ _01528_ _03107_ _03111_ _00192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05184__A3 _00720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05343__I cpu.PORTA_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09524_ _03640_ _04281_ _04559_ _04397_ _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06736_ _02204_ _02233_ _02234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09455_ cpu.orig_PC\[8\] _04354_ _04493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06667_ _02162_ _02164_ _02165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05618_ _01117_ _01087_ _01124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08406_ _03413_ _03616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07330__A1 _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09386_ _04347_ _04412_ _04426_ _04373_ _04427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06375__S _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06598_ _02090_ _02095_ _02096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_22_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08337_ _03513_ _03562_ _03563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05549_ _00678_ _01055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_62_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08268_ _02884_ _03503_ _03508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07633__A2 _02986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07219_ _02661_ _02687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08199_ _00728_ _03366_ _03367_ _03456_ _03457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_10230_ _00169_ clknet_leaf_116_wb_clk_i cpu.regs\[5\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_72_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09418__C _04340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Left_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10161_ _00100_ clknet_leaf_0_wb_clk_i cpu.regs\[13\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07149__A1 _02626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10092_ _00035_ clknet_leaf_102_wb_clk_i cpu.br_rel_dest\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08897__A1 _02626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06372__A2 _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05253__I _00788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05883__A1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08821__A1 cpu.timer_capture\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07624__A2 _02985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05635__A1 _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07908__I net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10428_ _00367_ clknet_leaf_27_wb_clk_i cpu.timer_div_counter\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_94_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10359_ _00298_ clknet_leaf_55_wb_clk_i cpu.orig_IO_addr_buff\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08888__A1 cpu.timer_div\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_69_Left_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07570_ _02930_ _02951_ _02959_ _00129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09998__C _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05163__I _00700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06521_ _01466_ _02003_ _02014_ _01484_ _02019_ _02020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_118_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09240_ _02792_ _04252_ _04285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06452_ _01951_ cpu.regs\[9\]\[6\] _01166_ _01952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06383_ net57 _01615_ _01616_ _01883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_103_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08407__C _03616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05403_ _00905_ _00912_ _00914_ _00915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09171_ _04215_ _04216_ _04217_ _04218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_113_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08122_ cpu.uart.div_counter\[5\] _03383_ _03395_ _03396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05334_ cpu.PORTB_DDR\[4\] net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XANTENNA__08812__A1 cpu.timer_capture\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07615__A2 _02985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08053_ _03323_ _03338_ _03339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_78_Left_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05626__A1 _01131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07004_ cpu.ROM_spi_dat_out\[7\] _02497_ _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05265_ net75 _00799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_113_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05196_ _00671_ _00733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09238__C _00761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05641__A4 _01126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09368__A2 _04408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08955_ _04043_ _04044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07906_ cpu.spi.div_counter\[7\] _03218_ _03219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input23_I io_in[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08886_ _02771_ _03987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08879__A1 cpu.timer_div\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07837_ _03155_ cpu.timer\[15\] _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07551__A1 _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07768_ cpu.spi.data_in_buff\[0\] _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_55_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09507_ _04521_ _04543_ _04484_ _00482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06719_ _00820_ _01014_ _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05073__I _00614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07699_ _03039_ _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_109_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09438_ _04470_ _04474_ _04476_ _04477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09369_ _02782_ _02386_ _04410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output91_I net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10213_ _00152_ clknet_leaf_115_wb_clk_i cpu.regs\[7\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06042__A1 _00794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10144_ _00083_ clknet_leaf_16_wb_clk_i _00001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10075_ _00018_ clknet_leaf_122_wb_clk_i cpu.regs\[9\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07463__I _02891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xwrapped_qcpu_110 io_out[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_69_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05711__I _01216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08294__I _03236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08270__A2 _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06281__B2 _01332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06281__A1 _01326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05050_ _00003_ _00593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_111_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06033__A1 _01498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07081__I0 _02361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06584__A2 _01996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08740_ _02707_ _03860_ _02714_ _03872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05952_ _00920_ _01353_ _01456_ _01341_ _01355_ _01457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_108_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05883_ net60 _01090_ _01388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08671_ _03816_ _03817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07622_ _01699_ _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10013__B _04340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07553_ _02949_ _02950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07484_ _02902_ _02905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06504_ _01990_ _02002_ _02003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09223_ _00778_ _00741_ _04268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06435_ _01340_ _01912_ _01915_ _01451_ _01934_ _01935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_32_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_86_Left_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_60_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09154_ _01923_ _01999_ _04199_ _04200_ _04201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_08105_ cpu.uart.div_counter\[1\] _03365_ _03382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06366_ _01579_ _01844_ _01862_ _01866_ _01867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_16_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09085_ cpu.last_addr\[1\] _04143_ _04147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06297_ _00967_ _01797_ _01798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05317_ _00805_ _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_32_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08036_ cpu.uart.div_counter\[5\] _01804_ _02848_ cpu.uart.div_counter\[2\] _03321_
+ _03322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_05248_ cpu.instr_cycle\[1\] _00784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05179_ cpu.base_address\[0\] _00716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09987_ _02459_ _04951_ _04952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_95_Left_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08379__I _03595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08938_ _01149_ _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_4_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08869_ cpu.timer_div\[0\] _03972_ _03974_ _03975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09003__I _04083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05531__I _00754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05838__A1 _00891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06015__A1 net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06566__A2 _02063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10127_ _00070_ clknet_leaf_12_wb_clk_i cpu.toggle_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07193__I _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10058_ cpu.regs\[15\]\[2\] _05014_ _05017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07126__C _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_69_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_69_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_46_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05829__A1 _00863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09848__I _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06220_ cpu.spi.divisor\[4\] _01628_ _01188_ _01722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_109_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08243__A2 _03368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06151_ _00859_ _01654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_14_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06254__A1 _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05102_ _00587_ _00641_ _00642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06082_ _01579_ _01568_ _01583_ _01585_ _01586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__10050__A2 _02932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09910_ _04887_ _04888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05033_ _00575_ _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_95_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09841_ _04836_ _00523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_95_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09772_ cpu.ROM_spi_cycle\[0\] _04749_ _03897_ _04782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06984_ _02471_ _02474_ _02477_ _02478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_08723_ _03845_ _03858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05935_ _01438_ _01439_ _01440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_96_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08654_ _03801_ _03804_ _03805_ _00367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05866_ _01308_ _01371_ _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_48_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08585_ _03729_ _03756_ _00347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07605_ cpu.regs\[8\]\[7\] _02969_ _02979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05797_ _01299_ _01301_ _01302_ _01303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07536_ cpu.regs\[11\]\[2\] _02936_ _02939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09206_ _01347_ _01020_ _01548_ _04252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_07467_ cpu.regs\[14\]\[1\] _02893_ _02895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07398_ cpu.uart.divisor\[13\] _02829_ _02830_ _02824_ _02831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06418_ _01915_ _01917_ _01918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09137_ _04180_ _04186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06349_ _01837_ _01850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09068_ cpu.regs\[3\]\[5\] _03649_ _04101_ _04132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06245__B2 _01452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08019_ _03304_ _03298_ _03305_ _03306_ _00231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_102_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09034__I1 cpu.ROM_addr_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output54_I net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06484__A1 cpu.toggle_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06293__S _00885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06236__A1 _01704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_116_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_116_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07916__I _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09336__C _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05436__I _00946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05720_ _01195_ _01224_ _01225_ _01226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_81_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05651_ _00738_ _00780_ _00685_ _01091_ _01157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_105_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08370_ _01078_ _03580_ _03588_ _03583_ _00300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_85_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05582_ _01044_ _01047_ _01087_ _01088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_07321_ _02768_ _00071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09661__A1 _00746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06475__A1 cpu.spi.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07252_ _01801_ _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07183_ cpu.uart.divisor\[4\] _02651_ _02655_ _02639_ _02656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06203_ _00967_ _01010_ _01705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06134_ _01241_ _01636_ _01637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06227__A1 cpu.timer_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06065_ _01553_ _01568_ _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_47_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09246__C _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07826__I cpu.timer_top\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09824_ _04823_ _04816_ _04824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07727__A1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09755_ _04756_ _04768_ _04769_ _00504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06967_ _02458_ _02461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09686_ _02039_ _04711_ _04712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08706_ _03835_ _03843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05918_ _01275_ _01423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06898_ _02373_ _02395_ _02075_ _02396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_68_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08637_ _02771_ _03794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05849_ _00720_ _01355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_64_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08568_ _03715_ _03744_ _03746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08499_ cpu.toggle_ctr\[11\] _03685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07519_ _02927_ _00110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06466__A1 cpu.PORTB_DDR\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10530_ _00468_ clknet_leaf_78_wb_clk_i cpu.last_addr\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_86_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10461_ _00400_ clknet_leaf_9_wb_clk_i cpu.timer_capture\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_45_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10392_ _00331_ clknet_leaf_14_wb_clk_i cpu.toggle_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_20_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05292__I2 _00823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07718__A1 _00787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06288__S _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06941__A2 _02407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09891__A1 _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08516__B _01170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06209__A1 cpu.PORTA_DDR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09946__A2 _00733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07646__I _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07870_ cpu.spi.div_counter\[7\] cpu.spi.divisor\[7\] _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06821_ _02309_ _02318_ _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_84_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_84_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08477__I _03653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_50_Left_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09540_ _00949_ _04505_ _04574_ _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06752_ _02248_ _02249_ _02250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05703_ _01203_ _01206_ _01208_ _01209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09471_ _04502_ _04504_ _04508_ _04370_ _04509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
Xclkbuf_leaf_13_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_13_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08422_ _02563_ _03619_ _03627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06683_ _02178_ _02179_ _02180_ _02181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_65_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05499__A2 _01005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_120_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06696__A1 _00605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05634_ _01127_ _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08353_ _03573_ _00703_ _03575_ _00296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_74_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05565_ _01065_ _01071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08284_ _02849_ _03510_ _03519_ _03520_ _03521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08988__A3 _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07304_ _02754_ _02750_ _02755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06448__A1 net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08145__C _03414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07235_ _02700_ _00053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05496_ _01003_ _01004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_81_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07166_ _01540_ _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08940__I _04028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_3_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06117_ _01217_ _01619_ _01620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07097_ net20 _02036_ _02583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06048_ _01325_ _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_100_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05076__I _00572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07999_ cpu.uart.dout\[1\] _03289_ _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09704__C _04684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06384__B1 _01882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09807_ _00737_ _00743_ net89 _04810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05187__A1 cpu.uart.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09738_ _04750_ _04755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_69_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09669_ _02483_ _04696_ _04697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05034__S1 _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06439__A1 _01360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10513_ _00451_ clknet_leaf_80_wb_clk_i cpu.ROM_addr_buff\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10444_ _00383_ clknet_leaf_29_wb_clk_i cpu.timer\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07939__B2 _03247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10375_ _00314_ clknet_leaf_87_wb_clk_i cpu.orig_PC\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09156__A3 _01784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_88_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05273__S1 _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05350_ _00715_ _00862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_112_Right_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_99_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05281_ _00586_ _00813_ _00593_ _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_113_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07020_ _02511_ _02512_ _02513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_23_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08971_ cpu.orig_IO_addr_buff\[2\] _04056_ _04057_ _02692_ _04058_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07922_ _02519_ _03232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08355__A1 _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07853_ cpu.timer\[8\] _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06804_ _02286_ _02301_ _02302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_07784_ cpu.spi.data_in_buff\[2\] _03108_ _03109_ _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_108_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09523_ _04281_ _04546_ _04559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06735_ _02212_ _02231_ _02232_ _02233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09454_ _04491_ _04492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06666_ _02140_ _02163_ _02164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05617_ _01117_ _01122_ _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08405_ cpu.orig_PC\[0\] _03611_ _03615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09385_ _04423_ _04425_ _04426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08336_ _02829_ _03557_ _03562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06597_ _02093_ _02094_ _02095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_22_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05548_ _01045_ _01054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_50_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08267_ _03226_ _02884_ _03496_ _03507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_61_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05479_ _00987_ _00988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07218_ _02684_ _02677_ _02678_ _02685_ _02686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08198_ _00767_ _03456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07149_ _02626_ _02620_ _02627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10160_ _00099_ clknet_leaf_2_wb_clk_i cpu.regs\[13\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10091_ _00034_ clknet_leaf_103_wb_clk_i cpu.br_rel_dest\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07149__A2 _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_76_Right_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_58_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05534__I _00756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09846__A1 _01063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_106_Left_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08845__I _03958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05883__A2 _01090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_85_Right_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05635__A2 _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10427_ _00366_ clknet_leaf_27_wb_clk_i cpu.timer_div_counter\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_115_Left_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10358_ _00297_ clknet_leaf_17_wb_clk_i cpu.orig_IO_addr_buff\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10289_ _00228_ clknet_leaf_45_wb_clk_i cpu.uart.dout\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06060__A2 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_94_Right_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06899__A1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09837__A1 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06520_ _01454_ _01998_ _02015_ _02018_ _02019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_06451_ _01950_ _01951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_113_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05402_ _00913_ _00914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06382_ cpu.PORTA_DDR\[6\] _01613_ _01882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_16_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09170_ _00590_ _02361_ _02416_ _02418_ _04217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_08121_ _03371_ _03394_ _03395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_98_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05333_ cpu.PORTA_DDR\[3\] net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_44_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07076__A1 _02561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08052_ _03327_ _03329_ _03334_ _03337_ _03338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_05264_ _00793_ _00798_ _00009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_71_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05626__A2 _01127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07003_ _02447_ _02497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_102_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05195_ _00700_ _00732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07379__A2 _02385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08954_ _04042_ _04043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06051__A2 _00944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07905_ cpu.spi.div_counter\[6\] _03216_ _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08885_ _02766_ _03983_ _03986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07836_ _03140_ _03154_ _03156_ _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input16_I io_in[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09828__A1 net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07551__A2 _02071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07767_ _03053_ _03095_ _03096_ _00189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_69_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09506_ _04487_ _04538_ _04539_ _04542_ _04049_ _04543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_06718_ _00834_ _00985_ _02216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07698_ _03038_ _03039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_109_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09437_ _04209_ _04463_ _04475_ _04327_ _04476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06649_ _02146_ _02145_ _02147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__05314__A1 _00566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09368_ _02548_ _04408_ _04409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08319_ _02862_ _03543_ _03544_ _03548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_09299_ _02810_ _04262_ _04343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07067__A1 _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05617__A2 _01122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06290__A2 _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10212_ _00151_ clknet_leaf_114_wb_clk_i cpu.regs\[7\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06042__A2 _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10143_ _00082_ clknet_leaf_105_wb_clk_i _00000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10074_ _00017_ clknet_leaf_122_wb_clk_i cpu.regs\[9\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09819__A1 _04819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_qcpu_100 io_oeb[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_qcpu_111 io_out[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_69_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06296__S _00870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06095__I _01157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input8_I io_in[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05951_ _00831_ _00919_ _01456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05882_ _01113_ _01384_ _01386_ _01387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_84_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08670_ _01111_ _02727_ _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08730__A1 cpu.timer_capture\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07621_ _02990_ _02985_ _02991_ _00148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_105_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07552_ _02948_ _02949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09286__A2 _03456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06503_ _00631_ _01840_ _02002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08418__C _03616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07483_ _02903_ _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09222_ _00739_ _04266_ _04267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06434_ _00656_ _01933_ _01934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06365_ _01451_ _01854_ _01863_ _01460_ _01865_ _01866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_09153_ _01745_ _01850_ _04200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08104_ _03375_ _03380_ _03381_ _00241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05316_ _00570_ _00846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_32_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09084_ cpu.ROM_addr_buff\[1\] _04145_ _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06296_ _01795_ _01796_ _00870_ _01797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08035_ _03320_ cpu.uart.divisor\[1\] _03316_ cpu.uart.div_counter\[0\] _03321_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05247_ _00750_ _00763_ _00768_ _00782_ _00783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_40_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07765__S _02401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05178_ cpu.base_address\[1\] _00715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09986_ _02457_ _04727_ _02456_ _04951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_4_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08937_ _04026_ _00429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08868_ _02726_ _03973_ _03974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07819_ _03138_ cpu.timer\[14\] cpu.timer\[13\] _03139_ _03140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_08799_ _01239_ _03921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08395__I _03595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08788__A1 cpu.timer_capture\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10126_ _00069_ clknet_leaf_11_wb_clk_i cpu.toggle_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07763__A2 _03092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10057_ _01494_ _05013_ _05016_ _00559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08712__A1 cpu.timer_capture\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05526__A1 _00656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07279__A1 _02644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_38_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_38_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_102_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06150_ _01378_ _01652_ _01653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_80_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05101_ cpu.regs\[12\]\[7\] cpu.regs\[13\]\[7\] cpu.regs\[14\]\[7\] cpu.regs\[15\]\[7\]
+ _00633_ _00634_ _00641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06081_ _01471_ _01584_ _01585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_37_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09864__I _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05169__I cpu.br_rel_dest\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05032_ _00574_ _00575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09840_ net66 _04828_ _04835_ _04833_ _04836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_1_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09771_ cpu.ROM_spi_cycle\[0\] _04749_ _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06983_ cpu.mem_cycle\[0\] _02054_ _02476_ _02477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__05765__A1 _01269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08722_ cpu.timer\[3\] _03850_ _03855_ _03834_ _03856_ _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05934_ cpu.br_rel_dest\[0\] _00818_ _01439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_37_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08653_ cpu.timer_div_counter\[0\] cpu.timer_div_counter\[1\] cpu.timer_div_counter\[2\]
+ _03805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05517__A1 _01020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05865_ _01309_ _01367_ _01369_ _01370_ _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_95_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07604_ _02978_ _00144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05632__I cpu.br_rel_dest\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05796_ _01140_ _01302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08584_ cpu.toggle_ctr\[14\] _03755_ _03756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_49_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07535_ _02921_ _02935_ _02938_ _00115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07466_ _01374_ _02892_ _02894_ _00090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09205_ _03456_ _04248_ _04250_ _04251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06417_ _01835_ _01916_ _01917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_17_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07397_ cpu.uart.receive_div_counter\[12\] _02830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_76_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09136_ cpu.TIE _04184_ _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06348_ _01326_ _01848_ _01849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09067_ _04131_ _00454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06279_ _01745_ _01779_ _01479_ _01781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08018_ _02617_ _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05079__I cpu.regs\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09195__A1 _01131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09969_ _04934_ _04935_ _04930_ _04936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_99_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09498__A2 _04033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output47_I net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09442__C _04340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09422__A2 _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08933__A1 _02847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10109_ _00052_ clknet_leaf_22_wb_clk_i cpu.timer_capture\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05650_ _01092_ _01156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_05581_ _01057_ _01086_ _01087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_58_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07320_ cpu.toggle_top\[13\] _02761_ _02767_ _02756_ _02768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_14_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07251_ cpu.timer\[6\] _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07182_ _02653_ _02654_ _02655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06202_ _01430_ _01704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_14_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06133_ cpu.timer_capture\[3\] _01236_ _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_113_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06064_ _01565_ _01567_ _01568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_22_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08924__A1 _02824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05738__A1 _01243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09823_ _00946_ _04823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09754_ cpu.ROM_spi_dat_out\[3\] _04760_ _03761_ _04769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06966_ _02456_ _02041_ _02458_ _02459_ _02460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__08938__I _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09685_ _04710_ _04711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08705_ _03839_ _03842_ _03646_ _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_69_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05917_ _01021_ _01268_ _01422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06897_ _02374_ _02392_ _02394_ _02395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_96_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08636_ _02766_ _03788_ _03793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05848_ _01345_ _01354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_64_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05910__A1 cpu.timer_top\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08567_ _03732_ _03744_ _03745_ _00340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05779_ _01279_ _01276_ _01285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_77_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08498_ cpu.toggle_ctr\[12\] _03684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07518_ _01789_ cpu.regs\[12\]\[4\] _02917_ _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_36_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07449_ cpu.uart.receive_counter\[2\] _02875_ _02880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_92_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10460_ _00399_ clknet_leaf_8_wb_clk_i cpu.timer_capture\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09119_ cpu.ROM_addr_buff\[11\] _04159_ _04171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10391_ _00330_ clknet_leaf_14_wb_clk_i cpu.toggle_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_20_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_75_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06921__I _00638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09168__B2 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05292__I3 cpu.regs\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09340__A1 _02561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06154__A1 net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07199__I _02668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10589_ _00527_ clknet_leaf_66_wb_clk_i net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07927__I _03236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09159__A1 _00997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08906__A1 _02636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05447__I _00956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06393__A1 cpu.spi.divisor\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06820_ _02309_ _02310_ _02311_ _02318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06751_ _02215_ _02218_ _02220_ _02249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_05702_ _01207_ _01208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_92_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09470_ _01020_ _04505_ _04507_ _04309_ _04508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_06682_ _00821_ _00835_ _00986_ _01016_ _02180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_08421_ _03625_ _03626_ _03610_ _00313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06145__B2 _00956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05633_ _01138_ _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_86_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_53_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_53_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08352_ cpu.had_int _03574_ cpu.needs_interrupt _03575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05564_ _01069_ _01051_ _01070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_74_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08283_ _02868_ _03520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07303_ _00946_ _02754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_46_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05495_ _00967_ _00983_ _01002_ _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_116_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07234_ cpu.timer_capture\[3\] _02674_ _02699_ _02687_ _02700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_73_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07165_ cpu.uart.divisor\[1\] _02641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_06116_ net62 _01089_ _01619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05503__S0 _00887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07096_ _02302_ _02342_ _02343_ _02582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_2_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06047_ _01550_ _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05357__I _00006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07998_ cpu.uart.receive_buff\[1\] _03291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06384__A1 net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05187__A2 cpu.spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09806_ _04793_ _04807_ _04808_ _04809_ _00746_ _00515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_09737_ _04754_ _00501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06949_ net20 _02075_ _02074_ _02444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09668_ _04691_ _04690_ _04696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09599_ cpu.orig_PC\[13\] _04033_ _04632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08619_ cpu.pwm_top\[0\] _03778_ _03780_ _03671_ _03781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_25_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_53_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05820__I _01325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10512_ _00450_ clknet_leaf_87_wb_clk_i cpu.ROM_addr_buff\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10443_ _00382_ clknet_leaf_26_wb_clk_i cpu.timer\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09389__B2 _04378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10374_ _00313_ clknet_leaf_86_wb_clk_i cpu.orig_PC\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06098__I _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05280_ cpu.regs\[12\]\[0\] cpu.regs\[13\]\[0\] cpu.regs\[14\]\[0\] cpu.regs\[15\]\[0\]
+ _00803_ _00573_ _00813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_3_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08970_ _04034_ _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_100_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_100_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07921_ _03230_ _03231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07852_ _03143_ _03150_ _03146_ _03172_ _03173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xinput1 io_in[0] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07392__I _02824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06803_ _02292_ _02299_ _02300_ _02301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07783_ _01403_ _03107_ _03110_ _00191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09522_ _04370_ _04553_ _04557_ _04558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06118__A1 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06734_ _02228_ _02229_ _02232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09453_ _04485_ _04489_ _04490_ _04491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06665_ _02160_ _02161_ _02163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05616_ _01066_ _01057_ _01122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09384_ _04353_ _04412_ _04424_ _04356_ _04425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_59_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08404_ _03613_ _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_19_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08335_ _02829_ _03557_ _03561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09112__I _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06596_ _00604_ _01956_ _02094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05547_ _01045_ _01048_ _01052_ _01053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_61_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08266_ _03506_ _00278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05478_ _00986_ _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08951__I _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08197_ _03453_ _03455_ _03381_ _00260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07217_ _02642_ _02679_ _02685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08043__A1 _02847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07148_ _01142_ _02626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_14_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07079_ _02541_ _02567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10090_ _00033_ clknet_leaf_101_wb_clk_i cpu.regs\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_58_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05580__A2 _01074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07857__A1 _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10426_ _00365_ clknet_leaf_27_wb_clk_i cpu.timer_div_counter\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_94_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10357_ _00296_ clknet_leaf_61_wb_clk_i cpu.needs_interrupt vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10288_ _00227_ clknet_leaf_66_wb_clk_i cpu.uart.dout\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06348__A1 _01326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06450_ _01949_ _01950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_118_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06520__A1 _01454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05401_ _00883_ _00913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_103_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06381_ cpu.uart.divisor\[6\] _01881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_44_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05332_ cpu.PORTB_DDR\[3\] net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_08120_ _03393_ _03389_ _03394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_71_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07076__A2 _02385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08051_ _02840_ cpu.uart.div_counter\[15\] _03335_ cpu.uart.divisor\[3\] _03336_
+ _03337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_05263_ _00784_ _00699_ _00797_ _00798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07002_ _02490_ _02493_ _02495_ _02496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_43_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05194_ _00698_ _00725_ _00730_ _00731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08953_ _04032_ _04042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07904_ _03203_ _03217_ _00205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08884_ _03985_ _00417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06339__A1 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07835_ _03155_ cpu.timer\[15\] cpu.timer\[14\] _03138_ _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_55_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07766_ _00851_ _03053_ _03096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07839__A1 cpu.timer_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07839__B2 cpu.timer_top\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09505_ _04455_ _04524_ _04540_ _04541_ _04542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06717_ _02213_ _02214_ _02215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_67_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09436_ cpu.orig_PC\[7\] _04043_ _04475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08500__A2 cpu.toggle_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07697_ _02067_ _02932_ _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_94_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06648_ _00834_ _01014_ _02146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_35_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09367_ _04407_ _04408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06579_ _02076_ _02077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08318_ _03510_ _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09298_ _04293_ _04332_ _04341_ _04342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08249_ _03495_ _03285_ _03496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07297__I _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10211_ _00150_ clknet_leaf_124_wb_clk_i cpu.regs\[7\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output77_I net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10142_ _00081_ clknet_leaf_101_wb_clk_i cpu.regs\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05250__A1 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10073_ _00016_ clknet_leaf_1_wb_clk_i cpu.regs\[9\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08856__I _03958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_qcpu_101 io_oeb[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_qcpu_112 io_oeb[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__06309__C _01108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09687__I _00790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09055__I0 cpu.regs\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10409_ _00348_ clknet_leaf_5_wb_clk_i cpu.toggle_ctr\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06569__A1 _01144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05950_ _00832_ _00929_ _01455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05881_ net40 _01385_ _01386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_108_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07620_ cpu.regs\[7\]\[2\] _02986_ _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_105_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06741__A1 _00919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07551_ _01165_ _02071_ _02948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_76_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08089__A4 _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06502_ _01999_ _02000_ _02001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07482_ _02902_ _02903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06286__I _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_66_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06219__C _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09221_ _00751_ _00767_ _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_44_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06433_ _01352_ _01800_ _01914_ _01350_ _01933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_17_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06364_ _01454_ _01836_ _01864_ _01865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09152_ _04196_ _01469_ _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08103_ _03226_ _03381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05315_ _00845_ net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_32_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09083_ _04137_ _04145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06295_ cpu.regs\[8\]\[6\] cpu.regs\[9\]\[6\] cpu.regs\[10\]\[6\] cpu.regs\[11\]\[6\]
+ _00888_ _00901_ _01796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_4_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08034_ cpu.uart.div_counter\[1\] _03320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_05246_ _00772_ _00777_ _00781_ _00782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_3_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05177_ _00709_ _00713_ _00714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_40_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09985_ _04680_ _04949_ _04915_ _04950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08936_ cpu.uart.divisor\[15\] _04013_ _04025_ _04020_ _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_4_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08867_ _03971_ _03973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07818_ cpu.timer_top\[13\] _03139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08798_ _03918_ _03920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_8_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_8_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07749_ _02374_ _03079_ _03080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_80_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08485__A1 _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09419_ _04293_ _04454_ _04458_ _04459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05299__A1 _00566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10044__A1 _04378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10044__B2 _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07460__A2 _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10125_ _00068_ clknet_leaf_11_wb_clk_i cpu.toggle_top\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07691__S _03026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10056_ cpu.regs\[15\]\[1\] _05014_ _05016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_100_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05526__A2 _01030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08228__A1 _02652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10035__A1 _01332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09976__A1 _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09028__I0 _00837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05100_ _00635_ _00639_ _00623_ _00640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06080_ _01580_ _01582_ _01584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_78_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_78_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05031_ _00573_ _00574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_111_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05214__A1 _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05065__I1 _00605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09770_ _04756_ _04779_ _04780_ _00508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_107_Right_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09880__I _04864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06982_ _02048_ _02475_ _02476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_111_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08721_ _03840_ _03856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05933_ _01034_ _00831_ _01438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08652_ cpu.timer_div_counter\[0\] cpu.timer_div_counter\[1\] cpu.timer_div_counter\[2\]
+ _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__05517__A2 _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06714__A1 _00930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07603_ _02945_ cpu.regs\[8\]\[6\] _02968_ _02978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05864_ _01306_ _01370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_37_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08583_ _03726_ _03754_ _03755_ _00346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05795_ _01300_ _01301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_66_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07534_ cpu.regs\[11\]\[1\] _02936_ _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07465_ cpu.regs\[14\]\[0\] _02893_ _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09204_ _03456_ _04248_ _04249_ _04250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06416_ _01836_ _01838_ _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07396_ cpu.uart.receive_div_counter\[13\] _02829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10026__A1 _00865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09967__B2 cpu.ROM_addr_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09967__A1 cpu.ROM_addr_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09135_ _04177_ _04183_ _04184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06347_ _01834_ _01846_ _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09066_ _04130_ cpu.ROM_addr_buff\[12\] _04126_ _04131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06278_ _01744_ _01779_ _01780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08017_ cpu.uart.dout\[6\] _03287_ _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05229_ _00753_ _00755_ _00757_ _00765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_13_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05205__A1 _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09968_ cpu.ROM_addr_buff\[9\] _02502_ _02477_ _04935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_99_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08919_ _04012_ _00425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09899_ _04018_ _04877_ _04880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06919__I _00621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10017__A1 cpu.orig_flags\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08630__A1 _02758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10108_ _00051_ clknet_leaf_22_wb_clk_i cpu.timer_capture\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10039_ _04986_ _02722_ _05002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_125_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_125_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_81_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05580_ _01071_ _01074_ _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08449__A1 _02393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07250_ _02713_ _00055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07181_ _02633_ _02654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06201_ _01167_ _01701_ _01703_ _00016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06132_ _01632_ _01634_ _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08621__A1 _03658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06063_ _01438_ _01439_ _01566_ _01567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09822_ _04822_ _00518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09753_ cpu.ROM_spi_dat_out\[2\] _04732_ _04767_ _04768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05294__S0 _00568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06965_ cpu.startup_cycle\[3\] cpu.startup_cycle\[2\] _02459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08704_ cpu.timer_capture\[0\] _03841_ _03842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09684_ _02045_ _02505_ _04710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08688__A1 _02658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05916_ cpu.toggle_top\[9\] _01259_ _01418_ _01420_ _01169_ _01421_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__07344__B _02567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06896_ _02393_ _02391_ _02394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08635_ _03792_ _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05847_ _01352_ _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_89_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08566_ cpu.toggle_ctr\[7\] _03743_ _03745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07360__A1 _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05778_ _01273_ _01278_ _01283_ _00920_ _01284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07517_ _02925_ _02918_ _02926_ _00109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08497_ _03678_ _03681_ _03682_ _03683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07448_ _02875_ _02879_ _00087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08860__A1 _02658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07663__A2 _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07379_ _02570_ _02385_ _02812_ _02816_ _02817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_09118_ _04169_ _04138_ _04170_ _03980_ _00466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_72_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10390_ _00329_ clknet_leaf_14_wb_clk_i cpu.toggle_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_20_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09049_ _04118_ cpu.ROM_addr_buff\[7\] _04115_ _04119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09168__A2 _02185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08679__A1 _02644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06154__A2 _00997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07351__A1 _02168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07103__A1 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08851__A1 cpu.spi.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10588_ _00526_ clknet_leaf_67_wb_clk_i net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07406__A2 cpu.uart.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09159__A2 _00988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05463__I _00972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06750_ _02246_ _02247_ _02248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_05701_ _01200_ _01207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06681_ _00800_ _01954_ _02179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08420_ cpu.orig_PC\[4\] _03607_ _03626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05632_ cpu.br_rel_dest\[3\] _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08351_ net17 _03574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_05563_ _00679_ _01069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_117_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08282_ cpu.uart.receive_div_counter\[2\] cpu.uart.receive_div_counter\[1\] cpu.uart.receive_div_counter\[0\]
+ _03519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__08842__A1 cpu.timer_capture\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07302_ _02753_ _00067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05494_ _00960_ _00980_ _01002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07233_ _02696_ _02677_ _02691_ _02698_ _02699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_61_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_93_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_93_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_46_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05656__A1 _01161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09398__A2 _00754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07164_ _02640_ _00042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_22_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_22_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_42_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06115_ net42 _01510_ _01614_ _01617_ _01089_ _01618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_42_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07095_ _02581_ _00032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_67_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05503__S1 _00900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06081__A1 _01471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06046_ _00845_ _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07997_ _03283_ _03288_ _03290_ _02628_ _00225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09805_ _03758_ _03760_ cpu.pwm_counter\[3\] _03763_ _04809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_09736_ _03120_ _04753_ _04754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06948_ _02064_ _02442_ _02443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09667_ cpu.mem_cycle\[4\] _04691_ _04690_ _04695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_69_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05373__I _00869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08618_ _02636_ _03779_ _03780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06879_ cpu.PC\[8\] _02377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07884__A2 _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09598_ _04623_ _04625_ _04630_ _00777_ _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09086__A1 _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08549_ cpu.toggle_ctr\[2\] _03730_ _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_TAPCELL_ROW_25_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10511_ _00449_ clknet_leaf_83_wb_clk_i cpu.ROM_addr_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05647__A1 _01029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10442_ _00381_ clknet_leaf_26_wb_clk_i cpu.timer\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08061__A2 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10373_ _00312_ clknet_leaf_89_wb_clk_i cpu.orig_PC\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09010__A1 _00865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09183__C _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07572__A1 _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05886__A1 _01090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05430__S0 _00878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08824__A1 _00989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05886__C _01390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07920_ cpu.spi.counter\[0\] _03200_ _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05810__A1 _01131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07851_ cpu.timer_top\[10\] _03170_ _03171_ cpu.timer_top\[9\] _03172_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput2 io_in[10] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07782_ cpu.spi.data_in_buff\[1\] _03108_ _03109_ _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06802_ _02297_ _02298_ _02300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09521_ _00952_ _04444_ _04556_ _04448_ _04557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06733_ _02230_ _02231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_108_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08718__B _03853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07315__A1 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07866__A2 cpu.spi.divisor\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09452_ _03057_ _04489_ _04490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06664_ _02160_ _02161_ _02162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09383_ cpu.orig_PC\[5\] _04354_ _04424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05615_ _01029_ _00759_ _01120_ _01121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_08403_ _02781_ _03613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06595_ _02091_ _02092_ _02093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08334_ _03553_ _03560_ _00292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05546_ _00649_ _01051_ _01052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_22_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07618__A2 _02985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08265_ cpu.uart.receive_buff\[7\] _03503_ _03497_ cpu.uart.receive_buff\[6\] _03506_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_61_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05477_ _00985_ _00986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08196_ _03454_ _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07216_ _02683_ _02684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07147_ _02610_ _02622_ _02625_ _02618_ _00040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_15_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05101__I0 cpu.regs\[12\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07078_ _02559_ _02565_ _02566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06029_ cpu.timer_top\[2\] _01382_ _01533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06357__A2 _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09719_ cpu.ROM_spi_dat_out\[0\] _04737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_97_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_6_0_wb_clk_i clknet_0_wb_clk_i clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_2_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09303__I _04292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_17_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10425_ _00364_ clknet_leaf_15_wb_clk_i cpu.pwm_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07093__I0 _01950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10356_ _00295_ clknet_leaf_34_wb_clk_i cpu.uart.receive_div_counter\[15\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_94_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10287_ _00226_ clknet_leaf_66_wb_clk_i cpu.uart.dout\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09534__A2 _04407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_29_Left_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_1_Left_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_75_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_56_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05400_ cpu.regs\[12\]\[1\] cpu.regs\[13\]\[1\] cpu.regs\[14\]\[1\] cpu.regs\[15\]\[1\]
+ _00899_ _00902_ _00912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XPHY_EDGE_ROW_38_Left_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_103_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06380_ cpu.spi.dout\[6\] _01880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09470__A1 _01020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05331_ _00860_ net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08050_ cpu.uart.divisor\[11\] cpu.uart.div_counter\[11\] _03336_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_98_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05262_ _00698_ _00704_ _00796_ _00797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__06284__A1 net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07001_ cpu.spi_clkdiv _02494_ _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05193_ _00729_ _00730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09816__C _04765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_47_Left_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08952_ _04040_ _04041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07903_ _03196_ _03216_ _03217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08883_ cpu.timer_div\[4\] _03976_ _03984_ _03956_ _03985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07834_ cpu.timer_top\[15\] _03155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07536__A1 cpu.regs\[11\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05398__I0 cpu.regs\[8\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07765_ _01699_ _03094_ _02401_ _03095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_69_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08448__B _03646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09504_ _04338_ _04541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06716_ _00800_ _01015_ _02214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07696_ _02997_ _03029_ _03037_ _00177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_56_Left_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09435_ _04312_ _04473_ _04474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06647_ cpu.regs\[1\]\[3\] _00985_ _02145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09366_ _03622_ _04348_ _04407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06578_ _01549_ _01030_ _01151_ _02076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_35_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08317_ _03522_ _03546_ _00289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_117_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09297_ _04333_ _04297_ _04337_ _04339_ _04340_ _04341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_34_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05529_ _01034_ _01035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08248_ _02867_ _03495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_62_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08179_ cpu.uart.counter\[0\] _03441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06027__A1 cpu.timer_capture\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_65_Left_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10210_ _00149_ clknet_4_0_0_wb_clk_i cpu.regs\[7\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06578__A2 _01030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10141_ _00080_ clknet_leaf_101_wb_clk_i cpu.regs\[1\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05826__I _01331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10072_ _00015_ clknet_leaf_1_wb_clk_i cpu.regs\[9\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_74_Left_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_qcpu_113 io_oeb[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xwrapped_qcpu_102 io_oeb[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_38_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09452__A1 _03057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09055__I1 _03637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09204__A1 _03456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10408_ _00347_ clknet_leaf_5_wb_clk_i cpu.toggle_ctr\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10339_ _00278_ clknet_leaf_43_wb_clk_i cpu.uart.receive_buff\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07766__A1 _00851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05880_ _01112_ _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_108_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07550_ _02930_ _02936_ _02947_ _00121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06567__I _01130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06501_ _01914_ _01917_ _01912_ _02000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09220_ _04264_ _04265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07481_ _01137_ _02889_ _02902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_29_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06432_ net96 _01931_ _01932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_60_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06363_ _01706_ _01351_ _01835_ _01339_ _00720_ _01864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_17_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09151_ _01476_ _01580_ _01670_ _04198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_32_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08102_ _03320_ _03365_ _03379_ _03380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09082_ _03360_ _04139_ _04144_ _00456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_83_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05314_ _00566_ _00839_ _00844_ _00845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_08033_ cpu.uart.divisor\[10\] _03318_ cpu.uart.div_counter\[8\] _02827_ _03319_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06294_ cpu.regs\[12\]\[6\] cpu.regs\[13\]\[6\] cpu.regs\[14\]\[6\] cpu.regs\[15\]\[6\]
+ _00898_ _00901_ _01795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_32_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05245_ _00778_ _00779_ _00780_ _00781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_24_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05176_ _00710_ _00712_ _00713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_4_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09984_ _02478_ _04944_ _04946_ _04948_ _04949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__05232__A2 _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08935_ _02775_ _04015_ _04025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input21_I io_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08866_ _03971_ _03972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07817_ cpu.timer_top\[14\] _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08797_ _03918_ _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08178__B _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07748_ _02389_ _03078_ _03079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_94_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07679_ _03027_ _03028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_109_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09418_ _04455_ _04433_ _04457_ _04339_ _04340_ _04458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_75_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09434__A1 _02626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09349_ _04299_ _04383_ _04390_ _04310_ _04391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_90_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10044__A2 _04985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09037__I1 cpu.ROM_addr_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10124_ _00067_ clknet_leaf_11_wb_clk_i cpu.toggle_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__06420__A1 _01437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08867__I _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10055_ _01373_ _05013_ _05015_ _00558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08173__A1 _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_82_Left_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_91_Left_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06239__B2 _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06239__A1 _01004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09028__I1 _02810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05030_ _00001_ _00573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07739__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06981_ _02056_ _02058_ _02475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__05065__I2 _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_47_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_47_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08720_ cpu.timer\[3\] _03854_ _03855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05932_ _01315_ _01437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08164__A1 _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08651_ _03802_ _03803_ _00366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05863_ net26 _01368_ _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07602_ _02977_ _00143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_37_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05794_ _01039_ _01041_ _01300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08582_ cpu.toggle_ctr\[13\] _03753_ _03755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_66_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07533_ _02914_ _02935_ _02937_ _00114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06478__A1 _01976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07464_ _02890_ _02893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09203_ _00764_ _04249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06415_ _01913_ _01914_ _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_29_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07395_ _02825_ cpu.uart.receive_div_counter\[12\] _02826_ _02827_ _02828_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09134_ _00728_ _04182_ _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06346_ _01834_ _01846_ _01847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10026__A2 _04985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09065_ cpu.regs\[3\]\[4\] _02393_ _04101_ _04130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06277_ _01689_ _01778_ _01779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08016_ cpu.uart.receive_buff\[6\] _03304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05228_ _00714_ _00658_ _00764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05159_ _00696_ _00697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05205__A2 _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05376__I _00887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09967_ cpu.ROM_addr_buff\[1\] _04927_ _02501_ cpu.ROM_addr_buff\[5\] cpu.ROM_addr_buff\[13\]
+ _02486_ _04934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08918_ cpu.uart.divisor\[11\] _04001_ _04011_ _04006_ _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09898_ _04879_ _00537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_99_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08849_ cpu.spi.divisor\[1\] _03960_ _03962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08458__A2 _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06469__A1 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10017__A2 _04032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07969__A1 _00788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08394__A1 _00794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10107_ _00050_ clknet_leaf_30_wb_clk_i cpu.timer_capture\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10038_ _04040_ _04992_ _04998_ _05000_ _05001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_98_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05380__B2 _00891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06200_ cpu.regs\[9\]\[3\] _01702_ _01703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07180_ _02652_ _02653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_54_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06131_ cpu.timer_div\[3\] _01406_ _01633_ _01634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06580__I _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06632__A1 _00638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06062_ _01034_ _00832_ _01566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_113_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05196__I _00671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09821_ net60 _04814_ _04820_ _04821_ _04822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05199__A1 _00671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09752_ _04741_ _04745_ _04715_ _04767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06964_ _02457_ _02450_ _02458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08703_ _03840_ _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05924__I _01354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09683_ _02040_ _04708_ _02506_ _02499_ _04709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_05915_ _01419_ _01173_ _01259_ _01420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06895_ _02375_ _02393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08634_ cpu.pwm_top\[4\] _03787_ _03791_ _03783_ _03792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05846_ _01351_ _01352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08565_ _03697_ _03698_ _03739_ _03744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_05777_ _01282_ _01283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07516_ cpu.regs\[12\]\[3\] _02917_ _02926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08496_ cpu.toggle_ctr\[11\] _01646_ _01538_ _03679_ _03682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_9_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07447_ _02873_ _02878_ cpu.uart.receive_counter\[1\] _02879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_107_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05674__A2 _01082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07378_ _02570_ _02815_ _02816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09117_ cpu.ROM_addr_buff\[10\] _04137_ _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06329_ _01281_ _01801_ _01829_ _01542_ _01830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_32_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09048_ cpu.regs\[2\]\[7\] _02588_ _04117_ _04118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_20_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06387__B1 _01884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output52_I net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06862__A1 _00605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05504__I3 cpu.regs\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10587_ _00525_ clknet_leaf_67_wb_clk_i net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09159__A3 _01018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_10_Left_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09216__I _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_2_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05700_ _01205_ _01206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06680_ _00835_ _00986_ _01016_ _00821_ _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05631_ _01130_ _01136_ _01137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__08276__B _02871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08350_ _00745_ _03573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_63_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05562_ _01061_ _01068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07301_ cpu.toggle_top\[9\] _02749_ _02752_ _02712_ _02753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_19_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06575__I _02072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08281_ _02833_ _02834_ _03518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05493_ _01001_ net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07232_ _00998_ _02697_ _02698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05656__A2 _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07163_ _02629_ _02634_ _02638_ _02639_ _02640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_42_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06114_ net82 _01615_ _01616_ _01617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_42_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07094_ _02416_ _02580_ _02544_ _02581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_62_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_62_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_41_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06045_ _01548_ _01549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_74_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07030__A1 _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09804_ cpu.pwm_counter\[5\] _03769_ cpu.pwm_counter\[7\] cpu.pwm_counter\[6\] _04808_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_07996_ cpu.uart.dout\[0\] _03289_ _03290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09858__A1 net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09735_ _04737_ _04751_ _04752_ _04753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08030__I _02629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06947_ _02429_ _02435_ _02441_ _02442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09666_ _04694_ _00490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_97_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08617_ _03777_ _03779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06878_ cpu.PC\[9\] _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09597_ _04621_ _04629_ _04440_ _04630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05829_ _00863_ _00867_ _01150_ _01335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_65_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08548_ _03725_ _03732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08479_ cpu.toggle_top\[4\] _03666_ _03668_ _03660_ _03669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07097__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10510_ _00448_ clknet_leaf_82_wb_clk_i cpu.ROM_addr_buff\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08833__A2 _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05647__A2 _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10441_ _00380_ clknet_leaf_19_wb_clk_i cpu.timer_top\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07249__C _02712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10372_ _00311_ clknet_leaf_86_wb_clk_i cpu.orig_PC\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09849__A1 _04815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07572__A2 _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09480__B _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05430__S1 _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05810__A2 _00816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07850_ cpu.timer\[9\] _03171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07781_ _00789_ _03109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_85_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08760__A1 cpu.timer_capture\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06801_ _02297_ _02298_ _02299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput3 io_in[11] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09520_ _04554_ _04555_ _04319_ _04556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06732_ _02228_ _02229_ _02230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_108_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09451_ _04408_ _04489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06663_ _02131_ _02132_ _02161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08402_ _01607_ _03589_ _03612_ _03591_ _00308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_59_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05614_ cpu.br_rel_dest\[7\] _00754_ _01120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09382_ _00763_ _04419_ _04422_ _04423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_47_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06594_ _00636_ _00986_ _02092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08333_ cpu.uart.receive_div_counter\[12\] _03547_ _03557_ _03559_ _03560_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05545_ _01050_ _01051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_22_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08264_ _03505_ _00277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_50_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05476_ _00984_ _00985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_116_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08028__B1 _01612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08195_ _03439_ _03450_ _03454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07215_ cpu.timer\[1\] _02683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07146_ _01877_ _02620_ _02625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07077_ _02560_ _02564_ _02374_ _02565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09240__A2 _04252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06028_ _01499_ _01234_ _01530_ _01531_ _01382_ _01532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09718_ _03227_ _04736_ _00500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07979_ _03269_ _03277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_58_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09649_ _04680_ _04681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_2_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10424_ _00363_ clknet_leaf_19_wb_clk_i cpu.pwm_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10355_ _00294_ clknet_leaf_34_wb_clk_i cpu.uart.receive_div_counter\[14\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_94_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10286_ _00225_ clknet_leaf_66_wb_clk_i cpu.uart.dout\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_2_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05330_ _00859_ _00860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06808__A1 _00822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05261_ _00794_ cpu.needs_interrupt _00795_ _00796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07481__A1 _01137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07000_ cpu.ROM_spi_cycle\[0\] _02447_ _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_72_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05192_ _00728_ _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_102_Left_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08951_ _01449_ _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07902_ _03206_ _03215_ _03216_ _00204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08882_ _02762_ _03983_ _03984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07833_ _03143_ _03151_ _03153_ _03154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06339__A3 _01758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_81_Right_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_55_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09404__I _04313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07764_ net20 _03054_ _03093_ _03094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09503_ _00823_ _04515_ _04540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06715_ _00820_ _02083_ _02213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07695_ cpu.regs\[4\]\[7\] _03027_ _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_69_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09434_ _02626_ _04444_ _04472_ _04448_ _04473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06646_ _02143_ _02144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_111_Left_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_35_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09365_ _02563_ _04344_ _04406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06577_ _02062_ _02075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08316_ _03543_ _03511_ _03545_ _03541_ _03546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09296_ _04194_ _04340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_47_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06763__I _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05528_ cpu.br_rel_dest\[1\] _01034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08247_ _03493_ _03494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_104_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_90_Right_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05459_ cpu.regs\[8\]\[3\] cpu.regs\[9\]\[3\] cpu.regs\[10\]\[3\] cpu.regs\[11\]\[3\]
+ _00962_ _00963_ _00969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05322__I1 _00850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08178_ cpu.uart.counter\[0\] _03439_ _03340_ _03440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_30_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07129_ _02611_ _02601_ _02612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_30_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10140_ _00079_ clknet_leaf_103_wb_clk_i cpu.regs\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10071_ _00014_ clknet_leaf_2_wb_clk_i cpu.regs\[9\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08724__A1 cpu.timer_capture\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09742__C _04684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_qcpu_114 io_oeb[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xwrapped_qcpu_103 io_oeb[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_97_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmax_cap98 _02279_ net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10536__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05289__I _00820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10407_ _00346_ clknet_leaf_4_wb_clk_i cpu.toggle_ctr\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10338_ _00277_ clknet_leaf_44_wb_clk_i cpu.uart.receive_buff\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_119_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_119_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10269_ _00208_ clknet_leaf_64_wb_clk_i cpu.spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_17_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06500_ _01993_ _01998_ _01999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07480_ _02033_ _02893_ _02901_ _00097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06431_ net95 _01762_ _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_60_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06362_ _01841_ _01762_ _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09150_ _04196_ _01359_ _00714_ _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08101_ _03378_ _03379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09081_ cpu.last_addr\[0\] _04143_ _04144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06293_ _01792_ _01793_ _00885_ _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06257__A2 _01758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05313_ _00566_ _00841_ _00843_ _00844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08032_ cpu.uart.div_counter\[10\] _03318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09894__I _04864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05244_ cpu.instr_buff\[14\] _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_4_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05175_ _00711_ cpu.instr_buff\[14\] _00712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09983_ _00670_ _04947_ _04701_ _04948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05768__A1 _00706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08934_ _04024_ _00428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_4_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08865_ _01073_ _01098_ _01235_ _02632_ _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__08182__A2 _03368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08796_ _01074_ _01235_ _02632_ _03918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_07816_ _03136_ _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input14_I io_in[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05662__I _01121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07747_ _03076_ _02388_ _03077_ _03078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05940__A1 _01437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07678_ _03026_ _03027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_80_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09417_ _02416_ _04375_ _04456_ _04457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06629_ _02110_ _02111_ _02127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09348_ _04387_ _04388_ _04389_ _04390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_62_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09279_ _04312_ _04322_ _04323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08945__A1 _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10123_ _00066_ clknet_leaf_11_wb_clk_i cpu.toggle_top\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10054_ cpu.regs\[15\]\[0\] _05014_ _05015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_7_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05782__I1 cpu.regs\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06487__A2 _01957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09189__A1 _01311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06980_ _02468_ _02059_ _02473_ _02474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__05065__I3 cpu.regs\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input6_I io_in[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05931_ _01434_ _01435_ _01305_ _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08650_ _03127_ cpu.timer_div_counter\[1\] _03803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05862_ _01157_ _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07601_ _02943_ cpu.regs\[8\]\[5\] _02968_ _02977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_37_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_87_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_87_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05922__A1 _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08581_ cpu.toggle_ctr\[13\] _03753_ _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05793_ _01269_ _01299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_66_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_16_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_16_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07532_ cpu.regs\[11\]\[0\] _02936_ _02937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_45_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07463_ _02891_ _02892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09202_ _00725_ _04247_ _04248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_57_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06414_ _00631_ _01800_ _01914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07394_ cpu.uart.divisor\[8\] _02827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_09133_ _04178_ _04180_ _04181_ _04182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06345_ _01770_ _01839_ _01845_ _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09064_ _04129_ _00453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06276_ _01752_ _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08015_ _03302_ _03298_ _03303_ _03296_ _00230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_71_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05227_ _00762_ _00763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05158_ _00695_ _00696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08927__A1 _04018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09129__I _04032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09966_ net72 _04933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07872__I cpu.spi.divisor\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08968__I _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05089_ _00599_ _00624_ _00629_ _00630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_09897_ cpu.PORTB_DDR\[4\] _04876_ _04878_ _04870_ _04879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08917_ _04010_ _04002_ _04011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08848_ _02726_ _03959_ _03961_ _00405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09352__A1 _01704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08779_ cpu.timer\[13\] _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_94_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06469__A2 _01390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07418__B2 _02847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07969__A2 _03223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08918__A1 cpu.uart.divisor\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09591__A1 _00772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10106_ _00049_ clknet_leaf_31_wb_clk_i cpu.uart.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10037_ _01466_ _04993_ _04999_ _01462_ _04196_ _05000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__05904__A1 cpu.timer_capture\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07657__A1 _01137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07022__I _02513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06130_ _01180_ _01633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06061_ _01563_ _01564_ _01565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_113_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08909__A1 _03658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09820_ _04683_ _04821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09582__A1 _00591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09751_ _04766_ _00503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06963_ cpu.startup_cycle\[6\] _02457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08702_ _01059_ _02747_ _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__09334__A1 _02108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05914_ cpu.toggle_top\[1\] _01419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09682_ _02449_ _02042_ _04705_ _04707_ _04708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_06894_ _02375_ _02391_ _02392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__06148__A1 _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08633_ _02762_ _03788_ _03791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05845_ _00657_ _01338_ _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_89_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08564_ _03732_ _03742_ _03743_ _00339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05776_ _01281_ _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09637__A2 cpu.ROM_addr_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07515_ _01700_ _02925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08495_ _03679_ _01538_ _03677_ _03680_ _03681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07446_ _02870_ _02877_ _02878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06320__A1 cpu.timer_capture\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07377_ _02405_ _02335_ _02814_ _02583_ _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_29_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07867__I cpu.spi.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09116_ cpu.last_addr\[10\] _04169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_79_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06328_ _01275_ _01828_ _01829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09047_ _04101_ _04117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_20_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06259_ _01139_ _01654_ _01761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__05387__I _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06387__A1 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08698__I _03835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09949_ _04703_ _02041_ _02454_ _02461_ _04918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__06139__A1 _01609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09750__C _04765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_36_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06311__A1 _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06862__A2 _01996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10586_ _00524_ clknet_leaf_68_wb_clk_i net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_23_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07811__A1 cpu.timer_div\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07811__B2 cpu.timer_div\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06378__A1 _01877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_75_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07878__B2 cpu.spi.divisor\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05889__B1 _01391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05630_ _01135_ _01136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_59_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05561_ _01066_ _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_63_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07300_ _02732_ _02750_ _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08280_ _02849_ _03517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05492_ _00990_ _01000_ _01001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07231_ _02676_ _02697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07162_ _02521_ _02639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06113_ _01509_ _01616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_41_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07802__A1 cpu.timer_div\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07093_ _01950_ _02579_ _02567_ _02580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06044_ _01356_ _01548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_2_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09803_ _04800_ _04803_ _04806_ _04807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06369__A1 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07995_ _03286_ _03289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09307__A1 _03623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09734_ _04743_ _04746_ _04749_ _02497_ _04752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
Xclkbuf_leaf_31_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_31_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06946_ _02415_ _02432_ _02433_ _02441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09665_ _04691_ _04643_ _04693_ _04684_ _04694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07869__B2 cpu.spi.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06877_ cpu.PC\[12\] _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08616_ _03777_ _03778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08530__A2 _01261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05828_ _01332_ _01333_ _01334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09596_ cpu.PC\[13\] _00925_ _04628_ _04629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08547_ _03729_ _03730_ _03731_ _00334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05759_ _01142_ _01154_ _01265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_25_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08478_ _02762_ _03667_ _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07429_ cpu.uart.receive_div_counter\[10\] _02862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05647__A3 _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10440_ _00379_ clknet_leaf_18_wb_clk_i cpu.timer_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10371_ _00310_ clknet_leaf_89_wb_clk_i cpu.orig_PC\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06006__I _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09546__A1 cpu.PC\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09761__B _03761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07572__A3 _01390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06532__A1 _01370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06532__B2 _02030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10569_ _00507_ clknet_leaf_75_wb_clk_i cpu.ROM_spi_dat_out\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07780_ _03105_ _03108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06800_ _02269_ _02270_ _02278_ _02298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xinput4 io_in[12] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06731_ _02193_ _02195_ _02229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_108_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09450_ _04266_ _04488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08401_ cpu.orig_flags\[3\] _03611_ _03612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06662_ _02144_ _02158_ _02159_ _02160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05613_ _01114_ _01118_ _01119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09381_ _00752_ _04314_ _04421_ _04321_ _04422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06593_ _00620_ _01016_ _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08332_ _02830_ _03558_ _03513_ _03559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_86_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05544_ cpu.IO_addr_buff\[3\] _01049_ _01050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_47_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08263_ cpu.uart.receive_buff\[6\] _03503_ _03497_ cpu.uart.receive_buff\[5\] _03505_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_50_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07214_ _02682_ _00050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_62_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05475_ _00980_ _00983_ _00883_ _00984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08194_ cpu.uart.counter\[3\] _03452_ _03453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07145_ _02607_ _02622_ _02624_ _02618_ _00039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_14_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07076_ _02561_ _02385_ _02563_ _02564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06027_ cpu.timer_capture\[2\] _01236_ _01234_ _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09528__A1 _00837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09137__I _04180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07978_ _03276_ _00220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09717_ cpu.spi_clkdiv _02497_ _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07880__I _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06929_ net12 _02404_ _02064_ _02406_ _02425_ _02426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_97_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08197__B _03381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09648_ _04656_ _04658_ _04659_ _04679_ _04680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_85_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06496__I _01994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09579_ _04347_ _04599_ _04612_ _04373_ _04613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08267__A1 _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07120__I _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10423_ _00362_ clknet_leaf_15_wb_clk_i cpu.pwm_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10354_ _00293_ clknet_leaf_36_wb_clk_i cpu.uart.receive_div_counter\[13\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09519__A1 _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10285_ _00224_ clknet_leaf_48_wb_clk_i cpu.spi.data_in_buff\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08886__I _02771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09491__B _04440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06505__A1 _01992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06355__B _01335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06808__A2 _00955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05260_ _00701_ net18 _00795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09058__I0 cpu.regs\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07481__A2 _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05191_ _00727_ _00728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08950_ _04029_ _04039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07901_ cpu.spi.div_counter\[5\] _03214_ _03216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08881_ _03971_ _03983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09930__A1 _02657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07832_ cpu.timer_top\[12\] _03141_ _03152_ _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06744__A1 _00918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05398__I2 cpu.regs\[10\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09502_ _04514_ _04524_ _04539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07763_ _03088_ _03092_ _03051_ _03093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_55_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07544__I0 _02943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07694_ _03036_ _00176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06714_ _00930_ _02207_ _02211_ _02212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__07205__I _02673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09433_ _04364_ _04462_ _04471_ _04446_ _04472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06645_ _02140_ _02142_ _02143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08249__A1 _03495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09364_ _04382_ _04405_ _04381_ _00477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08315_ _03543_ _03544_ _03545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06576_ _02072_ _02074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_35_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09295_ _04338_ _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05527_ _01032_ _01033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08246_ _02865_ _03284_ _03493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_105_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05458_ cpu.regs\[12\]\[3\] cpu.regs\[13\]\[3\] cpu.regs\[14\]\[3\] cpu.regs\[15\]\[3\]
+ _00962_ _00963_ _00968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08177_ _00726_ _03366_ _03367_ _00766_ _03439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_50_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05322__I2 _00851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05389_ _00900_ _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07128_ _01159_ _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_112_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05395__I _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07059_ _02381_ _02548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_7_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10070_ _00013_ clknet_leaf_2_wb_clk_i cpu.regs\[9\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_102_Right_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08639__C _03795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08488__A1 _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_qcpu_115 io_oeb[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xwrapped_qcpu_104 io_oeb[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_66_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10406_ _00345_ clknet_leaf_4_wb_clk_i cpu.toggle_ctr\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08412__A1 _02810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05226__A1 _00751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10337_ _00276_ clknet_leaf_45_wb_clk_i cpu.uart.receive_buff\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10268_ _00207_ clknet_leaf_63_wb_clk_i net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09912__A1 _04815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10199_ _00138_ clknet_leaf_0_wb_clk_i cpu.regs\[8\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08479__A1 cpu.toggle_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06430_ _00632_ _01929_ _01930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_57_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10038__A1 _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06361_ _01152_ _01839_ _01859_ _01861_ _01862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_32_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08100_ _03377_ _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09080_ _04142_ _04143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_83_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06292_ cpu.regs\[0\]\[6\] cpu.regs\[1\]\[6\] cpu.regs\[2\]\[6\] cpu.regs\[3\]\[6\]
+ _00888_ _00889_ _01793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_05312_ _00580_ _00842_ _00843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08031_ _02857_ cpu.uart.div_counter\[10\] cpu.uart.div_counter\[0\] _03316_ _03317_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_05243_ _00687_ _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_25_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05174_ cpu.instr_buff\[15\] _00711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05217__A1 _00655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09982_ _02485_ _02598_ _04947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08933_ _02847_ _04013_ _04023_ _04020_ _04024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_110_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09903__A1 _04022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08864_ _02670_ _03965_ _03970_ _00412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09415__I _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07765__I0 _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07815_ _03123_ _03124_ _03132_ _03135_ _03136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_08795_ _03917_ _00396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07746_ cpu.PC\[10\] _03077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_67_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09416_ _04335_ _04433_ _04456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07142__A1 _01704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07677_ _02915_ _02982_ _03026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_39_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08890__A1 _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10029__A1 _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06628_ _02122_ _02125_ _02126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06559_ _02056_ _02057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_81_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09347_ _04387_ _04388_ _04306_ _04389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09278_ _02611_ _04314_ _04320_ _04321_ _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_35_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08229_ cpu.uart.data_buff\[5\] _03475_ _03481_ _03462_ _03482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08945__A2 _01704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06405__B1 _01266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output75_I net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10122_ _00065_ clknet_leaf_19_wb_clk_i cpu.timer_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10053_ _05011_ _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05067__S0 _00572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06184__A2 _00956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07381__A1 _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05782__I2 cpu.regs\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08385__B _03570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08633__A1 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_111_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05930_ cpu.Z _01297_ _01435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05861_ _01329_ _01334_ _01364_ net90 _01366_ _01367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_08580_ _03726_ _03752_ _03753_ _00345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07600_ _02976_ _00142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_37_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05792_ _01284_ _01285_ _01296_ _01297_ _01298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_07531_ _02933_ _02936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08295__B _03529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08872__A1 _03658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07462_ _02890_ _02891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07393_ cpu.uart.receive_div_counter\[8\] _02826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09201_ _04243_ _04246_ _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_45_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06413_ _01912_ _01913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_56_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_56_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_60_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09132_ _00753_ _00758_ _04181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06344_ _01770_ _01844_ _01845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09063_ _04128_ cpu.ROM_addr_buff\[11\] _04126_ _04129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06275_ _01774_ _01776_ _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08014_ cpu.uart.dout\[5\] _03294_ _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05226_ _00751_ _00761_ _00762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05157_ _00694_ _00670_ _00695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_77_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09965_ _04932_ _00551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05205__A4 _00728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05088_ _00567_ _00626_ _00628_ _00629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09896_ _04014_ _04877_ _04878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08916_ _02647_ _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_99_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08847_ cpu.spi.divisor\[0\] _03960_ _03961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_26_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08778_ _03902_ _03903_ _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07115__A1 _00696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07729_ _00802_ _03053_ _03062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08863__A1 cpu.spi.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08615__A1 _01087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05429__A1 _00870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05848__I _01345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06929__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05583__I _01088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_65_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10105_ _00048_ clknet_leaf_32_wb_clk_i cpu.uart.divisor\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10036_ _04986_ _02016_ _04999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07106__A1 _01370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07106__B2 _02030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08854__A1 _02648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07303__I _00946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09658__C _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06060_ _01159_ net92 _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_113_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05840__A1 _00816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07593__A1 cpu.regs\[8\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_103_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_103_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09750_ cpu.ROM_spi_dat_out\[2\] _04760_ _04764_ _04765_ _04766_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06962_ cpu.startup_cycle\[4\] _02456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09681_ _04706_ _04707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08701_ cpu.timer\[0\] _03834_ _03836_ _03838_ _03839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05493__I _01001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05913_ _01415_ _01416_ _01417_ _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08632_ _03790_ _00360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06893_ _02390_ _02391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07345__A1 _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05844_ _01349_ _01338_ _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__09098__A1 cpu.ROM_addr_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08563_ _03699_ _03739_ _03743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05775_ _01279_ _01094_ _01280_ _01038_ _01281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_76_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08494_ cpu.toggle_ctr\[9\] _03680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07514_ _02923_ _02918_ _02924_ _00108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07445_ _02823_ _02876_ _02877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_71_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07376_ _02331_ _02813_ _02334_ _02814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09115_ _04166_ _04167_ _04168_ _00465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_72_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06327_ _01121_ _01826_ _01827_ _01266_ _01004_ _01828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_45_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09046_ _04116_ _00448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06258_ _01680_ _01683_ _01760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05209_ _00745_ _00746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05831__A1 _01299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07883__I _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06189_ _01680_ _01691_ _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09948_ _02475_ _04916_ _04917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07584__A1 _01833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09879_ _04864_ _04865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08533__B1 cpu.toggle_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09089__A1 _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output38_I net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08836__A1 cpu.timer_capture\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06448__B _01379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07123__I _02524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10585_ _00523_ clknet_leaf_68_wb_clk_i net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_36_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05822__A1 _01326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_1_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_1_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10136__D _00075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06202__I _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07327__A1 cpu.toggle_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10019_ _01354_ _01280_ _04981_ _04982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_98_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05560_ _01065_ _00648_ _01066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_25_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05491_ _00949_ _00974_ _00999_ _01000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07230_ cpu.timer\[3\] _02696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_109_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07161_ _02636_ _02637_ _02638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08055__A2 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06112_ _01210_ _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07092_ _02578_ _02579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06043_ _01305_ _01546_ _01547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_74_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09802_ cpu.pwm_top\[1\] _04797_ _04804_ cpu.pwm_top\[2\] _04805_ _04806_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_07994_ _03287_ _03288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09733_ _04750_ _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06112__I _01210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06945_ cpu.regs\[2\]\[7\] _02070_ _02440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09664_ _04642_ _04681_ _04692_ _04693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06876_ _01366_ _01156_ _01349_ _02374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_96_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08615_ _01087_ _02747_ _03777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09595_ _04626_ _04601_ _04627_ _04628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05827_ _01311_ _01319_ _01333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_71_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_71_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_85_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08818__A1 _00998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08546_ _03652_ cpu.toggle_ctr\[0\] cpu.toggle_ctr\[1\] _03731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05758_ _01261_ _01263_ _01264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05689_ _01194_ _01195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_92_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08477_ _03653_ _03667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07428_ _02847_ _02846_ _02860_ cpu.uart.divisor\[5\] _02861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07359_ _02546_ _02794_ _02798_ _02799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09243__B2 _04256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10370_ _00309_ clknet_leaf_89_wb_clk_i cpu.orig_PC\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09029_ _03997_ _04104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07557__A1 cpu.regs\[10\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07309__A1 _02758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06532__A2 _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_99_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_116_Right_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10568_ _00506_ clknet_leaf_75_wb_clk_i cpu.ROM_spi_dat_out\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10499_ _00437_ clknet_leaf_90_wb_clk_i cpu.IO_addr_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06220__A1 cpu.spi.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput5 io_in[13] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_79_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06730_ _02224_ _02226_ _02227_ _02228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_108_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06661_ _02156_ _02157_ _02159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08400_ _03586_ _03611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05612_ _01052_ _01117_ _01118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09380_ _04316_ _04411_ _04420_ _04319_ _04421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06592_ _02088_ _02089_ _02086_ _02090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_19_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08331_ _03554_ _03548_ _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05543_ cpu.IO_addr_buff\[2\] _01049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08262_ _03504_ _00276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05474_ _00981_ _00982_ _00869_ _00983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07698__I _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07213_ cpu.timer_capture\[0\] _02674_ _02681_ _02662_ _02682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_74_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08028__A2 _01962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08193_ _03449_ _03342_ _03451_ _03452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_54_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06039__A1 _00997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07144_ _00752_ _02621_ _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07075_ _02562_ _02563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06026_ cpu.timer_div\[2\] _01407_ _01527_ _01529_ _01182_ _01530_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_65_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06211__A1 net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07977_ cpu.spi.data_in_buff\[3\] _03270_ _03272_ cpu.spi.data_in_buff\[2\] _03276_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09716_ _04735_ _00499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_58_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06928_ _02407_ _02408_ _02424_ _02404_ _02425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_96_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09647_ cpu.last_addr\[13\] _04654_ _04660_ _04678_ _04679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_06859_ _00621_ _01956_ _02357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_2_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09578_ _04609_ _04611_ _04612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08529_ cpu.toggle_ctr\[8\] _03715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_93_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10422_ _00361_ clknet_leaf_15_wb_clk_i cpu.pwm_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10353_ _00292_ clknet_leaf_36_wb_clk_i cpu.uart.receive_div_counter\[12\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09519__A2 _00771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10284_ _00223_ clknet_leaf_64_wb_clk_i cpu.spi.data_in_buff\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09772__B _03897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08388__B _03570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07702__A1 _01373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09058__I1 _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05190_ _00726_ _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06371__B _01379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06292__I1 cpu.regs\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07900_ cpu.spi.div_counter\[5\] _03214_ _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08880_ _03982_ _00416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07831_ _03139_ cpu.timer\[13\] _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05547__A3 _01052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_16_Left_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05398__I3 cpu.regs\[11\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09501_ _04488_ _04524_ _04537_ _04511_ _04538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07762_ _02076_ _02391_ _03091_ _03092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_79_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07693_ _03011_ cpu.regs\[4\]\[6\] _03026_ _03036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06713_ _02209_ _02210_ _02211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_69_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09432_ _02587_ _04028_ _04471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06644_ _00621_ _00996_ _02141_ _02142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_82_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09363_ _04346_ _04400_ _04404_ _04405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06575_ _02072_ _02073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08314_ _02826_ _03537_ _03544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_47_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05526_ _00656_ _01030_ _01031_ _01032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_35_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09294_ _00764_ _04338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_25_Left_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08245_ _02873_ _03288_ _00271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05457_ _00907_ _00967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08176_ _03425_ _03438_ _00256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_105_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05388_ _00873_ _00900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_7_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05322__I3 cpu.regs\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07127_ _02527_ _02610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_70_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09148__I _04194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06432__A1 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07058_ _02076_ _02547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06009_ _01511_ _01512_ _01215_ _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_100_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_34_Left_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06196__B1 _01698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06291__S0 _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_qcpu_105 io_oeb[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__06499__A1 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09437__A1 _04209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_43_Left_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07131__I _02531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10405_ _00344_ clknet_leaf_4_wb_clk_i cpu.toggle_ctr\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05226__A2 _00761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10336_ _00275_ clknet_leaf_45_wb_clk_i cpu.uart.receive_buff\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_52_Left_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10267_ _00206_ clknet_leaf_28_wb_clk_i cpu.spi.div_counter\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08176__A1 _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10198_ _00137_ clknet_leaf_118_wb_clk_i cpu.regs\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_105_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07750__B _03064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_61_Left_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_75_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06360_ _01860_ _01861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06291_ cpu.regs\[4\]\[6\] cpu.regs\[5\]\[6\] cpu.regs\[6\]\[6\] cpu.regs\[7\]\[6\]
+ _00888_ _00889_ _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_05311_ cpu.regs\[8\]\[2\] cpu.regs\[9\]\[2\] cpu.regs\[10\]\[2\] cpu.regs\[11\]\[2\]
+ _00569_ _00574_ _00842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08030_ _02629_ _03316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput30 sram_out[4] net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05242_ _00711_ _00778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_5_0_wb_clk_i clknet_0_wb_clk_i clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__09600__A1 _04209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05173_ cpu.base_address\[5\] _00710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05496__I _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09981_ _02476_ _04945_ _02479_ _02486_ _04946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__05217__A2 _00658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08932_ _04022_ _04015_ _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08863_ cpu.spi.divisor\[7\] _03966_ _03970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07814_ cpu.timer_div\[6\] _03133_ cpu.timer_div_counter\[7\] _01976_ _03134_ _03135_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_08794_ cpu.timer_capture\[15\] _03843_ _03915_ _03916_ _03917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06120__I _01197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_16_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07745_ _02376_ _03076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09415_ _00740_ _04455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07676_ _02997_ _03017_ _03025_ _00169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06627_ _02123_ _02124_ _02125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06558_ cpu.mem_cycle\[3\] _02056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_74_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09346_ _02381_ _01430_ _04388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09277_ _04309_ _04321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06489_ _01021_ _01278_ _01432_ _01957_ _01791_ _01988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_7_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05509_ _01016_ _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08228_ _02652_ _03476_ _03480_ _03481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06790__I _00822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08159_ _00792_ _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06405__B2 _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10121_ _00064_ clknet_leaf_19_wb_clk_i cpu.timer_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_55_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output68_I net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10052_ _05012_ _05013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05067__S1 _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05782__I3 cpu.regs\[3\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06644__A1 _00621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06205__I _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10319_ _00258_ clknet_leaf_40_wb_clk_i cpu.uart.counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_111_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05860_ _01365_ _01366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_28_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05791_ _01146_ _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_37_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07530_ _02934_ _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_66_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07461_ _02071_ _02889_ _02890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07392_ _02824_ _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_91_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09200_ cpu.orig_PC\[0\] _04244_ _04245_ _04181_ _04246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_56_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06412_ _00630_ _01799_ _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09131_ _04179_ _04180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06343_ _01840_ _01843_ _01844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09821__A1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09062_ cpu.regs\[3\]\[3\] _03090_ _04117_ _04128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06274_ net94 _01775_ _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08013_ cpu.uart.receive_buff\[5\] _03302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_69_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_25_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_25_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05225_ _00752_ _00660_ _00760_ _00761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_05156_ _00669_ _00694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_77_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09964_ net65 _04922_ _04924_ _04931_ _03122_ _04932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_05087_ _00623_ _00627_ _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09888__A1 _04823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09895_ _04864_ _04877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08915_ _04009_ _00424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08846_ _03958_ _03960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05049__S1 _00575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08560__A1 _03738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08777_ cpu.timer_capture\[12\] _03883_ _03897_ _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05989_ _01493_ _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07728_ _01308_ _01371_ _02401_ _03061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07659_ _03015_ _03016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08933__C _04020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09329_ _04357_ _04371_ _04372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_11_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05429__A2 _00939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10104_ _00047_ clknet_leaf_32_wb_clk_i cpu.uart.divisor\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09780__B _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10035_ _01332_ _04997_ _04998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07106__A2 _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05117__A1 cpu.base_address\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05668__A2 _01111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07520__S _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07290__A1 _02665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06363__C _00720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05840__A2 _01345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06961_ _02449_ _02450_ _02041_ _02454_ _02455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_09680_ _02038_ _02039_ _04706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08700_ cpu.timer\[0\] _03837_ _03838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05912_ cpu.pwm_top\[1\] _01254_ _01255_ _01417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08631_ cpu.pwm_top\[3\] _03787_ _03789_ _03783_ _03790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06892_ cpu.PC\[11\] _02389_ _02390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_89_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05843_ _01347_ _01348_ _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_89_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08562_ _03699_ _03739_ _03742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05774_ _00707_ _01120_ _01280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08493_ cpu.toggle_ctr\[10\] _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07513_ cpu.regs\[12\]\[2\] _02919_ _02924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07444_ _02845_ _02864_ _02876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07375_ _02325_ _02330_ _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08325__I _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09114_ cpu.last_addr\[9\] _04157_ _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_79_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06326_ cpu.toggle_top\[13\] _01106_ _01827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09045_ _04113_ _04114_ _04115_ _04116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07281__A1 _02648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06257_ _00598_ _01758_ _01759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_103_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05208_ _00687_ _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06188_ _01591_ _01682_ _01691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05684__I cpu.spi.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05139_ cpu.IO_addr_buff\[7\] cpu.IO_addr_buff\[6\] cpu.IO_addr_buff\[5\] _00678_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XPHY_EDGE_ROW_8_Left_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09947_ _02052_ _02483_ _04916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07584__A2 _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09878_ _01122_ _04812_ _04864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_99_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08829_ _03904_ _03922_ _03945_ _03946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_68_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05859__I _00656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10584_ _00522_ clknet_leaf_68_wb_clk_i net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_63_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07647__I0 _03007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07024__A1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10018_ _01269_ _01265_ _04223_ _02721_ _04221_ _04981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_98_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07314__I _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05490_ _00992_ _00998_ _00959_ _00999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07160_ _02633_ _02637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06111_ cpu.PORTA_DDR\[3\] _01613_ _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_81_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07263__A1 cpu.timer_capture\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07091_ _02570_ _02572_ _02577_ _02578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06042_ _00794_ _01297_ _01544_ _01545_ _01546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_2_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07015__A1 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09801_ cpu.pwm_top\[3\] cpu.pwm_counter\[3\] _04805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07993_ _03286_ _03287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09732_ _02495_ _04749_ _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_5_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06944_ _02427_ _02438_ _02439_ _00023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09663_ _04691_ _02538_ _04692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06875_ _02077_ _02371_ _02372_ _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08614_ _03768_ _03776_ _00356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09594_ _04597_ _00952_ _04627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05826_ _01331_ _01332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07224__I _02673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08545_ cpu.toggle_clkdiv cpu.toggle_ctr\[1\] cpu.toggle_ctr\[0\] _03730_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_49_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05757_ _01262_ _01263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05688_ _00683_ _01194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_65_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08476_ _03653_ _03666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07427_ cpu.uart.receive_div_counter\[5\] _02860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06284__B _01380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_40_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_40_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_73_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07629__I0 _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07358_ _02797_ _02409_ _02798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06309_ net3 _01389_ _01807_ _01809_ _01108_ _01810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_103_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07289_ _02736_ _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09028_ _00837_ _02810_ _04102_ _04103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08754__A1 cpu.timer_capture\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output50_I net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05740__A1 _01063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07245__A1 _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10567_ _00505_ clknet_leaf_75_wb_clk_i cpu.ROM_spi_dat_out\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10498_ _00436_ clknet_leaf_55_wb_clk_i cpu.IO_addr_buff\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08993__A1 _01877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput6 io_in[14] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_108_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06660_ _02156_ _02157_ _02158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09170__A1 _00590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05611_ _01116_ _01117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_86_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05731__A1 cpu.timer_capture\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06591_ _00589_ _01956_ _02089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08330_ cpu.uart.receive_div_counter\[12\] _03554_ _03548_ _03557_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_86_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05542_ _01047_ _01048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_47_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08261_ cpu.uart.receive_buff\[5\] _03503_ _03497_ cpu.uart.receive_buff\[4\] _03504_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_86_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05473_ cpu.regs\[0\]\[4\] cpu.regs\[1\]\[4\] cpu.regs\[2\]\[4\] cpu.regs\[3\]\[4\]
+ _00877_ _00977_ _00982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_22_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07212_ _02675_ _02677_ _02678_ _02680_ _02681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08192_ _03450_ _03451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_89_Left_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_70_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07143_ _02595_ _02622_ _02623_ _02618_ _00038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_14_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07074_ cpu.PC\[5\] _02562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06025_ _01528_ _01383_ _01407_ _01529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__05448__B _00933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07219__I _02661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07976_ _03275_ _00219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09715_ _02457_ _04732_ _04733_ _04734_ _04735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XPHY_EDGE_ROW_98_Left_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_87_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06927_ _02423_ _02409_ _02424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09646_ _04662_ _04663_ _04664_ _04677_ _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__09161__A1 _01429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06279__B _01479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05970__A1 _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06858_ _00638_ _01017_ _02356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_2_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09577_ _04353_ _04599_ _04610_ _04356_ _04611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06789_ _00820_ _00849_ _00893_ _00953_ _02287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_05809_ _01313_ _01314_ _01315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_92_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08528_ _03697_ cpu.toggle_top\[7\] _03713_ _03714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08459_ _01052_ _02747_ _03653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_107_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10421_ _00360_ clknet_leaf_15_wb_clk_i cpu.pwm_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10352_ _00291_ clknet_leaf_36_wb_clk_i cpu.uart.receive_div_counter\[11\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10283_ _00222_ clknet_leaf_64_wb_clk_i cpu.spi.data_in_buff\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07292__C _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09152__A1 _04196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05713__A1 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07799__I _02735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06208__I cpu.uart.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05112__I net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10619_ _00557_ clknet_leaf_66_wb_clk_i net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_113_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08423__I _03595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06292__I2 cpu.regs\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07830_ _03146_ _03149_ _03150_ _03151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07761_ _03090_ _02389_ _03091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09500_ _04530_ _04534_ _04536_ _04537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06712_ _00589_ _00994_ _02210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05952__A1 _00920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07692_ _03035_ _00175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_69_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09431_ _00777_ _04468_ _04469_ _04470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06643_ _02138_ _02139_ _02141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09362_ _02530_ _04384_ _04402_ _04378_ _04403_ _04404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_47_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06574_ _02071_ _02067_ _02072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_08313_ cpu.uart.receive_div_counter\[9\] _03543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05525_ _00778_ _00741_ _01029_ _01031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_35_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09293_ _02078_ _04334_ _04336_ _04337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05307__I1 _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08244_ _03120_ _03451_ _03492_ _00270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_62_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05456_ _00964_ _00965_ _00897_ _00966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08175_ cpu.uart.has_byte _03437_ _03289_ _03438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05387_ _00898_ _00899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__08957__B2 _01022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07126_ _02607_ _02603_ _02609_ _02606_ _00035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__10064__I0 _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05957__I _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_45_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08709__A1 _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07057_ _02541_ _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06008_ net41 _01385_ _01512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_7_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05692__I _01197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07959_ cpu.spi.data_out_buff\[5\] _03231_ _03263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09134__A1 _00728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06291__S1 _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08936__C _04020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09629_ cpu.last_addr\[8\] _04651_ _04661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xwrapped_qcpu_106 io_oeb[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__06499__A2 _01997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_84_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10404_ _00343_ clknet_leaf_5_wb_clk_i cpu.toggle_ctr\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05867__I _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10335_ _00274_ clknet_leaf_45_wb_clk_i cpu.uart.receive_buff\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10266_ _00205_ clknet_leaf_33_wb_clk_i cpu.spi.div_counter\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10197_ _00136_ clknet_leaf_112_wb_clk_i cpu.regs\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05934__A1 cpu.br_rel_dest\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05107__I _00646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07439__A1 _00788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07322__I _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06111__A1 cpu.PORTA_DDR\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06290_ _01300_ _01140_ _01791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_05310_ _00586_ _00840_ _00841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput20 io_in[3] net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_116_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput31 sram_out[5] net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05241_ _00776_ _00777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09249__I _04292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05172_ cpu.base_address\[4\] _00709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_116_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09980_ _04640_ _02055_ _04945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08931_ _02715_ _04022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_110_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08862_ _02665_ _03965_ _03969_ _00411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_4_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07813_ _03128_ cpu.timer_div_counter\[2\] _03133_ cpu.timer_div\[6\] _03134_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08793_ _03794_ _03916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_74_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07744_ _02350_ _03074_ _02409_ _03075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07675_ cpu.regs\[5\]\[7\] _03015_ _03025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09414_ _04294_ _04433_ _04453_ _04331_ _04454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_48_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06626_ _02079_ _02080_ _02124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_109_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06557_ _02054_ _02055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_47_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09345_ _04385_ _04386_ _04387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_118_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09276_ _04316_ _04296_ _04318_ _04319_ _04320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06488_ _01423_ _01986_ _01987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_7_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05508_ _01015_ _01016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_35_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08227_ cpu.uart.data_buff\[6\] _03458_ _03480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05439_ _00718_ _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_90_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05861__B1 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_1_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08158_ _03423_ _03424_ _00252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08063__I _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08089_ _00727_ _03366_ _03367_ _00767_ _03368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
X_07109_ _02594_ _00033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_101_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10120_ _00063_ clknet_leaf_20_wb_clk_i cpu.timer_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10051_ _05011_ _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06169__A1 _00973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05916__A1 cpu.toggle_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10318_ _00257_ clknet_leaf_21_wb_clk_i cpu.uart.counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07518__S _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10249_ _00188_ clknet_leaf_103_wb_clk_i cpu.regs\[2\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05790_ _01285_ _01295_ _01296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_37_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07460_ _01145_ _01163_ _02888_ _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__09688__B _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07391_ cpu.uart.divisor\[12\] _02824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_60_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06411_ _00631_ _01840_ _01911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08085__A1 _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09130_ _01142_ _01154_ _00707_ _01279_ _04179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_06342_ _01841_ _01842_ _01843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09061_ _04127_ _00452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08012_ _03300_ _03298_ _03301_ _03296_ _00229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__07832__A1 cpu.timer_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06273_ _01693_ _01761_ _01775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05224_ _00759_ _00760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05300__I _00831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05155_ _00692_ _00693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06399__A1 _01879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09963_ _04926_ _04928_ _04930_ _04931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_77_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05086_ cpu.regs\[8\]\[6\] cpu.regs\[9\]\[6\] cpu.regs\[10\]\[6\] cpu.regs\[11\]\[6\]
+ _00617_ _00618_ _00627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07060__A2 _02385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_65_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_65_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08914_ cpu.uart.divisor\[10\] _04001_ _04008_ _04006_ _04009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_90_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09894_ _04864_ _04876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08845_ _03958_ _03959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08776_ cpu.timer\[12\] _03811_ _03841_ _03901_ _03902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08560__A2 _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input12_I io_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07727_ net1 _03054_ _03059_ _02074_ _03060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_05988_ _01381_ _01436_ _01491_ _01492_ _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_95_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07658_ _03014_ _03015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06609_ _02105_ _02106_ _02107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07589_ _02969_ _02970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09328_ _04363_ _04369_ _04370_ _04371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_80_Left_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09259_ cpu.PC\[2\] cpu.br_rel_dest\[2\] _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__05210__I _00746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09576__A1 cpu.orig_PC\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10103_ _00046_ clknet_leaf_31_wb_clk_i cpu.uart.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10034_ _04986_ _02013_ _04997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05880__I _01112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08067__A1 _03347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07814__B2 _01976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07814__A1 cpu.timer_div\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05428__I0 cpu.regs\[8\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07042__A2 _02531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06960_ _02452_ _02453_ _02454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA_input4_I io_in[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05911_ cpu.timer_top\[9\] _01175_ _01179_ _01416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06891_ cpu.PC\[10\] _02376_ _02388_ _02389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_08630_ _02758_ _03788_ _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05842_ _00716_ _01348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_89_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08561_ _03741_ _00338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05773_ _01040_ _01279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__06305__A1 net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08492_ cpu.toggle_ctr\[9\] _03677_ _01261_ cpu.toggle_ctr\[8\] _03678_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07512_ _01602_ _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07443_ cpu.uart.receive_counter\[0\] cpu.uart.receive_counter\[1\] _02865_ _02875_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_77_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07711__S _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_112_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_112_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_91_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09113_ cpu.ROM_addr_buff\[9\] _04159_ _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09211__B _04256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07374_ _02810_ _02796_ _02811_ _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_79_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06325_ cpu.toggle_top\[5\] _01643_ _01825_ _01257_ _01826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_88_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09044_ _03997_ _04115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_45_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06256_ _01757_ _01665_ _01662_ _01758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05207_ _00732_ _00737_ _00743_ _00744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09558__A1 _00851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06187_ _01670_ _01688_ _01480_ _01690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05138_ cpu.IO_addr_buff\[4\] _00677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__07033__A2 _02524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09946_ _02045_ _00733_ _04915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08781__A2 _03811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05069_ cpu.regs\[8\]\[5\] cpu.regs\[9\]\[5\] cpu.regs\[10\]\[5\] cpu.regs\[11\]\[5\]
+ _00600_ _00601_ _00611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09877_ _04863_ _00532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_79_Right_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08828_ _02708_ _03923_ _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08759_ _03885_ _03865_ _03866_ _03887_ _03881_ _03888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_95_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_109_Left_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10583_ _00521_ clknet_leaf_68_wb_clk_i net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_106_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_88_Right_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06036__I _00930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05875__I _01379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_118_Left_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07024__A2 _02516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07575__A3 _01153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05586__A2 _00655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_97_Right_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10017_ cpu.orig_flags\[0\] _04032_ _04977_ _04979_ _04980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_47_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08288__B2 _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09788__A1 _03227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06110_ _00674_ _00679_ _01243_ _01613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_07090_ _02573_ _02575_ _02576_ _02577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06041_ _00920_ _01432_ _01146_ _01545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_23_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07992_ _02876_ _03285_ _03286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09960__B2 cpu.ROM_addr_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09960__A1 cpu.ROM_addr_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09800_ _03763_ _04804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09731_ _04747_ _04748_ _04749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_66_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06943_ _01950_ _02401_ _02402_ cpu.regs\[2\]\[6\] _02439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_09662_ _02056_ _04691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06874_ _02166_ _02352_ _02370_ _02372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__06526__A1 _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07505__I _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08613_ cpu.pwm_counter\[7\] _03774_ _03776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09593_ _04597_ _00951_ _04626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05825_ _00657_ _01330_ _01331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08279__A1 _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08544_ _03725_ _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05756_ _01106_ _01262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_85_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05687_ _01100_ _01193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08475_ _03665_ _00328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_49_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07426_ _02856_ cpu.uart.receive_div_counter\[13\] _02835_ _02629_ _02858_ _02859_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_18_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07357_ _02796_ _02797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06308_ _01217_ _01808_ _01809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_80_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_80_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07288_ cpu.timer_top\[6\] _02740_ _02743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09027_ _04101_ _04102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__05695__I _01200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06239_ _01004_ _01353_ _01740_ _01350_ _01356_ _01741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_32_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09951__A1 net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09929_ _04902_ _00545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07415__I cpu.uart.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output43_I net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07565__I0 _02943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05879__I0 cpu.PORTA_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08690__A1 _02665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07150__I _02617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10566_ _00504_ clknet_leaf_76_wb_clk_i cpu.ROM_spi_dat_out\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10290__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10497_ _00435_ clknet_leaf_55_wb_clk_i cpu.IO_addr_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput7 io_in[15] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06508__A1 _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07325__I _02771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09170__A2 _02361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05610_ cpu.IO_addr_buff\[4\] _01115_ _01055_ _01116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_59_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06590_ _02086_ _02087_ _02088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05541_ _01046_ _01047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_74_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08260_ _03493_ _03503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08681__A1 _02648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05472_ cpu.regs\[4\]\[4\] cpu.regs\[5\]\[4\] cpu.regs\[6\]\[4\] cpu.regs\[7\]\[4\]
+ _00877_ _00977_ _00981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_116_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08191_ _03376_ _03323_ _03338_ _03450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_07211_ _01023_ _02679_ _02680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07142_ _01704_ _02621_ _02623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07073_ _02548_ _02561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_35_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06024_ cpu.spi.dout\[2\] _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_100_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07975_ cpu.spi.data_in_buff\[2\] _03270_ _03272_ cpu.spi.data_in_buff\[1\] _03275_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09714_ _02457_ _04729_ _00689_ _04734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_87_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07547__I0 _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06926_ _02410_ _02422_ _02423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09645_ _04114_ _04666_ _04675_ _04676_ _04677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_06857_ _02091_ _02092_ _02354_ _02355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05808_ _00717_ _00719_ _01314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09576_ cpu.orig_PC\[12\] _04354_ _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06788_ _02285_ _02281_ _02286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10059__A1 _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05739_ cpu.timer_capture\[8\] _01242_ _01244_ _01245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08527_ _03700_ _03711_ _03712_ _03713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08458_ _03652_ _00747_ _00324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_74_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07409_ _02840_ cpu.uart.receive_div_counter\[15\] _02841_ cpu.uart.divisor\[3\]
+ _02842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08389_ cpu.orig_flags\[0\] _03587_ _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10420_ _00359_ clknet_leaf_14_wb_clk_i cpu.pwm_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07838__C cpu.timer_top\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10351_ _00290_ clknet_leaf_37_wb_clk_i cpu.uart.receive_div_counter\[10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10282_ _00221_ clknet_leaf_49_wb_clk_i cpu.spi.data_in_buff\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07163__A1 _02629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05713__A2 _01215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07081__S _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10618_ _00556_ clknet_leaf_99_wb_clk_i cpu.C vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10549_ _00487_ clknet_leaf_72_wb_clk_i cpu.mem_cycle\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_51_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09915__A1 _04819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_119_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07760_ _03089_ _03090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06711_ _02208_ _00928_ _02207_ _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09430_ _04413_ _04462_ _04469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07691_ _03009_ cpu.regs\[4\]\[5\] _03026_ _03035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_69_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09270__I _04313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06642_ _00972_ _02138_ _02139_ _02140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__06901__A1 _01788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09361_ _04194_ _04403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06573_ _02066_ _02071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08312_ _03522_ _03542_ _00288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_82_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_19_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_19_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_59_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09292_ _04335_ _04297_ _04336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05524_ _00714_ _01029_ _01030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08243_ _03109_ _03368_ cpu.uart.data_buff\[9\] _03492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05307__I2 _00837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05455_ cpu.regs\[0\]\[3\] cpu.regs\[1\]\[3\] cpu.regs\[2\]\[3\] cpu.regs\[3\]\[3\]
+ _00962_ _00963_ _00965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08174_ cpu.uart.clr_hb _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_103_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05386_ _00878_ _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07125_ _02608_ _02602_ _02609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07056_ _01787_ _02545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06007_ _01507_ _01508_ _01510_ _01511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09906__A1 _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09445__I _00689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07958_ _03262_ _00214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07889_ cpu.spi.div_counter\[1\] _03205_ _03208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06909_ _02405_ _02406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_97_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09628_ _04169_ cpu.ROM_addr_buff\[10\] _04652_ _04660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08893__A1 _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_qcpu_107 io_oeb[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_54_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09559_ _04256_ _04571_ _04593_ _04339_ _04594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_77_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10403_ _00342_ clknet_leaf_6_wb_clk_i cpu.toggle_ctr\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05369__B _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10334_ _00273_ clknet_leaf_67_wb_clk_i cpu.uart.receive_buff\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05631__A1 _01130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07620__A2 _02986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10265_ _00204_ clknet_leaf_33_wb_clk_i cpu.spi.div_counter\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07584__B _02967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09373__A2 _00756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10196_ _00135_ clknet_leaf_113_wb_clk_i cpu.regs\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05785__I2 cpu.regs\[10\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09090__I _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07439__A2 _02871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08636__A1 _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput10 io_in[18] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput21 io_in[6] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05240_ _00775_ _00776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput32 sram_out[6] net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05171_ _00707_ _00708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_116_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08930_ _04021_ _00427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05793__I _01269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08861_ cpu.spi.divisor\[6\] _03966_ _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07812_ cpu.timer_div_counter\[6\] _03133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_4_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08792_ _03180_ _03914_ _03845_ _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07743_ _02234_ _02348_ _02349_ _03074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__08875__A1 _02692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07674_ _03024_ _00168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09413_ _04443_ _04450_ _04452_ _04453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06625_ _02120_ _02121_ _02123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_59_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06350__A2 _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06556_ _02053_ cpu.mem_cycle\[4\] _02054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05033__I _00575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09344_ cpu.PC\[3\] _01138_ _04360_ _04386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06487_ _01268_ _01957_ _01985_ _01986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09275_ _04269_ _04319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05507_ _01014_ _01015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_105_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08226_ _03479_ _00265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05438_ _00948_ net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08157_ _03324_ _03421_ _03237_ _03424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_95_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09052__A1 _02378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07108_ _02418_ _02593_ _02543_ _02594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05369_ _00006_ _00880_ _00007_ _00881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_08088_ _00681_ _03367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_30_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05613__A1 _01114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07039_ _02529_ _00028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_100_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10050_ _02889_ _02932_ _05011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09108__C _03980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05208__I _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05472__S0 _00877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05652__B _01157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07423__I cpu.uart.divisor\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06341__A2 _01758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08618__A1 _02636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05852__A1 _00868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10317_ _00256_ clknet_leaf_42_wb_clk_i cpu.uart.has_byte vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05455__I1 cpu.regs\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09346__A2 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10248_ _00187_ clknet_leaf_106_wb_clk_i cpu.regs\[2\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09813__I _01429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10179_ _00118_ clknet_leaf_123_wb_clk_i cpu.regs\[11\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08857__A1 cpu.spi.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05135__A3 _00661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06410_ _01306_ _01909_ _01910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07390_ cpu.uart.receive_counter\[0\] _02823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_45_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06341_ _00598_ _01758_ _01842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09060_ _04125_ cpu.ROM_addr_buff\[10\] _04126_ _04127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_71_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06272_ _01739_ _01693_ _01761_ _01774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_08011_ cpu.uart.dout\[4\] _03294_ _03301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_72_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05223_ _00753_ _00758_ _00759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_71_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05154_ _00691_ _00692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09962_ _04929_ _04930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_77_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05085_ _00587_ _00625_ _00626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08913_ _02754_ _04002_ _04008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_90_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09893_ _04875_ _00536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08844_ _03232_ _03367_ _01067_ _02746_ _03958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__05028__I _00570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08775_ _03832_ _03899_ _03900_ _03901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05987_ _01379_ _01492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xclkbuf_leaf_34_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_34_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07726_ _03056_ _03058_ _03054_ _03059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08848__A1 _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07657_ _01137_ _02982_ _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_94_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06608_ _02088_ _02089_ _02106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07588_ _02968_ _02969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09327_ _00762_ _04370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_48_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06539_ _02036_ _02037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_90_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09258_ _04300_ _04275_ _04301_ _04302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08209_ _02635_ _03455_ _03465_ _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09189_ _01311_ _00709_ _04234_ _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_16_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07587__A1 _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output73_I net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10102_ _00045_ clknet_leaf_31_wb_clk_i cpu.uart.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_101_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08000__A2 _03288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10033_ _01992_ _04992_ _04994_ _04995_ _04996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__07153__I _01091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05401__I _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09016__A1 _00992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05053__A2 _00582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06250__A1 net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09971__C _03347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05910_ cpu.timer_top\[1\] _01382_ _01410_ _01412_ _01414_ _01415_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_06890_ _02378_ _02387_ _02388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05841_ _01312_ _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08159__I _00792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08560_ _03738_ _03724_ _03739_ _03740_ _03741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_05772_ _01277_ _01278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_89_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08491_ cpu.toggle_top\[9\] _03677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07502__A1 _01130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07511_ _02921_ _02918_ _02922_ _00107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07442_ _02823_ _02865_ _02874_ _00086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07373_ _02382_ _02811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09112_ _03812_ _04166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06324_ _01171_ _01823_ _01824_ _01825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_45_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06069__A1 _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06069__B2 _01452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09043_ cpu.ROM_addr_buff\[6\] _04114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06255_ _01139_ net93 _01757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_111_Right_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05206_ _00704_ _00734_ _00742_ _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06186_ _01658_ _01688_ _01689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05137_ cpu.IO_addr_buff\[3\] _00676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07569__A1 cpu.regs\[10\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09945_ _04910_ _02455_ _02482_ _04914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05068_ _00587_ _00609_ _00610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09876_ net58 _04853_ _04862_ _04858_ _04863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09030__I1 cpu.ROM_addr_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08518__B1 _01498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08827_ _03944_ _00401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08758_ _03885_ _03886_ _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_68_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08689_ cpu.timer_top\[14\] _03825_ _03829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09494__A1 _03637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07709_ _03007_ cpu.regs\[3\]\[4\] _03039_ _03046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_95_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09246__A1 _02797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10582_ _00520_ clknet_leaf_69_wb_clk_i net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_63_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06480__A1 cpu.timer_capture\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06232__B2 _00973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05586__A3 _01091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09021__I1 cpu.ROM_addr_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10016_ _02614_ _02109_ _04217_ _04978_ _04979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06535__A2 _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09485__A1 _03065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07611__I _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05897__I1 cpu.spi.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09237__A1 _04281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06471__A1 _01962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08442__I _03595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_25_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06040_ _01423_ _01541_ _01543_ _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07058__I _02076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07991_ cpu.uart.receiving _03284_ _03285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09730_ _00691_ _02492_ _04748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_66_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06942_ _02406_ _02436_ _02437_ _02438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09173__B1 _04180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09661_ _00746_ _04689_ _04690_ _00489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06873_ _02166_ _02352_ _02370_ _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_08612_ _03773_ _03775_ _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09592_ _03649_ _00772_ _04505_ _04624_ _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05824_ _01314_ _01330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08543_ _03727_ _03728_ _00333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05755_ cpu.toggle_top\[8\] _01261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_106_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05686_ _01190_ _01191_ _01189_ _01192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08474_ cpu.toggle_top\[3\] _03654_ _03664_ _03660_ _03665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_18_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07425_ _02857_ cpu.uart.receive_div_counter\[10\] _02849_ _02848_ _02858_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_clkbuf_leaf_64_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07356_ _02795_ _02796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06307_ net64 _01514_ _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07287_ _02658_ _02739_ _02742_ _02737_ _00063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_115_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09026_ _00700_ _04101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06238_ _00596_ _01003_ _01740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_103_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06169_ _00973_ _01352_ _01656_ _01340_ _01355_ _01672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06214__A1 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09928_ cpu.PORTA_DDR\[4\] _04899_ _04901_ _04893_ _04902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09859_ _04850_ _00527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_output36_I net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10565_ _00503_ clknet_leaf_75_wb_clk_i cpu.ROM_spi_dat_out\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10496_ _00434_ clknet_leaf_56_wb_clk_i cpu.IO_addr_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_109_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput8 io_in[16] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07705__A1 cpu.regs\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09170__A3 _02416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05540_ _00677_ _00678_ _01046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10068__A2 _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05471_ _00978_ _00979_ _00869_ _00980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08190_ cpu.uart.counter\[2\] _03449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07210_ _02676_ _02679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07141_ _02621_ _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05796__I _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07072_ _02386_ _02560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06023_ _01525_ _01526_ _01189_ _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_2_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07974_ _03274_ _00218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09713_ _04727_ _04724_ _04723_ _04733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_87_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06925_ _02412_ _02421_ _02422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09644_ cpu.last_addr\[5\] cpu.ROM_addr_buff\[5\] _04649_ _04676_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__09161__A3 _02668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06856_ _02093_ _02094_ _02354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_93_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05807_ _01312_ _00716_ _01313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05036__I _00002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09575_ _00763_ _04604_ _04608_ _04609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06787_ _02266_ _02271_ _02285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05738_ _01243_ _01104_ _01244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08526_ _03697_ cpu.toggle_top\[7\] _03712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05669_ _01174_ _01175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08457_ cpu.toggle_clkdiv _03652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_37_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07408_ cpu.uart.receive_div_counter\[3\] _02841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_18_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08388_ _03601_ _03602_ _03570_ _00304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_61_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07339_ _02542_ _02780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_33_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10350_ _00289_ clknet_leaf_36_wb_clk_i cpu.uart.receive_div_counter\[9\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05238__A2 _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06435__B2 _01451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10281_ _00220_ clknet_leaf_47_wb_clk_i cpu.spi.data_in_buff\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09009_ _03987_ _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_14_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08188__B2 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07627__S _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06294__S0 _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08112__A1 _00793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09860__A1 _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06674__A1 _02168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10617_ _00555_ clknet_leaf_74_wb_clk_i net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10548_ _00486_ clknet_leaf_84_wb_clk_i cpu.PC\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_52_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10479_ _00418_ clknet_leaf_20_wb_clk_i cpu.timer_div\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_71_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06710_ _00620_ _00927_ _02208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07690_ _03034_ _00174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_87_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06641_ _00620_ _00954_ _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_63_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09360_ _00590_ _04334_ _04401_ _04402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06572_ _02069_ _02070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08311_ _02826_ _03511_ _03540_ _03541_ _03542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_82_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09291_ _04252_ _04335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05523_ _01028_ _01029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_35_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08242_ _02606_ _03490_ _03491_ _00269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05454_ cpu.regs\[4\]\[3\] cpu.regs\[5\]\[3\] cpu.regs\[6\]\[3\] cpu.regs\[7\]\[3\]
+ _00962_ _00963_ _00964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05307__I3 cpu.regs\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08173_ _03425_ _03436_ _00255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_103_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05385_ _00886_ _00897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_6_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07124_ _01035_ _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07055_ _02543_ _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06006_ _01509_ _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_100_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07917__A1 _00746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07957_ cpu.spi.data_out_buff\[5\] _03255_ _03261_ _03258_ _03262_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06908_ _02035_ _02405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08342__A1 _02871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07888_ cpu.spi.div_counter\[1\] _03205_ _03207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09627_ cpu.last_addr\[11\] cpu.ROM_addr_buff\[11\] _04653_ _04659_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_54_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06839_ _02335_ _02336_ _02337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xwrapped_qcpu_108 io_out[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09558_ _00851_ _04515_ _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08509_ _03689_ _03692_ _03694_ _03695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09489_ _04497_ _04498_ _04525_ _04526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_53_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_12_Left_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10402_ _00341_ clknet_leaf_5_wb_clk_i cpu.toggle_ctr\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06408__A1 _01018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10333_ _00272_ clknet_leaf_67_wb_clk_i cpu.uart.receive_buff\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10264_ _00203_ clknet_leaf_33_wb_clk_i cpu.spi.div_counter\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10195_ _00134_ clknet_leaf_111_wb_clk_i cpu.regs\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05785__I3 cpu.regs\[11\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_21_Left_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_105_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06195__I0 net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09833__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06647__A1 cpu.regs\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput11 io_in[19] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput22 io_in[7] net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput33 sram_out[7] net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05170_ _00706_ _00707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_12_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08860_ _02658_ _03965_ _03968_ _00410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07811_ cpu.timer_div\[1\] _03125_ _03126_ cpu.timer_div\[5\] _03131_ _03132_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_4_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_106_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_106_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_74_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08791_ cpu.timer\[15\] _03913_ _03914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07742_ _03073_ _00187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07673_ _03011_ cpu.regs\[5\]\[6\] _03014_ _03024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09412_ _04324_ _04433_ _04451_ _04327_ _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06624_ _02120_ _02121_ _02122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10079__D _00022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09343_ _02382_ _01138_ _04385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09824__A1 _04823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06555_ _02052_ _02053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_118_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09274_ _02802_ _04317_ _04318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06486_ _01271_ _01958_ _01983_ _01984_ _01267_ _01985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_05506_ _01010_ _01013_ _00883_ _01014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08225_ cpu.uart.data_buff\[4\] _03475_ _03478_ _03467_ _03479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05437_ _00925_ _00933_ _00947_ _00948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_7_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08156_ _03324_ _03383_ _03422_ _03390_ _03423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_99_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05368_ cpu.regs\[4\]\[0\] cpu.regs\[5\]\[0\] cpu.regs\[6\]\[0\] cpu.regs\[7\]\[0\]
+ _00878_ _00879_ _00880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_15_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07063__A1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07107_ _02546_ _02591_ _02592_ _02593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_113_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08087_ _00650_ _03366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05299_ _00566_ _00825_ _00830_ _00831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_07038_ _00780_ _02514_ _02528_ _02522_ _02529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_101_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08989_ cpu.IO_addr_buff\[5\] _04066_ _04072_ _04069_ _04073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05472__S1 _00977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09815__A1 _04815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_4_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_4_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10316_ _00255_ clknet_leaf_38_wb_clk_i cpu.uart.div_counter\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_21_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05455__I2 cpu.regs\[2\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10247_ _00186_ clknet_leaf_106_wb_clk_i cpu.regs\[2\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07601__I0 _02943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_111_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10178_ _00117_ clknet_leaf_125_wb_clk_i cpu.regs\[11\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08306__A1 _03495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05134__I _00672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05391__I1 cpu.regs\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06340_ _00614_ _01841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07293__A1 _01091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06271_ _01769_ _01772_ _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08010_ cpu.uart.receive_buff\[4\] _03300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05222_ _00755_ _00757_ _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05153_ _00665_ _00668_ _00691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_69_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09961_ _00665_ _04929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_77_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05084_ cpu.regs\[12\]\[6\] cpu.regs\[13\]\[6\] cpu.regs\[14\]\[6\] cpu.regs\[15\]\[6\]
+ _00600_ _00601_ _00625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08912_ _04007_ _00423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_90_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09892_ cpu.PORTB_DDR\[3\] _04865_ _04874_ _04870_ _04875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_85_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08843_ _03957_ _00404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_109_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08774_ _03894_ _03890_ cpu.timer\[12\] _03900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05986_ _01309_ _01489_ _01490_ _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__07524__I _02032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06571__A3 _02068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07725_ _02077_ _03057_ _03058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__06859__A1 _00621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07656_ _02997_ _03002_ _03013_ _00161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_74_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_74_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06607_ _02103_ _02104_ _02101_ _02105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_07587_ _01165_ _02915_ _02968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_75_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09326_ _02615_ _04239_ _04367_ _04368_ _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_47_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05979__I _01331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06538_ _02035_ _02036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10537__D _00475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09257_ _02384_ _01034_ _04301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06469_ net5 _01390_ _01110_ _01967_ _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_90_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08208_ cpu.uart.data_buff\[2\] _03464_ _03465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09188_ cpu.Z _00709_ _04234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08139_ _03400_ _03409_ _00248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07036__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05598__A1 _01054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07587__A2 _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10101_ _00044_ clknet_leaf_31_wb_clk_i cpu.uart.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output66_I net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10032_ _01991_ _02005_ _04995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_4_0_wb_clk_i clknet_0_wb_clk_i clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_39_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07275__A1 cpu.timer_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_15_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_113_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05428__I2 cpu.regs\[10\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05589__A1 _01090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06250__A2 _00973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05840_ _00816_ _01345_ _01346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__07750__A2 _03080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05771_ _01270_ _01276_ _01277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07510_ cpu.regs\[12\]\[1\] _02919_ _02922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08490_ _03676_ _00332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07441_ _02869_ _02873_ _02823_ _02874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_54_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07502__A2 _01135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07372_ _02802_ _02810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_84_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09111_ _04150_ _04164_ _04165_ _00464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06323_ cpu.pwm_top\[5\] _01178_ _01824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09042_ cpu.regs\[2\]\[6\] _02586_ _04102_ _04113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06254_ _01675_ _01755_ _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05205_ _00740_ _00741_ _00701_ _00728_ _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_53_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06185_ _01594_ _01687_ _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_25_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05136_ _00674_ _00675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08766__A1 _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_121_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_121_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_96_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09944_ _04713_ _04913_ _00549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05067_ cpu.regs\[12\]\[5\] cpu.regs\[13\]\[5\] cpu.regs\[14\]\[5\] cpu.regs\[15\]\[5\]
+ _00572_ _00576_ _00609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_0_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09875_ _04837_ _04854_ _04862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08826_ cpu.timer_capture\[12\] _03941_ _03943_ _03939_ _03944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__09191__A1 _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_93_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08757_ cpu.timer\[8\] _03879_ _03886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05969_ _01462_ _01464_ _01466_ _01440_ _01473_ _01474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08688_ _02658_ _03824_ _03828_ _03827_ _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09494__A2 _04028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07708_ _01700_ _03040_ _03045_ _00181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07639_ _02980_ _03001_ _03003_ _00154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09309_ _04351_ _04352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10581_ _00519_ clknet_leaf_70_wb_clk_i net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_90_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05363__S0 _00872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07009__A1 cpu.ROM_addr_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05658__B _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10015_ _04214_ _04215_ _04216_ _04978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05743__A1 cpu.timer_top\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_4_Left_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08996__A1 _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07990_ cpu.uart.receive_counter\[0\] cpu.uart.receive_counter\[1\] cpu.uart.receive_counter\[3\]
+ cpu.uart.receive_counter\[2\] _03284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_06941_ _02404_ _02407_ _02437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09660_ _02484_ _02537_ _04641_ _04690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__09173__B2 _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08611_ _03738_ _03774_ _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06872_ _02367_ _02369_ _02370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_82_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09591_ _00772_ _04621_ _04624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05823_ _01311_ _01322_ _01328_ _01329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_89_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08542_ _03652_ cpu.toggle_ctr\[0\] _03728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05754_ _01170_ _01173_ _01251_ _01256_ _01259_ _01260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_85_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08473_ _02758_ _03655_ _03664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07424_ cpu.uart.divisor\[10\] _02857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_92_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05685_ _01097_ _01191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_59_Left_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07239__A1 _00989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07355_ _02384_ _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06306_ net44 _01616_ _01805_ _01806_ _01514_ _01807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_93_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07286_ cpu.timer_top\[5\] _02740_ _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08987__B2 _01018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09025_ _04100_ _00443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06237_ _00597_ _01739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_60_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06168_ _01670_ _01671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06214__A2 _01390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Left_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06099_ _01602_ _01603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05119_ _00656_ _00657_ _00658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_09927_ _02652_ _04900_ _04901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09858_ net81 _04841_ _04849_ _04847_ _04850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08911__A1 _02853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09789_ net73 _04793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08809_ _03921_ _03930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_68_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08808__I _03918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_77_Left_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09219__A2 _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10564_ _00502_ clknet_leaf_76_wb_clk_i cpu.ROM_spi_dat_out\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07159__I _02635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10495_ _00433_ clknet_leaf_55_wb_clk_i cpu.IO_addr_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06012__B _01053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05407__I _00918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07705__A2 _03041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput9 io_in[17] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05716__B2 _01221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09170__A4 _02418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09458__A2 _01036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07622__I _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05470_ cpu.regs\[8\]\[4\] cpu.regs\[9\]\[4\] cpu.regs\[10\]\[4\] cpu.regs\[11\]\[4\]
+ _00871_ _00977_ _00979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_117_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07140_ _02620_ _02621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07071_ _02037_ _02340_ _02557_ _02558_ _02559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_23_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06022_ cpu.spi.divisor\[2\] _01191_ _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08197__A2 _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09712_ _04731_ _04732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07973_ cpu.spi.data_in_buff\[1\] _03270_ _03272_ cpu.spi.data_in_buff\[0\] _03274_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09146__A1 _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06924_ _02414_ _02420_ _02421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05317__I _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05707__A1 net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09643_ cpu.ROM_addr_buff\[6\] _04666_ _04673_ _04674_ _04675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_87_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06855_ _02098_ _02113_ _02353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09574_ _00769_ _04314_ _04607_ _04321_ _04608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05806_ _00715_ _01312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08525_ _03699_ cpu.toggle_top\[6\] cpu.toggle_top\[5\] _03701_ _03710_ _03711_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06786_ _02260_ _02283_ _02284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05737_ _01068_ _01058_ _01243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_38_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08456_ _03354_ _03574_ _00323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05668_ _01104_ _01111_ _01174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07407_ cpu.uart.divisor\[15\] _02840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_08387_ cpu.orig_IO_addr_buff\[7\] _03596_ _03602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05599_ _01068_ _01050_ _01105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07338_ _02613_ _02778_ _02616_ _02779_ _00077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__05987__I _01379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07269_ _02728_ _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10280_ _00219_ clknet_leaf_47_wb_clk_i cpu.spi.data_in_buff\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09008_ _02524_ _04085_ _04088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06294__S1 _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06611__I _02108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_85_Left_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08360__A2 _03581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06371__A1 net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10616_ _00554_ clknet_leaf_72_wb_clk_i net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_94_Left_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_107_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10547_ _00485_ clknet_leaf_84_wb_clk_i cpu.PC\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10478_ _00417_ clknet_leaf_21_wb_clk_i cpu.timer_div\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06640_ _00822_ _01995_ _02138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05165__A2 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06571_ _02037_ _02064_ _02068_ _02069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_08310_ _02868_ _03541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05522_ _00651_ _01027_ _01028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09290_ _04253_ _04334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08241_ cpu.uart.data_buff\[8\] _03459_ _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05453_ _00901_ _00963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08172_ cpu.uart.div_counter\[15\] _03432_ _03435_ _03436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_103_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05384_ _00868_ _00895_ _00896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07123_ _02524_ _02607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_112_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07054_ _02534_ _02077_ _02540_ _02542_ _02543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
Xclkbuf_leaf_99_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_99_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_28_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_28_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06005_ _01043_ _01047_ _01122_ _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__07917__A2 cpu.spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05928__A1 _01429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07956_ _02657_ _03241_ _03260_ _03261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08590__A2 _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input28_I sram_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06907_ _02075_ _02404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_106_Right_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07887_ _03202_ _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_69_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09626_ cpu.last_addr\[12\] cpu.ROM_addr_buff\[12\] _04657_ _04658_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_69_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06838_ _02331_ _02323_ _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05400__I0 cpu.regs\[12\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_qcpu_109 io_out[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09557_ _04514_ _04571_ _04592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06769_ _02263_ _02265_ _02267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08508_ cpu.toggle_ctr\[15\] _03693_ _03690_ cpu.toggle_ctr\[14\] _03694_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_38_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09488_ _04499_ _04525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08439_ _03638_ _03639_ _03630_ _00318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_65_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05510__I _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10401_ _00340_ clknet_leaf_7_wb_clk_i cpu.toggle_ctr\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10332_ _00271_ clknet_leaf_43_wb_clk_i cpu.uart.receiving vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output96_I net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10263_ _00202_ clknet_leaf_33_wb_clk_i cpu.spi.div_counter\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10194_ _00133_ clknet_leaf_1_wb_clk_i cpu.regs\[0\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09652__I _04683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07844__B2 _01802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07844__A1 _01879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput12 io_in[1] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_114_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput23 io_in[8] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_12_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07775__C _02628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05473__I3 cpu.regs\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07810_ cpu.timer_div\[5\] _03126_ cpu.timer_div_counter\[7\] _01976_ _03130_ _03131_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08790_ _03908_ _03837_ _03909_ _03913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_4_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06583__A1 _00972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07741_ _03063_ _03072_ _03073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07672_ _03023_ _00167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07082__I _02569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09411_ cpu.orig_PC\[6\] _04043_ _04451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06623_ _02103_ _02104_ _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06554_ cpu.mem_cycle\[5\] _02052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09342_ _04383_ _04384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05505_ _01011_ _01012_ _00885_ _01013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06485_ cpu.toggle_top\[15\] _01263_ _01958_ _01984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09273_ _04027_ _04317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08224_ _00975_ _03476_ _03477_ _03478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05436_ _00946_ _00947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__05330__I _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08155_ _03324_ _03421_ _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_95_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09588__A1 cpu.PC\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05367_ _00873_ _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_113_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07106_ _01370_ _01989_ _02028_ _02030_ _02542_ _02592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08086_ cpu.uart.div_counter\[0\] _03365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05298_ _00003_ _00827_ _00829_ _00830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_100_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07037_ _02515_ _02527_ _02528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08988_ _00749_ _04029_ _04040_ _04071_ _04059_ _04072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__06574__A1 _02071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07939_ cpu.spi.data_out_buff\[1\] _03234_ _03245_ _03247_ _03248_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06326__A1 cpu.toggle_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09609_ _02510_ _03995_ _00736_ _04641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08079__A1 _03354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06764__C _02261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10315_ _00254_ clknet_leaf_32_wb_clk_i cpu.uart.div_counter\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05455__I3 cpu.regs\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10246_ _00185_ clknet_leaf_109_wb_clk_i cpu.regs\[3\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06014__B1 _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10177_ _00116_ clknet_leaf_126_wb_clk_i cpu.regs\[11\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06317__A1 cpu.timer_div\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09503__A1 _00823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_44_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06270_ _01770_ _01751_ _01771_ _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05150__I _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05221_ cpu.br_rel_dest\[5\] _00756_ _00757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_8_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08242__A1 _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05152_ _00689_ _00690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08461__I _03653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09960_ cpu.ROM_addr_buff\[0\] _04927_ _02501_ cpu.ROM_addr_buff\[4\] cpu.ROM_addr_buff\[8\]
+ _02502_ _04928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_TAPCELL_ROW_77_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05083_ _00619_ _00622_ _00623_ _00624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08911_ _02853_ _04001_ _04005_ _04006_ _04007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_90_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09042__I0 cpu.regs\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09891_ _04010_ _04866_ _04874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_83_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08842_ cpu.timer_capture\[15\] _03941_ _03955_ _03956_ _03957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08773_ cpu.timer\[12\] _03894_ _03890_ _03899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_05985_ net27 _01309_ _01490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07724_ _02378_ _02585_ _03057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_79_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07655_ cpu.regs\[6\]\[7\] _03000_ _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_40_Left_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06606_ _00850_ _01955_ _02104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07540__I _01788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07586_ _02033_ _02967_ _00137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07108__I0 _02418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07808__A1 cpu.timer_div\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07808__B2 cpu.timer_div\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09325_ _00775_ _04368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06537_ _00708_ _01270_ _01039_ _02035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_06468_ _01218_ _01965_ _01966_ _01967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_62_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08481__A1 _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09256_ cpu.PC\[1\] cpu.br_rel_dest\[1\] _04300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_43_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_43_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08207_ _03450_ _03464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05419_ _00929_ _00930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_16_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05295__A1 _00002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06399_ _01879_ _01639_ _01897_ _01898_ _01413_ _01899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_50_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09467__I _04313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09187_ _04232_ _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08138_ _03407_ _03403_ _03408_ _03401_ _03409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07036__A2 _02516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08069_ _03221_ cpu.spi.counter\[1\] _03352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10100_ _00043_ clknet_leaf_31_wb_clk_i cpu.uart.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06795__A1 _00801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10031_ _01992_ _04993_ _04994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output59_I net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08224__A1 _00975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09972__A1 _04114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10031__A1 _01992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05428__I3 cpu.regs\[11\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10229_ _00168_ clknet_leaf_115_wb_clk_i cpu.regs\[5\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05770_ _01275_ _01276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05145__I _00683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_0_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07440_ _02872_ _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07371_ _02809_ _00080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09110_ cpu.last_addr\[8\] _04157_ _04165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06322_ cpu.timer_top\[13\] _01413_ _01124_ _01822_ _01823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_44_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09041_ _04112_ _00447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06253_ _01744_ _01753_ _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05204_ _00653_ _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06184_ _01551_ _00956_ _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_25_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05135_ cpu.instr_cycle\[2\] _00651_ _00661_ _00673_ _00674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_52_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10022__A1 _01299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09943_ cpu.ROM_spi_mode _04912_ _04913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05066_ _00602_ _00607_ _00583_ _00608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09874_ _04861_ _00531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08518__A2 _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06529__A1 _01031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08825_ _03141_ _03928_ _03929_ _03942_ _03943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA_input10_I io_in[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08756_ cpu.timer\[9\] _03885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05968_ _01467_ _01450_ _01472_ _01473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_95_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05899_ _01403_ _01383_ _01404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_68_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08687_ cpu.timer_top\[13\] _03825_ _03828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07707_ cpu.regs\[3\]\[3\] _03039_ _03045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07638_ cpu.regs\[6\]\[0\] _03002_ _03003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05060__S0 _00600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07569_ cpu.regs\[10\]\[7\] _02949_ _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09308_ _04349_ _04350_ _04351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10580_ _00518_ clknet_leaf_68_wb_clk_i net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_106_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09239_ _00751_ _00761_ _04280_ _04283_ _04284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__05363__S1 _00874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10013__A1 _00655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10014_ _04211_ _04977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_116_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_63_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07180__I _02652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08445__A1 _03090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_75_Right_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10193__D _00132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_105_Left_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06940_ _02429_ _02435_ _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input2_I io_in[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09173__A2 _04209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06871_ _02081_ _02136_ _02368_ _02369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08610_ cpu.pwm_counter\[6\] _03772_ _03774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05822_ _01326_ _01327_ _01328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_84_Right_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09590_ _00778_ _00773_ _04623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06931__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08541_ _03726_ _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05753_ _01258_ _01259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05684_ cpu.spi.divisor\[0\] _01190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_85_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08684__A1 cpu.timer_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08472_ _03663_ _00327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07487__A2 _02905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05603__I _01108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07423_ cpu.uart.divisor\[13\] _02856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_106_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_114_Left_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07354_ _02406_ _02791_ _02793_ _02558_ _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06305_ net56 _01615_ _01509_ _01806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07285_ _02653_ _02739_ _02741_ _02737_ _00062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_45_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_93_Right_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09024_ _04099_ cpu.ROM_addr_buff\[1\] _03998_ _04100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06236_ _01704_ _01302_ _01736_ _01737_ _01738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_14_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06167_ _01658_ _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06098_ _01601_ _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05118_ cpu.base_address\[1\] cpu.base_address\[0\] _00657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_09926_ _04887_ _04900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05049_ cpu.regs\[0\]\[4\] _00590_ _00591_ cpu.regs\[3\]\[4\] _00571_ _00575_ _00592_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__05273__I1 _00801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05422__A1 _00896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07265__I _02635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09164__A2 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09857_ _04823_ _04842_ _04849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07175__A1 _02648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09788_ _03227_ _04792_ _00514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08808_ _03918_ _03929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06922__A1 _02418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08739_ cpu.timer\[6\] cpu.timer\[5\] _03860_ _03871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_68_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08675__A1 _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05513__I _00868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06150__A2 _01652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08427__A1 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10563_ _00501_ clknet_leaf_74_wb_clk_i cpu.ROM_spi_dat_out\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09927__A1 _02652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10494_ _00432_ clknet_leaf_55_wb_clk_i cpu.IO_addr_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08418__A1 _03623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09091__A1 cpu.ROM_addr_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07070_ net12 _02405_ _02551_ _02558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06021_ _01096_ _01076_ _01500_ _01524_ _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__05652__A1 _00720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09394__A2 _00706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09711_ _02505_ _04731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07972_ _03097_ _03270_ _03272_ _03273_ _00217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06923_ _02091_ _02415_ _02417_ _02419_ _02420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_87_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09642_ cpu.last_addr\[4\] cpu.ROM_addr_buff\[4\] _04648_ _04674_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06854_ _02203_ _02350_ _02351_ _02352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09573_ _04505_ _04606_ _04607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06785_ _02272_ _02281_ _02282_ _02283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05805_ _01310_ _01311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05736_ _01241_ _01242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08524_ _03705_ _03708_ _03709_ _03710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05333__I cpu.PORTA_DDR\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08455_ _03650_ _03651_ _03646_ _00322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05667_ _01172_ _01173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07406_ cpu.uart.receive_div_counter\[4\] cpu.uart.divisor\[4\] _02839_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05598_ _01054_ _01103_ _01104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08386_ cpu.IO_addr_buff\[7\] _03598_ _03601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_21_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09082__A1 _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07337_ _02610_ _02778_ _02612_ _02779_ _00076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_9_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07268_ _02728_ _02729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07632__A2 _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06219_ cpu.uart.dout\[4\] _01195_ _01718_ _01720_ _01102_ _01721_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__09909__A1 _01059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07199_ _02668_ _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09007_ _04087_ _00438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09909_ _01059_ _04812_ _04887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08896__A1 _00700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output41_I net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05243__I _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07320__A1 cpu.toggle_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10615_ _00553_ clknet_leaf_74_wb_clk_i net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_3_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05309__S1 _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10546_ _00484_ clknet_leaf_84_wb_clk_i cpu.PC\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07623__A2 _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10477_ _00416_ clknet_leaf_21_wb_clk_i cpu.timer_div\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09376__A2 _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06570_ _02066_ _02067_ _02068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07789__B _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_82_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05521_ _01025_ _01026_ _01027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08240_ cpu.uart.data_buff\[9\] _03451_ _03489_ _03490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05452_ _00961_ _00962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_117_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08171_ cpu.uart.div_counter\[15\] _03404_ _03430_ _03435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_6_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07301__C _02712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05383_ _00894_ _00895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07122_ _02595_ _02603_ _02604_ _02606_ _00034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_103_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07614__A2 _02986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07053_ _02541_ _02542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_113_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06004_ net81 _00675_ _01069_ _01243_ _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_23_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_68_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_68_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07955_ cpu.spi.data_out_buff\[4\] _03231_ _03260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08878__A1 _02758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06906_ _01874_ _02401_ _02402_ _00606_ _02403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_09625_ cpu.last_addr\[11\] _04653_ _04657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07886_ _03203_ _03204_ _03205_ _00199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_54_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06837_ _02325_ _02334_ _02335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_78_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09556_ _04488_ _04571_ _04590_ _04511_ _04591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06768_ _00927_ _02263_ _02265_ _02266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_05719_ cpu.uart.dout\[0\] _00012_ _01225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09487_ _04523_ _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08507_ cpu.toggle_top\[15\] _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_38_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06699_ _02193_ _02195_ _02196_ _02197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__05998__I _01197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08438_ cpu.orig_PC\[9\] _03628_ _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08369_ cpu.orig_IO_addr_buff\[3\] _03587_ _03588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08802__A1 _02635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10400_ _00339_ clknet_leaf_7_wb_clk_i cpu.toggle_ctr\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10331_ _00270_ clknet_leaf_58_wb_clk_i cpu.uart.data_buff\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output89_I net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10262_ _00201_ clknet_leaf_33_wb_clk_i cpu.spi.div_counter\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07369__A1 _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10193_ _00132_ clknet_leaf_107_wb_clk_i cpu.regs\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06041__A1 _00920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08869__A1 cpu.timer_div\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_34_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05701__I _01200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05855__A1 _00992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput13 io_in[20] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput24 io_in[9] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_52_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10529_ _00467_ clknet_leaf_78_wb_clk_i cpu.last_addr\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05148__I _00685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_73_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07080__I0 _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07740_ _01493_ _02073_ _03070_ _03071_ _03052_ _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__06335__A2 _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07671_ _03009_ cpu.regs\[5\]\[5\] _03014_ _03023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07532__A1 cpu.regs\[11\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09410_ _04312_ _04449_ _04450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06622_ _02117_ _02118_ _02119_ _02120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06553_ _02050_ _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_90_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09341_ _02381_ _04349_ _04383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_114_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05504_ cpu.regs\[0\]\[5\] cpu.regs\[1\]\[5\] cpu.regs\[2\]\[5\] cpu.regs\[3\]\[5\]
+ _00871_ _00900_ _01012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_118_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06484_ cpu.toggle_top\[7\] _01255_ _01982_ _01258_ _01983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_09272_ _04315_ _04316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_115_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_115_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08223_ cpu.uart.data_buff\[5\] _03464_ _03477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05435_ _00945_ _00946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08154_ cpu.uart.div_counter\[11\] _03415_ _03421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08922__I _04000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05366_ _00877_ _00878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08085_ _03360_ _03363_ _03364_ _00238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07105_ _02407_ _02584_ _02590_ _02591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07036_ net19 _02516_ _02527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05297_ _00579_ _00828_ _00829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08987_ cpu.orig_IO_addr_buff\[5\] _04056_ _04057_ _01018_ _04071_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07938_ _03246_ _03247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_98_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07869_ cpu.spi.div_counter\[3\] _03187_ _03188_ cpu.spi.divisor\[4\] _03189_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__06326__A2 _01106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09608_ _02466_ _04640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_104_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09539_ _04446_ _04573_ _04574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_118_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09579__A2 _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06262__A1 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07054__A3 _02540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10314_ _00253_ clknet_leaf_38_wb_clk_i cpu.uart.div_counter\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10245_ _00184_ clknet_leaf_114_wb_clk_i cpu.regs\[3\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06014__A1 _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10176_ _00115_ clknet_leaf_3_wb_clk_i cpu.regs\[11\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06565__A2 _01156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07762__A1 _02076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05391__I3 cpu.regs\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05828__A1 _01332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05220_ cpu.br_rel_dest\[4\] _00756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05151_ _00688_ _00689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_8_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05082_ _00583_ _00623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09890_ _04873_ _00535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_100_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08910_ _03987_ _04006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_90_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09042__I1 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08841_ _03794_ _03956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09506__C _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07753__A1 _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08772_ _03896_ _03898_ _00392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05984_ _01448_ _01475_ _01488_ net91 _01366_ _01489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_07723_ _02570_ _02346_ _03055_ _03056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07654_ _03012_ _00160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06605_ _02101_ _02102_ _02103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07585_ _01910_ _01948_ _02967_ _00136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09324_ _04239_ _04366_ _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06536_ _01375_ _02033_ _02034_ _00020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06467_ net67 _01515_ _01966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09255_ _04298_ _04299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_8_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08206_ _03461_ _03463_ _00261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05418_ _00928_ _00929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06398_ cpu.timer_capture\[14\] _01233_ _01247_ _01898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09186_ _00710_ _00774_ _04232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08137_ _03407_ _03404_ _03408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05349_ _00861_ net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08068_ cpu.spi.counter\[1\] _03349_ _03351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_83_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_83_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06172__I _01471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07019_ _00697_ _02060_ _02061_ _02512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_12_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_12_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09483__I _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10030_ _01990_ _02002_ _04993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_110_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05516__I _01022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05251__I _00685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07178__I _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06235__A1 _00974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09024__I1 cpu.ROM_addr_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09607__B _00690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10228_ _00167_ clknet_leaf_114_wb_clk_i cpu.regs\[5\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10159_ _00098_ clknet_leaf_2_wb_clk_i cpu.regs\[13\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07370_ _02808_ _02078_ _02789_ _02809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07797__B _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06321_ _01802_ _01247_ _01820_ _01821_ _01413_ _01822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09040_ _04111_ cpu.ROM_addr_buff\[5\] _04104_ _04112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06252_ _01745_ _01753_ _01754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05203_ _00739_ _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06183_ _01674_ _01679_ _01685_ _01686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05134_ _00672_ _00673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06226__A1 _01708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09942_ _02463_ _02042_ _04910_ _04911_ _04912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_96_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05065_ cpu.regs\[0\]\[5\] _00605_ _00606_ cpu.regs\[3\]\[5\] _00600_ _00601_ _00607_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_110_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09873_ net57 _04853_ _04860_ _04858_ _04861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06529__A2 _02027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08824_ _00989_ _03930_ _03942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08755_ _03882_ _03884_ _00389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05967_ _01468_ _01471_ _01472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07706_ _01602_ _03040_ _03044_ _00180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05898_ cpu.spi.dout\[1\] _01403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_68_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08686_ _02653_ _03824_ _03826_ _03827_ _00377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_95_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07637_ _02999_ _03002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05060__S1 _00601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07568_ _02958_ _00128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09307_ _03623_ _04348_ _04350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06519_ _01451_ _01999_ _02017_ _01461_ _02018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_118_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06465__A1 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07499_ cpu.regs\[13\]\[7\] _02903_ _02913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09238_ cpu.orig_PC\[1\] _04281_ _04282_ _00761_ _04283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_35_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09169_ _02611_ _02261_ _02109_ _02614_ _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_4_8_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output71_I net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09167__B1 _02261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10013_ _00655_ _01453_ _04340_ _04976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08390__A1 _01311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08557__I _02521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07956__A1 _02657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07708__A1 _01700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05431__A2 _00941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06870_ _02114_ _02135_ _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_66_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05821_ _01310_ _01322_ _01327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08540_ _03725_ _03726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05752_ _01257_ _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05683_ _01188_ _01189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08471_ cpu.toggle_top\[2\] _03654_ _03662_ _03660_ _03663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_49_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10011__B net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09881__A1 _04815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07422_ _02851_ _02852_ _02854_ _02855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_85_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07353_ _02792_ _01022_ _01540_ _02327_ _02793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06304_ cpu.PORTA_DDR\[5\] _01613_ _01805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_73_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07284_ cpu.timer_top\[4\] _02740_ _02741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09023_ _00823_ _02797_ _00732_ _04099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06235_ _00974_ _01285_ _01302_ _01301_ _01737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_103_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07947__B2 _03247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06166_ _01655_ _01668_ _01669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06097_ _01497_ _01547_ _01600_ _01492_ _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_05117_ cpu.base_address\[3\] cpu.base_address\[2\] _00656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_09925_ _04887_ _04899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05048_ cpu.regs\[2\]\[4\] _00591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__05273__I2 _00802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09856_ _04848_ _00526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08807_ _03921_ _03928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09787_ net74 _03724_ _04792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06999_ _02491_ _02492_ _02493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_99_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06922__A2 _01957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08738_ _03868_ _03870_ _00386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08669_ _03802_ _03815_ _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09872__A1 _04022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10562_ _00500_ clknet_leaf_73_wb_clk_i cpu.spi_clkdiv vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06438__B2 _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06438__A1 _01484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10493_ _00431_ clknet_leaf_17_wb_clk_i cpu.IO_addr_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06429__A1 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06020_ _01501_ _01523_ _01193_ _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07567__S _02948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05652__A2 _01156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07971_ net16 _03273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09710_ _04728_ _04730_ _00498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06922_ _02418_ _01957_ _02091_ _02419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09641_ _04668_ _04670_ _04671_ _04672_ _04673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_87_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05168__A1 _00690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06853_ _02137_ _02165_ _02351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_117_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09572_ _02375_ _00772_ _04605_ _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06784_ _02279_ _02280_ _02282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05804_ cpu.C _01310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_05735_ _01240_ _01241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08523_ _03701_ cpu.toggle_top\[5\] cpu.toggle_top\[4\] _03706_ _03709_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_93_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07034__C _02522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08454_ cpu.orig_PC\[13\] _03642_ _03651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05666_ _01171_ _01172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07405_ cpu.uart.divisor\[11\] cpu.uart.receive_div_counter\[11\] _02838_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05597_ _01056_ _01055_ _01103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08385_ _03599_ _03600_ _03570_ _00303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07336_ _02607_ _02778_ _02609_ _02779_ _00075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_21_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07267_ _01243_ _02727_ _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09006_ _01020_ _04084_ _04086_ _04020_ _04087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_103_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06218_ _01522_ _01719_ _01720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07198_ _01295_ _02668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06149_ _01607_ _01301_ _01650_ _01651_ _01652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_13_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09908_ _04886_ _00540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09839_ _04022_ _04829_ _04835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_29_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_24_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05706__I0 cpu.PORTA_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10614_ _00552_ clknet_leaf_74_wb_clk_i net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10545_ _00483_ clknet_leaf_97_wb_clk_i cpu.PC\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10476_ _00415_ clknet_leaf_21_wb_clk_i cpu.timer_div\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07186__I _02657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_63_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_69_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05434__I _00944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05520_ cpu.instr_cycle\[2\] cpu.instr_cycle\[3\] cpu.instr_cycle\[1\] _00673_ _01026_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_05451_ _00898_ _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_27_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08170_ _03433_ _03434_ _03381_ _00254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07862__A3 _00765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07121_ _02605_ _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05382_ _00893_ _00894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_27_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07052_ _01137_ _02067_ _02541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_30_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06003_ _01196_ _01048_ _01063_ cpu.PORTA_DDR\[2\] _01507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_51_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05609__I _00675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07954_ _03259_ _00213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07885_ cpu.spi.div_counter\[0\] _03184_ _03205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06905_ _02069_ _02402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09624_ cpu.ROM_addr_buff\[13\] _04655_ _04656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06836_ _02168_ _02333_ _02329_ _02334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_37_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05344__I cpu.PORTA_DDR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_37_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_37_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09827__A1 _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09555_ _04587_ _04589_ _04590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06767_ _00876_ _00881_ _00884_ _00891_ _02264_ _02265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_05718_ _01198_ _01222_ _01223_ _01224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08506_ cpu.toggle_ctr\[14\] _03690_ _03691_ _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09486_ _03076_ _04489_ _04522_ _04523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06698_ _02191_ _02192_ _02196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07689__I0 _03007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_108_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08437_ _03637_ _03633_ _03638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05649_ _01154_ _01155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__05313__A1 _00566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08368_ _03586_ _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08299_ cpu.uart.receive_div_counter\[5\] _03525_ _03532_ _03533_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07319_ _02766_ _02763_ _02767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10330_ _00269_ clknet_leaf_54_wb_clk_i cpu.uart.data_buff\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10261_ _00200_ clknet_leaf_33_wb_clk_i cpu.spi.div_counter\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10192_ _00131_ clknet_leaf_11_wb_clk_i cpu.regs\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_6_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05254__I _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09597__S _04440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput14 io_in[21] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput25 rst_n net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_10528_ _00466_ clknet_leaf_81_wb_clk_i cpu.last_addr\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_12_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10459_ _00398_ clknet_leaf_7_wb_clk_i cpu.timer_capture\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_20_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06688__C _02185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07670_ _03022_ _00166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06621_ _02115_ _02116_ _02119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06552_ cpu.mem_cycle\[0\] _02050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09340_ _02561_ _04344_ _04382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09271_ _01149_ _04315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05503_ cpu.regs\[4\]\[5\] cpu.regs\[5\]\[5\] cpu.regs\[6\]\[5\] cpu.regs\[7\]\[5\]
+ _00887_ _00900_ _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_114_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08222_ _03454_ _03476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06483_ _01959_ _01253_ _01981_ _01172_ _01982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_74_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05434_ _00944_ _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_31_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08153_ _03400_ _03420_ _00251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05365_ _00004_ _00877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_99_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08084_ _03238_ _03200_ _03364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08796__A1 _01074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07104_ _02585_ _02589_ _02407_ _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07035_ _02526_ _00027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05296_ cpu.regs\[8\]\[1\] cpu.regs\[9\]\[1\] cpu.regs\[10\]\[1\] cpu.regs\[11\]\[1\]
+ _00568_ _00804_ _00828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_113_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05339__I cpu.PORTA_DDR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07220__A1 cpu.timer_capture\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08986_ _04055_ _04070_ _00434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input33_I sram_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07937_ _02660_ _03246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07554__I _02948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07868_ cpu.spi.div_counter\[4\] _03188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_39_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07799_ _02735_ _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09607_ _04619_ _04639_ _00690_ _00486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06819_ _02316_ _02305_ _02317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09538_ _04315_ _04570_ _04572_ _04573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07287__A1 _02658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09469_ _04364_ _04491_ _04506_ _04313_ _04507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_109_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10313_ _00252_ clknet_leaf_31_wb_clk_i cpu.uart.div_counter\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_115_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08539__A1 _03232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10244_ _00183_ clknet_leaf_113_wb_clk_i cpu.regs\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__06014__A2 _01053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07211__A1 _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10175_ _00114_ clknet_leaf_126_wb_clk_i cpu.regs\[11\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07762__A2 _02391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09019__A2 _00802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05150_ _00687_ _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_100_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05159__I _00696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05081_ cpu.regs\[0\]\[6\] _00621_ cpu.regs\[2\]\[6\] cpu.regs\[3\]\[6\] _00617_
+ _00618_ _00622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_21_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08840_ _03920_ _03954_ _03955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08771_ cpu.timer_capture\[11\] _03883_ _03897_ _03898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05983_ _01478_ _01482_ _01487_ _01488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07722_ _02284_ _02344_ _02345_ _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__08702__A1 _01059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07653_ _03011_ cpu.regs\[6\]\[6\] _02999_ _03012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_88_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06604_ _02099_ _02100_ _02102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09323_ _02811_ _04364_ _04365_ _04366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07584_ _01833_ _01872_ _02967_ _00135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_34_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06535_ cpu.regs\[9\]\[7\] _01702_ _02034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06466_ cpu.PORTB_DDR\[7\] _01385_ _01964_ _01215_ _01965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_63_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09254_ _04278_ _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08205_ _03462_ cpu.uart.data_buff\[1\] _03451_ _03463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09185_ _03604_ _04195_ _04230_ _04231_ _00472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05417_ _00927_ _00928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08136_ cpu.uart.div_counter\[8\] _03407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06397_ cpu.timer_capture\[6\] _01181_ _01894_ _01896_ _01241_ _01897_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_05348_ net75 cpu.ROM_spi_mode _00861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07441__A1 _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08067_ _03347_ _03239_ _03350_ _00234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05279_ _00580_ _00811_ _00812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07018_ _00736_ _02510_ _02511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_101_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_52_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_52_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08969_ _04043_ _04056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09004__I _04083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07432__A1 _00787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05294__I0 cpu.regs\[12\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10227_ _00166_ clknet_leaf_116_wb_clk_i cpu.regs\[5\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08932__A1 _04022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07194__I _02664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10158_ _00097_ clknet_leaf_1_wb_clk_i cpu.regs\[14\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10089_ _00032_ clknet_leaf_112_wb_clk_i cpu.regs\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06171__A1 _01452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06171__B2 _01466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06320_ cpu.timer_capture\[13\] _01232_ _01247_ _01821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08753__I _03835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06251_ _01678_ _01752_ _01753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05202_ _00738_ _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06182_ _01152_ _01660_ _01684_ _01462_ _01685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_25_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05133_ net71 _00665_ _00668_ _00671_ _00672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_09941_ _02449_ _04704_ _04911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05064_ cpu.regs\[2\]\[5\] _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09517__C _00776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05985__A1 net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09872_ _04022_ _04854_ _04860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08923__A1 _04014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08823_ _03918_ _03941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08754_ cpu.timer_capture\[8\] _03883_ _03869_ _03884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05966_ _01470_ _01471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07705_ cpu.regs\[3\]\[2\] _03041_ _03044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05897_ _01401_ cpu.spi.divisor\[1\] _01191_ _01402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08685_ _02736_ _03827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07636_ _03000_ _03001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05352__I _00863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07567_ _02945_ cpu.regs\[10\]\[6\] _02948_ _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09306_ _03623_ _04348_ _04349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_8_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06518_ net97 _02016_ _02017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_118_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09237_ _04281_ _04265_ _04282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07498_ _02912_ _00104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06449_ _01910_ _01948_ _01949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09168_ _01304_ _02185_ _04213_ _02608_ _04215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08119_ cpu.uart.div_counter\[5\] _03393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09099_ _04141_ _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09167__A1 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output64_I net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09167__B2 _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10012_ _04965_ _04972_ _04975_ _03347_ _00555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08914__A1 cpu.uart.divisor\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09642__A2 cpu.ROM_addr_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07189__I _02660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05211__B _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07405__A1 cpu.uart.divisor\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05865__C _01370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09158__B2 _02027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05820_ _01325_ _01326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_19_Left_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05751_ _01117_ _01204_ _01257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_106_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05682_ _01187_ _01188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08470_ _02754_ _03655_ _03662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06144__A1 _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07421_ _02853_ cpu.uart.receive_div_counter\[9\] _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_106_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07352_ _02288_ _02792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06303_ cpu.uart.divisor\[5\] _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_73_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07283_ _02728_ _02740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_28_Left_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09022_ _04098_ _00442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06234_ _01707_ _01282_ _01426_ _01735_ _01736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_3_0_wb_clk_i clknet_0_wb_clk_i clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_06165_ _01437_ _01660_ _01667_ _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05116_ cpu.instr_buff\[15\] _00653_ cpu.base_address\[5\] _00654_ _00655_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_40_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06096_ net28 _01598_ _01599_ _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09924_ _04898_ _00544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05047_ _00589_ _00590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_0_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05273__I3 cpu.regs\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09855_ net80 _04841_ _04845_ _04847_ _04848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08806_ _03927_ _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_37_Left_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09786_ _04784_ _04791_ _00513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06998_ cpu.spi_clkdiv _02046_ _02492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_14_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08737_ cpu.timer_capture\[5\] _03858_ _03869_ _03870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06922__A3 _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05949_ _01151_ _01453_ _01454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08668_ cpu.timer_div_counter\[7\] _03814_ _03815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06135__A1 cpu.timer_capture\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07619_ _01601_ _02990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08599_ cpu.pwm_counter\[3\] _03765_ _03766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_24_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_46_Left_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10561_ _00499_ clknet_leaf_76_wb_clk_i cpu.startup_cycle\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_91_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10492_ _00430_ clknet_leaf_18_wb_clk_i cpu.IO_addr_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09388__A1 _02361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08061__C _00239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_53_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05257__I _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_55_Left_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07673__S _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08363__A2 _03581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_101_Right_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06126__A1 cpu.spi.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_64_Left_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_92_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05876__B _01380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07970_ _03271_ _03272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_73_Left_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06921_ _00638_ _02418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09640_ cpu.last_addr\[2\] cpu.ROM_addr_buff\[2\] _04647_ _04672_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_87_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06852_ _02234_ _02348_ _02349_ _02350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__06365__A1 _01451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_109_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_109_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09571_ _00771_ _04598_ _04605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06783_ net98 _02280_ _02281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05803_ _01157_ _01309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_89_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05734_ _01115_ _01239_ _01240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08522_ _03706_ cpu.toggle_top\[4\] cpu.toggle_top\[3\] _03707_ _03708_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_26_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08453_ _03649_ _03581_ _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07404_ _02832_ cpu.uart.divisor\[7\] _02641_ _02833_ _02836_ _02837_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09530__C _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05665_ _01118_ _01171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05596_ _01101_ _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08384_ cpu.orig_IO_addr_buff\[6\] _03596_ _03600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05630__I _01135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07335_ _02595_ _02778_ _02604_ _02779_ _00074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_98_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07266_ _01103_ _02631_ _02727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_5_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06217_ cpu.uart.divisor\[12\] _01503_ _01719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09005_ _02517_ _04085_ _04086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07197_ _02667_ _00048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06148_ _00957_ _01285_ _01301_ _01651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06079_ _01580_ _01582_ _01583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09907_ cpu.PORTB_DDR\[7\] _04876_ _04885_ _04881_ _04886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07493__S _02903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05077__I _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09838_ _04834_ _00522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_29_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09769_ cpu.ROM_spi_dat_out\[7\] _04751_ _00790_ _04780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_57_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10613_ _00551_ clknet_leaf_73_wb_clk_i net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07608__A1 _01144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10544_ _00482_ clknet_leaf_97_wb_clk_i cpu.PC\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10475_ _00414_ clknet_leaf_30_wb_clk_i cpu.timer_div\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06831__A2 _00929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08033__B2 _02827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08033__A1 cpu.uart.divisor\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_7_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_7_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_9_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06595__A1 _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06898__A2 _02395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07847__A1 _01960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05450_ _00914_ _00960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_90_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05381_ _00892_ _00893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07120_ _00779_ _02605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07051_ _02535_ _02536_ _00693_ _02539_ _02540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XPHY_EDGE_ROW_81_Left_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_70_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06002_ net23 _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_93_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06586__A1 cpu.regs\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07953_ cpu.spi.data_out_buff\[4\] _03255_ _03257_ _03258_ _03259_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07884_ cpu.spi.div_counter\[0\] _03184_ _03204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06904_ _02068_ _02401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_97_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09623_ cpu.last_addr\[13\] _04654_ _04655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06835_ _02326_ _02328_ _02333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05625__I cpu.br_rel_dest\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09554_ _04324_ _04571_ _04588_ _04397_ _04589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06766_ _00588_ _02264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_05717_ cpu.uart.divisor\[8\] _01198_ _01223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07838__A1 cpu.timer_top\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08505_ _03687_ cpu.toggle_top\[13\] _03691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09485_ _03065_ _04489_ _04522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06697_ _02176_ _02194_ _02195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08157__B _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_77_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_77_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_78_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05648_ _01037_ _01154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08436_ _03076_ _03637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_34_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08367_ _03578_ _03586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05360__I _00871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07318_ _02708_ _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05579_ _01053_ _01084_ _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_18_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08298_ _03495_ _03531_ _03532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08671__I _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07066__A2 _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07249_ cpu.timer_capture\[5\] _02701_ _02711_ _02712_ _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_10260_ _00199_ clknet_leaf_35_wb_clk_i cpu.spi.div_counter\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09763__A1 _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10191_ _00130_ clknet_leaf_107_wb_clk_i cpu.regs\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_6_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08846__I _03958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05471__S _00869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07829__A1 _01609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput15 io_in[23] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput26 sram_out[0] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_91_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10527_ _00465_ clknet_leaf_80_wb_clk_i cpu.last_addr\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10061__A1 _01700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10458_ _00397_ clknet_leaf_25_wb_clk_i cpu.timer_capture\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10389_ _00328_ clknet_leaf_11_wb_clk_i cpu.toggle_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06620_ _00835_ _01955_ _02118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07660__I _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06551_ _02048_ _02049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_90_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06482_ cpu.timer_top\[15\] _01414_ _01253_ _01980_ _01981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_09270_ _04313_ _04314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05502_ _01008_ _01009_ _00885_ _01010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08221_ _03459_ _03475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05180__I cpu.base_address\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05433_ _00938_ _00943_ _00944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_90_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08705__B _03646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08152_ cpu.uart.div_counter\[11\] _03370_ _03419_ _03379_ _03420_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_71_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08491__I cpu.toggle_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05364_ _00870_ _00875_ _00876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_113_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08083_ cpu.spi.counter\[4\] _03362_ _03363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07103_ _02586_ _02560_ _02588_ _02589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05295_ _00002_ _00826_ _00827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07034_ _00773_ _02514_ _02525_ _02522_ _02526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_43_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_124_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_124_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08985_ _01056_ _04066_ _04068_ _04069_ _04070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07936_ _00922_ _03242_ _03244_ _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input26_I sram_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07867_ cpu.spi.divisor\[3\] _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07798_ _01961_ _03113_ _03119_ _00197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09606_ _04293_ _04635_ _04638_ _04639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06818_ _02308_ _02312_ _02313_ _02316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_104_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09537_ _03089_ _04027_ _04572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06749_ _02236_ _02237_ _02247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_93_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09468_ _04485_ _04315_ _04506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05090__I _00630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08419_ _02561_ _03619_ _03625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09399_ _04437_ _04438_ _04439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08236__A1 _02664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10312_ _00251_ clknet_leaf_38_wb_clk_i cpu.uart.div_counter\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output94_I net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09736__A1 _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09036__I0 _00591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08539__A2 _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10243_ _00182_ clknet_leaf_109_wb_clk_i cpu.regs\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10174_ _00113_ clknet_leaf_124_wb_clk_i cpu.regs\[12\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05265__I net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05525__A2 _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09975__A1 net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06789__A1 _00820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05080_ _00620_ _00621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06005__A3 _01122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08770_ _03121_ _03897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05982_ _01463_ _01483_ _01486_ _01487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07721_ _03051_ _03054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07652_ _01949_ _03011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06603_ _02099_ _02100_ _02101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07583_ _02545_ _02967_ _00134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_87_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09322_ _04315_ _04351_ _04365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06534_ _02032_ _02033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08466__A1 _03658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06465_ net38 _01211_ _01963_ _01385_ _01964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_75_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09253_ _04296_ _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08204_ _03246_ _03462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08218__A1 _00947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06396_ _01181_ _01895_ _01896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09184_ _02605_ _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_8_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05416_ _00926_ _00927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08135_ _03400_ _03406_ _00247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_105_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05347_ cpu.PORTB_DDR\[2\] net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_90_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08066_ _03221_ _03349_ _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05278_ cpu.regs\[8\]\[0\] cpu.regs\[9\]\[0\] cpu.regs\[10\]\[0\] cpu.regs\[11\]\[0\]
+ _00569_ _00805_ _00811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_31_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09718__A1 _03227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07017_ _00671_ _00795_ _02510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08170__B _03381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08941__A2 _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08968_ _03552_ _04055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07919_ _03182_ _03229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08899_ _02660_ _00737_ _03996_ _03997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
Xclkbuf_leaf_92_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_92_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_94_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_21_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_21_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_78_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08209__A1 _02635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05691__A1 _01196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09709__A1 _03738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09185__A2 _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10226_ _00165_ clknet_leaf_109_wb_clk_i cpu.regs\[5\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10157_ _00096_ clknet_leaf_121_wb_clk_i cpu.regs\[14\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06943__A1 _01950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06943__B2 cpu.regs\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10088_ _00031_ clknet_leaf_111_wb_clk_i cpu.regs\[1\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07499__A2 _02903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06250_ net93 _00973_ _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_79_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05201_ cpu.instr_buff\[15\] _00738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06181_ _01680_ _01683_ _01684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_25_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05132_ _00669_ _00670_ _00671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_52_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09940_ _02448_ _04910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05063_ _00604_ _00605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_115_Right_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09871_ _04859_ _00530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_110_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07187__A1 _02658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08822_ _03940_ _00400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08753_ _03835_ _03883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05965_ _01150_ _01469_ _01470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07704_ _01494_ _03040_ _03043_ _00179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05896_ _01193_ _01399_ _01400_ _01401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08684_ cpu.timer_top\[12\] _03825_ _03826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07635_ _02999_ _03000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08944__I _04032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07566_ _02957_ _00127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09305_ _02383_ _02384_ _02781_ _04348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06517_ _00616_ _00632_ _01762_ _02016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_35_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09236_ _04244_ _04281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07497_ _01951_ cpu.regs\[13\]\[6\] _02902_ _02912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06448_ net32 _01368_ _01379_ _01947_ _01948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_90_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06379_ cpu.timer_top\[6\] _01879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09167_ _02608_ _04213_ _02261_ _02611_ _04214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_08118_ _03391_ _03392_ _00244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09098_ cpu.ROM_addr_buff\[5\] _04145_ _04156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08611__A1 _03738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_43_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08049_ cpu.uart.div_counter\[3\] _03335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_102_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10011_ _04965_ _04974_ net77 _04975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_47_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08678__A1 cpu.timer_top\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06153__A2 _00972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06374__I _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08850__A1 _02732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_82_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05967__A2 _01471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10209_ _00148_ clknet_leaf_108_wb_clk_i cpu.regs\[7\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05275__S0 _00803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05750_ cpu.pwm_top\[0\] _01254_ _01255_ _01256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_89_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05453__I _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05681_ _01096_ _01186_ _01187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_82_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07420_ cpu.uart.divisor\[9\] _02853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_85_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07351_ _02168_ _02329_ _02791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06302_ cpu.spi.dout\[5\] _01803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_85_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07282_ _02728_ _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09021_ _04097_ cpu.ROM_addr_buff\[0\] _03998_ _04098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06233_ _01423_ _01734_ _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06164_ _01554_ _01666_ _01667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05115_ cpu.base_address\[4\] _00654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_41_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06095_ _01157_ _01599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08004__I _02617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09923_ cpu.PORTA_DDR\[3\] _04888_ _04897_ _04893_ _04898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05046_ _00588_ _00589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09854_ _04846_ _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_4_12_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08805_ cpu.timer_capture\[8\] _03919_ _03926_ _03916_ _03927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_09785_ cpu.ROM_spi_cycle\[4\] _04790_ _04791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06997_ _02047_ _00733_ _02491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08736_ _03121_ _03869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05948_ _00991_ _00924_ _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05879_ cpu.PORTA_DDR\[1\] net80 _01211_ _01384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08667_ cpu.timer_div_counter\[6\] _03809_ _03814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_71_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07618_ _02988_ _02985_ _02989_ _00147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08598_ _03573_ _03764_ _03765_ _00351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_49_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07549_ cpu.regs\[11\]\[7\] _02934_ _02947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_101_Left_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10560_ _00498_ clknet_leaf_77_wb_clk_i cpu.startup_cycle\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_24_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10491_ _00429_ clknet_leaf_50_wb_clk_i cpu.uart.divisor\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09219_ _02795_ _03614_ _04264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_80_Right_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06071__A1 _01377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08899__A1 _02660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05474__S _00869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07571__A1 _01084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07323__A1 _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07874__A2 cpu.spi.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09076__A1 cpu.ROM_addr_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09000__A1 _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06920_ _02416_ _01997_ _02417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06851_ _02201_ _02202_ _02349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09570_ _04413_ _04602_ _04603_ _04368_ _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06782_ _02250_ _02251_ _02280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05802_ _01298_ _01303_ _01307_ _01308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05733_ _01081_ _01186_ _01239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08521_ cpu.toggle_ctr\[3\] _03707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08452_ cpu.PC\[13\] _03649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07403_ cpu.uart.receive_div_counter\[1\] _02641_ _02629_ _02835_ _02836_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__07865__A2 cpu.spi.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05664_ cpu.toggle_top\[0\] _01170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__05876__A1 _01377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05595_ _01097_ _01100_ _01101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_08383_ cpu.IO_addr_buff\[6\] _03598_ _03599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07331__C _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08814__A1 _02692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07334_ _02605_ _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07617__A2 _02986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07265_ _02635_ _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06216_ _01710_ _01208_ _01716_ _01717_ _01623_ _01718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_84_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08443__B _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09004_ _04083_ _04085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07196_ cpu.uart.divisor\[6\] _02651_ _02666_ _02662_ _02667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08042__A2 cpu.uart.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06147_ _00988_ _01282_ _01426_ _01649_ _01650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__05358__I _00869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06078_ _01468_ _01581_ _01582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09906_ _04837_ _04877_ _04885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05029_ _00571_ _00572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09837_ net64 _04828_ _04832_ _04833_ _04834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09768_ cpu.ROM_spi_dat_out\[6\] _04732_ _04767_ _04779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_57_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08719_ cpu.timer\[2\] cpu.timer\[1\] cpu.timer\[0\] _03854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09699_ _03227_ _04721_ _00496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08502__B1 cpu.toggle_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10612_ _00550_ clknet_leaf_77_wb_clk_i net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__08805__A1 cpu.timer_capture\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07608__A2 _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05619__A1 _01121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10543_ _00481_ clknet_leaf_97_wb_clk_i cpu.PC\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_118_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10474_ _00413_ clknet_leaf_51_wb_clk_i cpu.timer_div\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_118_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09230__A1 cpu.PC\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06595__A2 _02092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07483__I _02903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09533__A2 _04408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06099__I _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07151__C _02628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05380_ _00876_ _00881_ _00884_ _00891_ _00892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_82_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07050_ _02057_ _02055_ _02538_ _02539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_3_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06283__A1 _01031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07658__I _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06001_ cpu.uart.divisor\[2\] _01208_ _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09221__A1 _00751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06035__A1 _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05469__S0 _00871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08710__C _03795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09806__C _00746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07952_ _03246_ _03258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05906__I cpu.timer_capture\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07883_ _03202_ _03203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09524__A2 _04281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06903_ _02070_ _02399_ _02400_ _00021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09622_ cpu.last_addr\[12\] cpu.last_addr\[11\] _04653_ _04654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06834_ _02323_ _02331_ _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_37_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09553_ cpu.orig_PC\[11\] _04178_ _04588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08504_ cpu.toggle_top\[14\] _03690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06765_ _02262_ _02263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05716_ cpu.uart.divisor\[0\] _01202_ _01209_ _01221_ _01222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09484_ _03637_ _04520_ _04521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06696_ _00605_ _00995_ _02175_ _02194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08435_ _02378_ _03592_ _03636_ _03616_ _00317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_19_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05647_ _01029_ _01149_ _01152_ _01128_ _01153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_08366_ _01049_ _03580_ _03585_ _03583_ _00299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08952__I _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05578_ _01054_ _01083_ _01084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07317_ _02765_ _00070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08297_ _02860_ _03527_ _03531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_61_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06274__A1 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07248_ _02661_ _02712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07179_ _01005_ _02652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09212__A1 _04256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10190_ _00129_ clknet_leaf_125_wb_clk_i cpu.regs\[10\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07774__A1 cpu.spi.dout\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09515__A2 _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06329__A2 _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput16 io_in[26] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput27 sram_out[1] net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10526_ _00464_ clknet_leaf_79_wb_clk_i cpu.last_addr\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06265__A1 _01360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10457_ _00396_ clknet_leaf_24_wb_clk_i cpu.timer\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10388_ _00327_ clknet_leaf_9_wb_clk_i cpu.toggle_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06568__A2 _01135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06550_ cpu.mem_cycle\[1\] _02048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06481_ _01960_ _01248_ _01978_ _01979_ _01640_ _01980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05501_ cpu.regs\[8\]\[5\] cpu.regs\[9\]\[5\] cpu.regs\[10\]\[5\] cpu.regs\[11\]\[5\]
+ _00887_ _00900_ _01009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_114_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09690__A1 _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08220_ _03474_ _00264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05432_ _00940_ _00942_ _00943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08151_ cpu.uart.div_counter\[11\] _03415_ _03419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08245__A2 _03288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05363_ cpu.regs\[0\]\[0\] cpu.regs\[1\]\[0\] cpu.regs\[2\]\[0\] cpu.regs\[3\]\[0\]
+ _00872_ _00874_ _00875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_08082_ _03361_ _03222_ _03357_ _03362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_71_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07102_ _02587_ _02588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05294_ cpu.regs\[12\]\[1\] cpu.regs\[13\]\[1\] cpu.regs\[14\]\[1\] cpu.regs\[15\]\[1\]
+ _00568_ _00804_ _00826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07033_ _02515_ _02524_ _02525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06008__A1 net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09045__I1 _04114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08984_ _02630_ _04069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07935_ cpu.spi.data_out_buff\[0\] _03243_ _03244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05636__I _01036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07866_ cpu.spi.div_counter\[5\] cpu.spi.divisor\[5\] _03186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09605_ _04333_ _04622_ _04637_ _04541_ _04403_ _04638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_39_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input19_I io_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07797_ cpu.spi.data_in_buff\[7\] _03106_ _03116_ _03119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06817_ _02305_ _02314_ _02315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_104_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09536_ _04570_ _04571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06748_ _02213_ _02214_ _02246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__05371__I _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09467_ _04313_ _04505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08418_ _03623_ _03592_ _03624_ _03616_ _00312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06679_ _02173_ _02176_ _02177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_81_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08682__I _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09398_ cpu.PC\[6\] _00754_ _04438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08349_ _03553_ _03572_ _00295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10311_ _00250_ clknet_leaf_39_wb_clk_i cpu.uart.div_counter\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_115_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09036__I1 _02561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10242_ _00181_ clknet_4_2_0_wb_clk_i cpu.regs\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_100_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10173_ _00112_ clknet_leaf_120_wb_clk_i cpu.regs\[12\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05525__A3 _01029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09672__A1 _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08592__I _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06238__A1 _00596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10509_ _00447_ clknet_leaf_82_wb_clk_i cpu.ROM_addr_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_110_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07738__A1 _03064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05981_ _01484_ _01485_ _01486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07720_ _03052_ _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07651_ _03010_ _00159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06287__I _01788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06602_ _00589_ _01015_ _02100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07582_ _02965_ _02967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05191__I _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09321_ _04027_ _04364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06533_ _02031_ _02032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06464_ net58 _01615_ _01963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09252_ _02802_ _04295_ _04296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_8_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08203_ cpu.uart.data_buff\[0\] _03460_ _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08218__A2 _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06395_ cpu.timer_div\[6\] _01631_ _01895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08435__C _03616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09183_ _04197_ _04205_ _04228_ _04229_ _04195_ _04230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05415_ _00904_ _00908_ _00915_ _00911_ _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_08134_ _03332_ _03403_ _03405_ _03406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05346_ cpu.PORTB_DDR\[1\] net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_16_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08065_ _03238_ _03348_ _03349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_clkbuf_leaf_33_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08451__B _03646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05277_ _00807_ _00809_ _00810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07016_ _00793_ _02509_ _00025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_113_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07729__A1 _00802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05366__I _00877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08967_ _03768_ _04054_ _00431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07918_ _03227_ _03102_ _03228_ _00208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08898_ _00734_ _03995_ _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07849_ cpu.timer\[10\] _03170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06197__I _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09519_ _03641_ _00771_ _04555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_72_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_61_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_61_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_14_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08209__A2 _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09301__I _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10016__A2 _02109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07432__A3 _02845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06640__A1 _00822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10225_ _00164_ clknet_leaf_108_wb_clk_i cpu.regs\[5\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10156_ _00095_ clknet_leaf_121_wb_clk_i cpu.regs\[14\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06943__A2 _02401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10087_ _00030_ clknet_leaf_111_wb_clk_i cpu.regs\[1\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09645__A1 _04114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05506__I0 _01010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05200_ _00733_ _00736_ _00737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06180_ _01681_ _01682_ _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05131_ cpu.mem_cycle\[1\] cpu.mem_cycle\[0\] _00670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_80_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05062_ _00603_ _00604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09870_ net56 _04853_ _04857_ _04858_ _04859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_0_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08821_ cpu.timer_capture\[11\] _03919_ _03938_ _03939_ _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08752_ _03174_ _03865_ _03866_ _03880_ _03881_ _03882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05964_ _01347_ _00866_ _01469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08683_ _03816_ _03825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07703_ cpu.regs\[3\]\[1\] _03041_ _03043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09884__A1 _04819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05895_ cpu.uart.has_byte _01193_ _01400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07634_ _02071_ _02982_ _02999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_75_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07565_ _02943_ cpu.regs\[10\]\[5\] _02948_ _02957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09304_ _04266_ _04347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07496_ _02911_ _00103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06516_ _01295_ _01352_ _01993_ _01340_ _01355_ _02015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_106_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09235_ _04233_ _04273_ _04277_ _04279_ _04280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06447_ _01599_ _01946_ _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09166_ _02792_ _04213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06378_ _01877_ _01302_ _01878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08117_ cpu.uart.div_counter\[4\] _03388_ _03237_ _03392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09097_ _04153_ _04138_ _04155_ _03980_ _00460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_71_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05329_ _00593_ _00853_ _00858_ _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_112_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08048_ _02824_ _03330_ _03331_ _01881_ _03333_ _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_10010_ _04745_ _04973_ _04971_ _04974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_8_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05096__I cpu.regs\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09999_ _00694_ _04681_ _04687_ _04963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_98_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08200__I _03450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09875__A1 _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06689__A1 cpu.regs\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09966__I net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10208_ _00147_ clknet_leaf_12_wb_clk_i cpu.regs\[7\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10139_ _00078_ clknet_leaf_103_wb_clk_i cpu.regs\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05275__S1 _00573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05680_ _01176_ _01186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07350_ _02790_ _00078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_116_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06301_ cpu.timer_top\[5\] _01802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_72_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07281_ _02648_ _02729_ _02738_ _02737_ _00061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09020_ _03614_ _04095_ _04096_ _04097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06232_ _01168_ _01732_ _01733_ _01267_ _00973_ _01734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_5_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06163_ _01663_ _01665_ _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_25_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05114_ cpu.instr_buff\[14\] _00653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_40_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06094_ _01549_ _01551_ _01597_ _01598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09922_ _00975_ _04889_ _04897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05045_ cpu.regs\[1\]\[4\] _00588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09853_ _02520_ _04846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09784_ cpu.ROM_spi_cycle\[3\] _04787_ _04790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08804_ _03920_ _03925_ _03926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06996_ _02448_ _02489_ _02490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08735_ _02707_ _03865_ _03866_ _03867_ _03856_ _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09857__A1 _04823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05947_ _01451_ _01452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08666_ cpu.timer_div_counter\[6\] _03809_ _03813_ _00371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05878_ _01189_ _01383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__08955__I _04043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08597_ cpu.pwm_counter\[0\] cpu.pwm_counter\[1\] cpu.pwm_counter\[2\] _03765_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_07617_ cpu.regs\[7\]\[1\] _02986_ _02989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07548_ _02946_ _00120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_63_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07479_ cpu.regs\[14\]\[7\] _02891_ _02901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10490_ _00428_ clknet_leaf_41_wb_clk_i cpu.uart.divisor\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09218_ _04260_ _04263_ _03853_ _00473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09149_ _01548_ _04196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_102_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06071__A2 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09026__I _00700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06850_ _02259_ _02346_ _02347_ _02348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__05464__I _00973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05801_ _01304_ _01305_ _01306_ _01307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09839__A1 _04022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06781_ _02248_ _02274_ _02275_ _02276_ _02277_ _02278_ _02279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
X_05732_ _01182_ _01231_ _01234_ _01237_ _01238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_08520_ cpu.toggle_ctr\[4\] _03706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08451_ _03647_ _03648_ _03646_ _00321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05663_ _01168_ _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07402_ _02834_ _02835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_58_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05594_ _01096_ _01099_ _01100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08382_ _03579_ _03598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07333_ _02602_ _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_98_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07264_ _02725_ _00057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08724__B _03529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_118_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_118_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06215_ net10 _01206_ _01201_ _01717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_104_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09003_ _04083_ _04084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07195_ _02665_ _02654_ _02666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05639__I _01144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06146_ _01276_ _01648_ _01649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06077_ net91 _00919_ _01581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09905_ _04884_ _00539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05028_ _00570_ _00571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09836_ _04683_ _04833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05374__I _00885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09767_ _04778_ _00507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06979_ _02472_ _02050_ _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_57_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09698_ _02452_ _04719_ _04721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08718_ _03848_ _03852_ _03853_ _00383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_69_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_107_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08649_ cpu.timer_div_counter\[0\] _03802_ _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_1_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10611_ _00549_ clknet_leaf_77_wb_clk_i cpu.ROM_spi_mode vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_37_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10542_ _00480_ clknet_leaf_97_wb_clk_i cpu.PC\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10473_ _00412_ clknet_leaf_31_wb_clk_i cpu.spi.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09230__A2 cpu.br_rel_dest\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07241__A1 cpu.timer_capture\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05993__B _01380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05284__I _00816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06000_ cpu.uart.divisor\[10\] _01503_ _01504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_70_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06283__A2 _01784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09221__A2 _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07232__A1 _00998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05469__S1 _00977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07951_ _02652_ _03242_ _03256_ _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06902_ _00591_ _02070_ _02400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07882_ _03184_ _03201_ _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09621_ _04169_ _04652_ _04653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06833_ _02325_ _02330_ _02331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09552_ _04312_ _04586_ _04587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06764_ _00935_ _00937_ _00942_ _00940_ _02261_ _02262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_05715_ _01214_ _01219_ _01220_ _01110_ _01221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_54_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07299__A1 _01261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08503_ _03683_ _03686_ _03688_ _03689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09483_ _04261_ _04520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08496__B1 _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06695_ _02191_ _02192_ _02193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08434_ cpu.orig_PC\[8\] _03611_ _03636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05646_ _01150_ _01151_ _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_05577_ _01055_ _01064_ _01072_ _01082_ _01083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_08365_ cpu.orig_IO_addr_buff\[2\] _03581_ _03585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07316_ cpu.toggle_top\[12\] _02761_ _02764_ _02756_ _02765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_116_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08296_ _03528_ _03530_ _00284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_104_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07247_ _02678_ _02710_ _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07178_ _02633_ _02651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06129_ cpu.spi.dout\[3\] _01611_ _01630_ _01631_ _01632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_41_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_86_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_86_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08971__B2 _02692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_15_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_15_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_6_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09819_ _04819_ _04816_ _04820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput17 io_in[28] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput28 sram_out[2] net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_64_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10525_ _00463_ clknet_leaf_81_wb_clk_i cpu.last_addr\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10456_ _00395_ clknet_leaf_24_wb_clk_i cpu.timer\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10387_ _00326_ clknet_leaf_10_wb_clk_i cpu.toggle_top\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10300__D _00239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06480_ cpu.timer_capture\[15\] _01233_ _01639_ _01979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05500_ cpu.regs\[12\]\[5\] cpu.regs\[13\]\[5\] cpu.regs\[14\]\[5\] cpu.regs\[15\]\[5\]
+ _00887_ _00879_ _01008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_114_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05431_ _00905_ _00941_ _00913_ _00942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_08150_ _03400_ _03418_ _00250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08274__B _03381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07101_ _02379_ _02587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05362_ _00873_ _00874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_113_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08081_ _03098_ _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05293_ _00819_ _00824_ _00579_ _00825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_113_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_23_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07032_ net12 _02516_ _02524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_3_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08983_ _01279_ _04039_ _04041_ _04067_ _04059_ _04068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_11_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07934_ _03230_ _03243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07865_ cpu.spi.div_counter\[0\] cpu.spi.divisor\[0\] _03185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_98_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09604_ _00606_ _04614_ _04636_ _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07796_ _01880_ _03113_ _03118_ _00196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06816_ _02308_ _02312_ _02313_ _02314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_104_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09535_ _03089_ _04568_ _04569_ _04570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_39_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06747_ _02239_ _02244_ _02245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09466_ _00777_ _04503_ _04504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06678_ _00604_ _00995_ _02175_ _02176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_19_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_62_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08417_ cpu.orig_PC\[3\] _03611_ _03624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05378__S0 _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05629_ _01033_ _01132_ _01134_ _01135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_62_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09397_ cpu.PC\[6\] _01037_ _04437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_19_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08348_ cpu.uart.receive_div_counter\[15\] _03567_ _03571_ _03572_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_34_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07444__A1 _02845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08279_ _03425_ _03516_ _00281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_73_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10310_ _00249_ clknet_leaf_38_wb_clk_i cpu.uart.div_counter\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10241_ _00180_ clknet_leaf_107_wb_clk_i cpu.regs\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_100_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05758__A1 _01261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10172_ _00111_ clknet_leaf_122_wb_clk_i cpu.regs\[12\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05302__S0 _00570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05930__A1 cpu.Z vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06238__A2 _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10508_ _00446_ clknet_leaf_82_wb_clk_i cpu.ROM_addr_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09188__A1 cpu.Z vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10439_ _00378_ clknet_leaf_19_wb_clk_i cpu.timer_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_107_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08935__A1 _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05980_ _01463_ _01483_ _01485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09360__A1 _00590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07650_ _03009_ cpu.regs\[6\]\[5\] _02999_ _03010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07910__A2 _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06601_ _00603_ _02083_ _02099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07581_ _01701_ _02966_ _00133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09879__I _04864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09320_ _04358_ _04361_ _04362_ _04363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06532_ _01370_ _01989_ _02028_ _02030_ _02031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_34_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09251_ _02795_ _02782_ _04295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06463_ cpu.uart.divisor\[7\] _01962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_08202_ _03459_ _03460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06394_ _01880_ _01188_ _01892_ _01893_ _01184_ _01894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_09182_ _03604_ _04031_ _04197_ _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05414_ _00924_ _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_8_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08133_ _03332_ _03404_ _03397_ _03405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__07426__B2 _02629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05345_ cpu.PORTB_DDR\[0\] net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_43_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08064_ _03222_ _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_70_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07015_ net54 _02496_ _02508_ _02509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09179__A1 cpu.Z vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05276_ _00002_ _00808_ _00003_ _00809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_101_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08023__I net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input31_I sram_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08966_ _01073_ _04038_ _04053_ _04050_ _04054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07917_ _00746_ cpu.spi.busy _03228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08897_ _02626_ _01155_ _00722_ _03994_ _03995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_98_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07848_ cpu.timer_top\[7\] _02720_ _03168_ _03169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06165__A1 _01437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07779_ _03106_ _03107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09103__A1 _04114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09789__I net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09518_ _04028_ _04546_ _04554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09449_ _04338_ _04487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07432__A4 _02864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_30_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_30_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_50_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08917__A1 _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10224_ _00163_ clknet_leaf_12_wb_clk_i cpu.regs\[5\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10155_ _00094_ clknet_leaf_123_wb_clk_i cpu.regs\[14\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10086_ _00029_ clknet_leaf_92_wb_clk_i cpu.instr_buff\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07353__B1 _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05903__A1 cpu.timer_div\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05130_ cpu.mem_cycle\[5\] cpu.mem_cycle\[4\] cpu.mem_cycle\[3\] cpu.mem_cycle\[2\]
+ _00669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_52_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05061_ cpu.regs\[1\]\[5\] _00603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08384__A2 _03596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08820_ _03794_ _03939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06395__A1 cpu.timer_div\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08751_ _03840_ _03881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05963_ _01467_ _01450_ _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05894_ _01195_ _01397_ _01398_ _01399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08682_ _03816_ _03824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_49_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06147__A1 _00988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07702_ _01373_ _03040_ _03042_ _00178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07633_ _02997_ _02986_ _02998_ _00153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09636__A2 cpu.ROM_addr_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07564_ _02956_ _00126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09303_ _04292_ _04346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07495_ _01875_ cpu.regs\[13\]\[5\] _02902_ _02911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06515_ net97 _02013_ _02014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08018__I _02617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09234_ _04278_ _04265_ _04233_ _04279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06446_ net96 _01365_ _01945_ _01946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_118_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05122__A2 _00655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09165_ _01304_ _02185_ _02109_ _02615_ _04212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_8_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08116_ cpu.uart.div_counter\[4\] _03374_ _03389_ _03390_ _03391_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06377_ _01155_ _01877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09096_ cpu.ROM_addr_buff\[4\] _04154_ _04155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05328_ _00855_ _00857_ _00593_ _00858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08047_ _03332_ _01962_ cpu.uart.divisor\[1\] _03320_ _03333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_05259_ cpu.IE _00794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_31_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09572__A1 _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09998_ _04942_ _04960_ _04962_ _04231_ _00554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_08949_ _04037_ _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06138__A1 cpu.timer_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06689__A2 _01994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07810__B2 _01976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07810__A1 cpu.timer_div\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10207_ _00146_ clknet_leaf_13_wb_clk_i cpu.regs\[7\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10138_ _00077_ clknet_leaf_106_wb_clk_i _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10069_ _02032_ _05014_ _05022_ _00565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07280_ cpu.timer_top\[3\] _02730_ _02738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06300_ _01800_ _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_73_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06231_ cpu.toggle_top\[12\] _01262_ _01733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_31_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09097__C _03980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06162_ _01563_ _01567_ _01664_ _01665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_111_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05113_ cpu.br_rel_dest\[5\] _00652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_13_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06093_ _01552_ _01571_ _01588_ _01596_ _01597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_111_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09921_ _04896_ _00543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05044_ _00586_ _00587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09852_ _04819_ _04842_ _04845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09783_ cpu.ROM_spi_cycle\[3\] _04787_ _04789_ _00512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08803_ _03174_ _03922_ _03924_ _03925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06995_ _02455_ _02460_ _02465_ _02488_ _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_08734_ _02707_ _03860_ _03867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09306__A1 _03623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05946_ _01338_ _01359_ _01451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08665_ cpu.timer_div_counter\[6\] _03809_ _03811_ _03812_ _03813_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05877_ _01248_ _01382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09560__C _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09609__A2 _03995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08596_ _03759_ _03760_ _03763_ _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07616_ _01493_ _02988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_62_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07547_ _02945_ cpu.regs\[11\]\[6\] _02933_ _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_52_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07478_ _02900_ _00096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09217_ _02783_ _04262_ _04263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06429_ net95 _01774_ _01929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09148_ _04194_ _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06491__I _00646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09079_ _04141_ _04142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_15_Left_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output62_I net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_24_Left_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09470__C _04309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06531__A1 _01370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09977__I net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08881__I _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_33_Left_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_112_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06598__A1 _02090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_42_Left_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05800_ _01033_ _01306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06780_ _02246_ _02247_ _02274_ _02278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_117_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05731_ cpu.timer_capture\[0\] _01236_ _01237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_77_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08450_ cpu.orig_PC\[12\] _03642_ _03648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05662_ _01121_ _01168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06576__I _02072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07401_ cpu.uart.receive_div_counter\[0\] _02834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08381_ _03593_ _03597_ _03570_ _00302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05480__I _00988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05593_ _01071_ _01098_ _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_46_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07332_ _02777_ _00073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_51_Left_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07078__A2 _02565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07263_ cpu.timer_capture\[7\] _02701_ _02724_ _02712_ _02725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_61_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06214_ net2 _01390_ _01713_ _01715_ _01110_ _01716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__08027__B2 _01881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09002_ _02536_ _03050_ _04082_ _02511_ _04083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_07194_ _02664_ _02665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_60_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09775__A1 _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10047__B _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07200__I _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06145_ _01168_ _01645_ _01647_ _01267_ _00956_ _01648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_41_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07625__I1 cpu.regs\[7\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06076_ _01558_ _01580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09904_ cpu.PORTB_DDR\[6\] _04876_ _04883_ _04881_ _04884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05261__A1 _00794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05027_ _00569_ _00570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09835_ _04018_ _04829_ _04832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09766_ cpu.ROM_spi_dat_out\[6\] _04760_ _04777_ _04765_ _04778_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06978_ cpu.mem_cycle\[1\] _02472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_57_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09697_ _04720_ _00495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08717_ _03609_ _03853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05929_ _01424_ _01428_ _01433_ _01434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_107_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08648_ _03801_ _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08502__A2 cpu.toggle_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06513__A1 _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05390__I _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08579_ cpu.toggle_ctr\[12\] _03751_ _03753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_37_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10610_ _00548_ clknet_leaf_57_wb_clk_i cpu.PORTA_DDR\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10541_ _00479_ clknet_leaf_93_wb_clk_i cpu.PC\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10472_ _00411_ clknet_leaf_30_wb_clk_i cpu.spi.divisor\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07110__I _02517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09518__A1 _04028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08876__I _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_4_2_0_wb_clk_i clknet_0_wb_clk_i clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_83_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_13_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05491__A1 _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07950_ cpu.spi.data_out_buff\[3\] _03243_ _03256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06901_ _01788_ _02073_ _02398_ _02399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07881_ _03105_ _03200_ _03201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09620_ cpu.last_addr\[9\] cpu.last_addr\[8\] _04651_ _04652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06832_ _02326_ _02328_ _02329_ _02330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09551_ _04368_ _04575_ _04584_ _04585_ _04586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06763_ _00834_ _02261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_05714_ net21 _01053_ _01220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_54_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08502_ _03687_ cpu.toggle_top\[13\] cpu.toggle_top\[12\] _03684_ _03688_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_66_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09482_ _04486_ _04519_ _04484_ _00481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06694_ _02153_ _02154_ _02192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_52_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08433_ _03634_ _03635_ _03630_ _00316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05645_ _00715_ _00866_ _01151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_05576_ _01076_ _01081_ _01082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08364_ _01071_ _03580_ _03584_ _03583_ _00298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_62_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07315_ _02762_ _02763_ _02764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10055__A1 _01373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08295_ cpu.uart.receive_div_counter\[4\] _03526_ _03529_ _03530_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07246_ _02707_ _02703_ _02709_ _02710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09048__I0 cpu.regs\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07471__A2 _02891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07177_ _02650_ _00045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06128_ _01183_ _01631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06059_ _01160_ _01550_ _01563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_6_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09920__A1 cpu.PORTA_DDR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09818_ _00921_ _04819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05537__A2 net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_91_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09749_ _04683_ _04765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_55_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_55_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_96_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08239__A1 _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput18 io_in[29] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_52_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput29 sram_out[3] net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10524_ _00462_ clknet_leaf_81_wb_clk_i cpu.last_addr\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09039__I0 _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10455_ _00394_ clknet_leaf_24_wb_clk_i cpu.timer\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10386_ _00325_ clknet_leaf_10_wb_clk_i cpu.toggle_top\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05225__A1 _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05084__S0 _00600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08478__A1 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05430_ cpu.regs\[12\]\[2\] cpu.regs\[13\]\[2\] cpu.regs\[14\]\[2\] cpu.regs\[15\]\[2\]
+ _00878_ _00879_ _00941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_55_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10037__A1 _01466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10037__B2 _01462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05361_ _00005_ _00873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07100_ _02571_ _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_99_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08080_ _03346_ _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_82_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05292_ cpu.regs\[0\]\[1\] _00822_ _00823_ cpu.regs\[3\]\[1\] _00568_ _00804_ _00824_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07031_ _02523_ _00026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08402__A1 _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08982_ cpu.orig_IO_addr_buff\[4\] _04056_ _04057_ _00989_ _04067_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05311__S1 _00574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07933_ _03241_ _03242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07864_ _00686_ _03183_ _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_97_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09603_ _04614_ _04622_ _04636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_39_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06815_ _02309_ _02310_ _02311_ _02313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07795_ cpu.spi.data_in_buff\[6\] _03106_ _03116_ _03118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_104_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09534_ _02390_ _04407_ _04569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06746_ _02242_ _02243_ _02244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_66_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09465_ _04413_ _04491_ _04503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06677_ _02173_ _02174_ _02175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_19_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08416_ _03622_ _03623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05378__S1 _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05628_ _01133_ _01128_ _01134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09396_ _04434_ _04435_ _04436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08347_ cpu.uart.receive_div_counter\[15\] _03513_ _03565_ _03571_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_74_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05559_ cpu.IO_addr_buff\[1\] _01065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07444__A2 _02864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08278_ _02833_ _03514_ _03515_ _02869_ _03516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08641__A1 _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_102_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_102_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_104_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07229_ _02695_ _00052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10240_ _00179_ clknet_leaf_107_wb_clk_i cpu.regs\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_100_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10171_ _00110_ clknet_leaf_123_wb_clk_i cpu.regs\[12\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05302__S1 _00574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_110_Right_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06707__A1 cpu.regs\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07263__C _02712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07380__A1 _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05930__A2 _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05694__A1 _01196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10019__A1 _01354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_7_Left_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10507_ _00445_ clknet_leaf_82_wb_clk_i cpu.ROM_addr_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_110_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10438_ _00377_ clknet_leaf_19_wb_clk_i cpu.timer_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05049__I1 _00590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10369_ _00308_ clknet_leaf_90_wb_clk_i cpu.orig_flags\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09653__C _04684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06600_ _02082_ _02097_ _02098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07580_ _01603_ _02966_ _00132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10502__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06531_ _01370_ _02029_ _02030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09250_ _04266_ _04294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_0_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_0_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06462_ cpu.spi.dout\[7\] _01961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08201_ _03457_ _03458_ _03232_ _03459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_44_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06393_ cpu.spi.divisor\[6\] _01628_ _01610_ _01893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_56_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09181_ _04181_ _04208_ _04220_ _04227_ _04228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_7_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05413_ _00719_ _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08132_ _03371_ _03404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09895__I _04864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05344_ cpu.PORTA_DDR\[2\] net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_43_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08063_ _03346_ _03347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05437__A1 _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05275_ cpu.regs\[4\]\[0\] cpu.regs\[5\]\[0\] cpu.regs\[6\]\[0\] cpu.regs\[7\]\[0\]
+ _00803_ _00573_ _00808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_113_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07014_ _02496_ _02498_ _02507_ _02508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_71_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05988__A2 _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08965_ _01377_ _04039_ _04041_ _04052_ _04047_ _04053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05296__S0 _00568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07916_ _03226_ _03227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_110_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input24_I io_in[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08896_ _00700_ _01025_ _00757_ _03994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_07847_ _01960_ cpu.timer\[7\] _03167_ _03168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07778_ _03105_ _03106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_65_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09517_ _04358_ _04546_ _04552_ _00776_ _04553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06729_ _02222_ _02223_ _02227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08862__A1 _02665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09448_ _04485_ _04344_ _04486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07665__A2 _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09379_ _02562_ _04317_ _04420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07417__A2 _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08642__C _03795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08090__A2 _03368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output92_I net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09754__B _03761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10223_ _00162_ clknet_leaf_13_wb_clk_i cpu.regs\[5\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06928__A1 _02407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_70_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_70_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05287__S0 _00803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10154_ _00093_ clknet_leaf_0_wb_clk_i cpu.regs\[14\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10085_ _00028_ clknet_leaf_92_wb_clk_i cpu.instr_buff\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06669__I _00801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07353__B2 _02327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07105__A1 _02407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08853__A1 cpu.spi.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07656__A2 _03002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07168__C _00791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05060_ cpu.regs\[4\]\[5\] cpu.regs\[5\]\[5\] cpu.regs\[6\]\[5\] cpu.regs\[7\]\[5\]
+ _00600_ _00601_ _00602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_111_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09581__A2 _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08750_ _03174_ _03879_ _03880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05483__I _00991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06579__I _02076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05962_ net90 _01354_ _01467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05893_ cpu.uart.dout\[1\] _00012_ _01398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08681_ _02648_ _03817_ _03823_ _03820_ _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_49_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07344__A1 _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07701_ cpu.regs\[3\]\[0\] _03041_ _03042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07912__B _03223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07632_ cpu.regs\[7\]\[7\] _02984_ _02998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09302_ _02811_ _04344_ _04345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07563_ _02941_ cpu.regs\[10\]\[4\] _02949_ _02956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08844__A1 _03232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07494_ _02910_ _00102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06514_ _00616_ _00632_ _01774_ _02013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_118_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09233_ _00991_ _04235_ _04278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06445_ _01922_ _01928_ _01938_ _01944_ _01945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_28_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_15_0_wb_clk_i clknet_0_wb_clk_i clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_90_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05122__A3 _00658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09164_ _00748_ _01430_ _04210_ _04211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_8_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08115_ _03377_ _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06376_ _01876_ _00018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09095_ _04136_ _04154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05327_ _00581_ _00856_ _00857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05258_ _00792_ _00793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08046_ cpu.uart.div_counter\[7\] _03332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06083__B2 _01462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06083__A1 _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05189_ cpu.instr_cycle\[2\] _00726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08969__I _04043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05830__A1 _01269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09572__A2 _00772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09997_ _04910_ _04961_ _04960_ _02494_ _04962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_08948_ _04030_ _04036_ _02630_ _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05393__I _00006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08879_ cpu.timer_div\[3\] _03976_ _03981_ _03956_ _03982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_98_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_88_Left_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07638__A2 _03002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06310__A2 _01205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_97_Left_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09012__A1 _02527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10206_ _00145_ clknet_leaf_124_wb_clk_i cpu.regs\[8\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07574__A1 _01175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10137_ _00076_ clknet_leaf_106_wb_clk_i _00006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10068_ cpu.regs\[15\]\[7\] _05012_ _05022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08523__B1 cpu.toggle_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07877__A2 cpu.spi.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08826__A1 cpu.timer_capture\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07023__I _00733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06230_ cpu.toggle_top\[4\] _01255_ _01731_ _01258_ _01732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_26_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06161_ _01160_ _01551_ _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_25_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05112_ net25 _00651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06092_ _01590_ _01592_ _01594_ _01595_ _01596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_09920_ cpu.PORTA_DDR\[2\] _04888_ _04895_ _04893_ _04896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05812__A1 _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05043_ _00002_ _00586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09851_ _04844_ _00525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_111_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09782_ cpu.ROM_spi_cycle\[3\] _04787_ _00790_ _04789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06994_ _02478_ _02480_ _02487_ _02488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08802_ _02635_ _03923_ _03924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08733_ _03833_ _03866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05945_ _01441_ _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06102__I cpu.br_rel_dest\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08664_ _02660_ _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05876_ _01377_ _01378_ _01380_ _01381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08595_ cpu.pwm_counter\[2\] _03763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05423__S0 _00872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07615_ _02980_ _02985_ _02987_ _00146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07546_ _01949_ _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_24_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09216_ _04261_ _04262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_52_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07477_ _01951_ cpu.regs\[14\]\[6\] _02890_ _02900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_106_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06428_ _01479_ _01926_ _01927_ _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09147_ _00727_ _03594_ _04194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06359_ _01837_ _01858_ _01470_ _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07089__B _02063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09078_ _00693_ _04140_ _04141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08029_ _02853_ _03310_ _03311_ cpu.uart.divisor\[2\] _03314_ _03315_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_73_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05582__A3 _01087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07271__C _00791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08284__A2 _03510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08036__A2 _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09233__A1 _00991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06770__A2 _00917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05730_ _01054_ _01076_ _01235_ _01236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__05761__I _01266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_42_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05661_ _01166_ _01167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07400_ cpu.uart.receive_div_counter\[1\] _02833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08380_ cpu.orig_IO_addr_buff\[5\] _03596_ _03597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05592_ _00648_ _01098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07331_ cpu.toggle_top\[15\] _02761_ _02776_ _02773_ _02777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_42_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07262_ _02720_ _02703_ _02691_ _02723_ _02724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06213_ _01218_ _01714_ _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09001_ _00697_ _03050_ _04082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07193_ _01801_ _02664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06144_ _01646_ _01262_ _01647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06075_ _01465_ _01579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09903_ _04022_ _04877_ _04883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09408__I _04309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05026_ _00568_ _00569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09834_ _04831_ _00521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_81_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09765_ _04755_ _04776_ _04777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06977_ _02466_ _02469_ _02470_ _02471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_29_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09696_ _03247_ _04717_ _04719_ _04720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_08716_ _03836_ _03850_ _03851_ _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_57_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05928_ _01429_ _01432_ _01146_ _01433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_107_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08647_ _03121_ _03800_ _03801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_1_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05859_ _00656_ _01365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08578_ cpu.toggle_ctr\[12\] _03751_ _03752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_37_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07529_ _02933_ _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10540_ _00478_ clknet_4_9_0_wb_clk_i cpu.PC\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10471_ _00410_ clknet_leaf_28_wb_clk_i cpu.spi.divisor\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06029__A1 cpu.timer_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07701__A1 cpu.regs\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_126_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05491__A2 _00974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_9_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05756__I _01106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06900_ _02074_ _02397_ _02398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07880_ _03199_ _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06831_ _02288_ _00929_ _02329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_37_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09550_ _04358_ _04570_ _00776_ _04585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06762_ _02245_ _02257_ _02260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05713_ net59 _01215_ _01218_ _01219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09481_ _04487_ _04512_ _04517_ _04518_ _04519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_54_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08501_ cpu.toggle_ctr\[13\] _03687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08432_ cpu.orig_PC\[7\] _03628_ _03635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08496__A2 _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06693_ _02183_ _02190_ _02191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05644_ _00717_ _00950_ _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_05575_ _01080_ _01081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08363_ cpu.orig_IO_addr_buff\[1\] _03581_ _03584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_34_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08294_ _03236_ _03529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_85_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07314_ _02748_ _02763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06259__A1 _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07245_ _02708_ _02697_ _02709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09048__I1 _02588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07176_ cpu.uart.divisor\[3\] _02634_ _02649_ _02639_ _02650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_14_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06127_ _01627_ _01629_ _01188_ _01630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05234__A2 _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06431__A1 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06058_ _01559_ _01561_ _01562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_111_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_70_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09817_ _04818_ _00517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09748_ _04751_ _04763_ _04764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05537__A3 _00661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09679_ _04704_ _04705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_96_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_24_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_24_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08645__C _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput19 io_in[2] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_91_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10523_ _00461_ clknet_leaf_82_wb_clk_i cpu.last_addr\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09039__I1 _02563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10454_ _00393_ clknet_leaf_24_wb_clk_i cpu.timer\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_70_Left_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10385_ _00324_ clknet_leaf_8_wb_clk_i cpu.toggle_clkdiv vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06422__A1 _01325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05084__S1 _00601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05784__I0 cpu.regs\[12\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06489__B2 _01957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06489__A1 _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05360_ _00871_ _00872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_31_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05291_ cpu.regs\[2\]\[1\] _00823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_113_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07030_ _00769_ _02514_ _02518_ _02522_ _02523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_2_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06091__B _01479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08981_ _04037_ _04066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07932_ _03229_ _03239_ _03241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08797__I _03918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07863_ _03104_ _03182_ _03183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09602_ _04294_ _04622_ _04634_ _04331_ _04635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_39_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06814_ _02309_ _02310_ _02311_ _02312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_07794_ _01803_ _03107_ _03117_ _00195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_64_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09533_ _02389_ _04408_ _04568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_104_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06745_ _02108_ _00995_ _02243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06676_ _00637_ _00929_ _02172_ _02174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_19_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09464_ _04497_ _04500_ _04501_ _04502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_93_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09395_ cpu.PC\[5\] cpu.br_rel_dest\[5\] _04416_ _04435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05627_ _01040_ _01133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08415_ _02382_ _03622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_117_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08346_ _03568_ _03569_ _03570_ _00294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_62_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05558_ _01056_ _01059_ _01063_ _01064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08277_ _02833_ _02835_ _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_61_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05489_ _00997_ _00998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07228_ cpu.timer_capture\[2\] _02674_ _02694_ _02687_ _02695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_6_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07159_ _02635_ _02636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06404__A1 cpu.toggle_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10170_ _00109_ clknet_leaf_126_wb_clk_i cpu.regs\[12\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05143__A1 _00675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_69_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09409__A1 _01877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05694__A2 _01199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06891__A1 cpu.PC\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10506_ _00444_ clknet_leaf_83_wb_clk_i cpu.ROM_addr_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_52_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10437_ _00376_ clknet_leaf_23_wb_clk_i cpu.timer_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_78_Right_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10368_ _00307_ clknet_leaf_86_wb_clk_i cpu.orig_flags\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05049__I2 _00591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10299_ _00238_ clknet_leaf_63_wb_clk_i cpu.spi.counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_108_Left_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09896__A1 _04014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07026__I _00685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_87_Right_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06530_ net33 _01309_ _02029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08285__C _03414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06461_ cpu.timer_top\[7\] _01960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_47_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08200_ _03450_ _03458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05412_ _00923_ net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_44_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_117_Left_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06392_ cpu.uart.dout\[6\] _01194_ _01889_ _01891_ _01101_ _01892_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_09180_ _04222_ _04226_ _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_44_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08131_ _03371_ _03401_ _03402_ _03403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05343_ cpu.PORTA_DDR\[1\] net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_71_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08062_ _02735_ _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05437__A2 _00933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05274_ _00579_ _00806_ _00807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07013_ _02499_ _02504_ _02460_ _02506_ _02507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XPHY_EDGE_ROW_96_Right_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08964_ cpu.orig_IO_addr_buff\[1\] _04044_ _04045_ _02642_ _04052_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_110_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07915_ _00688_ _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05944__I _01360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08895_ _03993_ _00420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07846_ _03164_ _03165_ _03166_ _03167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input17_I io_in[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07777_ _03104_ _03105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09516_ _04306_ _04551_ _04552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06728_ _02225_ _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_93_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09447_ cpu.PC\[8\] _04485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_39_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06659_ _02123_ _02124_ _02157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09378_ _04413_ _04417_ _04418_ _04368_ _04419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08329_ _03553_ _03556_ _00291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09811__A1 _01087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10222_ _00161_ clknet_leaf_116_wb_clk_i cpu.regs\[6\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05287__S1 _00573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06928__A2 _02408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10153_ _00092_ clknet_leaf_2_wb_clk_i cpu.regs\[14\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09878__A1 _01122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07274__C _00791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10084_ _00027_ clknet_leaf_92_wb_clk_i cpu.base_address\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05364__A1 _00870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07353__A2 _01022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06864__A1 _02361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07041__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05278__S1 _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input9_I io_in[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05961_ _01465_ _01466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07700_ _03038_ _03041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05892_ _01396_ cpu.uart.divisor\[9\] _01198_ _01397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08680_ cpu.timer_top\[11\] _03818_ _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_49_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07912__C _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07631_ _02031_ _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07562_ _02925_ _02950_ _02955_ _00125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09301_ _04261_ _04344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06513_ _01675_ _02011_ _02012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07493_ _01789_ cpu.regs\[13\]\[4\] _02903_ _02910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09232_ _04274_ _04276_ _04277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06444_ _01939_ _01943_ _01944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05658__A2 _01153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09163_ _01953_ _01154_ _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_8_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06375_ _01875_ cpu.regs\[9\]\[5\] _01702_ _01876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08114_ cpu.uart.div_counter\[4\] _03388_ _03389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05326_ cpu.regs\[8\]\[3\] cpu.regs\[9\]\[3\] cpu.regs\[10\]\[3\] cpu.regs\[11\]\[3\]
+ _00846_ _00847_ _00856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09094_ cpu.last_addr\[4\] _04153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_114_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05257_ _00745_ _00792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08045_ cpu.uart.div_counter\[6\] _03331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07280__A1 cpu.timer_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05188_ _00723_ _00724_ _00725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__07032__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09996_ _04929_ _04944_ _04957_ _04961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07583__A2 _02967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08947_ _04031_ _04035_ _04036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08878_ _02758_ _03973_ _03981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07829_ _01609_ cpu.timer\[11\] cpu.timer\[10\] _03147_ _03150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_79_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05849__I _00720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07271__A1 _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10205_ _00144_ clknet_leaf_119_wb_clk_i cpu.regs\[8\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08771__A1 cpu.timer_capture\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07574__A2 _01215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10136_ _00075_ clknet_leaf_112_wb_clk_i _00005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_89_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10067_ _05021_ _00564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_32_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06160_ _01661_ _01662_ _01663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05111_ _00649_ _00650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06091_ _01580_ _01593_ _01479_ _01595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05042_ _00583_ _00584_ _00585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_111_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09850_ net79 _04841_ _04843_ _04833_ _04844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_clkbuf_leaf_71_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09781_ _04787_ _04788_ _00511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06993_ _00695_ _02482_ _02486_ _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08801_ _03921_ _03923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07923__B _03232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08732_ _03137_ _03865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05944_ _01360_ _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08663_ _03137_ _03811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05875_ _01379_ _01380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08594_ _03759_ _03760_ _03762_ _00350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05423__S1 _00874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07614_ cpu.regs\[7\]\[0\] _02986_ _02987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_62_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07545_ _02944_ _00119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07476_ _02899_ _00095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_24_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09215_ _01026_ _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06427_ _01923_ _01925_ _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09146_ _04074_ _04193_ _00471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06358_ _01850_ _01858_ _01859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09077_ _00669_ _04134_ _04140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09585__B _00690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06289_ _01790_ _00017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05309_ cpu.regs\[12\]\[2\] cpu.regs\[13\]\[2\] cpu.regs\[14\]\[2\] cpu.regs\[15\]\[2\]
+ _00569_ _00805_ _00840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08028_ cpu.uart.div_counter\[7\] _01962_ _01612_ cpu.uart.div_counter\[3\] _03313_
+ _03314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xclkbuf_leaf_49_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_49_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_4_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09979_ _04916_ _02599_ _04943_ _04640_ _04944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_98_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06516__B1 _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_105_Right_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_84_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_116_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09479__C _04292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08992__B2 _01957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10119_ _00062_ clknet_leaf_20_wb_clk_i cpu.timer_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05660_ _01137_ _01165_ _01166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05591_ _01096_ _01075_ _01097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__05730__A1 _01054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07330_ _02775_ _02763_ _02776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07261_ _02679_ _02722_ _02723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09000_ _04074_ _04081_ _00437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05489__I _00997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06212_ net63 _01515_ _01714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_98_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07192_ _02663_ _00047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06143_ cpu.toggle_top\[11\] _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_13_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08983__A1 _01279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06074_ _01574_ _01577_ _01578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05797__A1 _01299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09902_ _04882_ _00538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05025_ _00000_ _00568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09833_ net63 _04828_ _04830_ _04821_ _04831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06113__I _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07209__I _02673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09764_ cpu.ROM_spi_dat_out\[5\] _04731_ _04762_ _04775_ _04776_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06976_ _02056_ _02058_ _02470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_29_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09695_ _02453_ _04718_ _02039_ _02447_ _04719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_96_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08715_ _02684_ _03838_ _02690_ _03851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_57_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05927_ _01430_ _01431_ _01432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_107_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08646_ _03137_ _03800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09160__A1 _00921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05858_ _01337_ _01342_ _01357_ _01363_ _01364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__05721__A1 cpu.uart.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08577_ _03726_ _03750_ _03751_ _00344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05789_ _01294_ _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_37_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07528_ _01165_ _02932_ _02933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_106_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07459_ _01148_ _01153_ _02888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_91_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10470_ _00409_ clknet_leaf_31_wb_clk_i cpu.spi.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_51_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07226__A1 _02692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09129_ _04032_ _04178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_32_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05862__I _01157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05960__A1 _00863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07701__A2 _03041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07217__A1 _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09206__A2 _01020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10599_ _00537_ clknet_leaf_71_wb_clk_i cpu.PORTB_DDR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08965__A1 _01377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05779__A1 _01279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07029__I _02521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10210__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06830_ _02078_ _00895_ _00955_ _02327_ _02328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06761_ _02235_ _02258_ _02259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05951__A1 _00831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05712_ _01217_ _01218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09142__A1 _00946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09480_ _02530_ _04492_ _04195_ _04518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_54_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08500_ _03684_ cpu.toggle_top\[12\] cpu.toggle_top\[11\] _03685_ _03686_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06692_ _02184_ _02189_ _02190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08431_ _02588_ _03633_ _03634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05643_ _00654_ _00713_ _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05574_ _01077_ _01079_ _01080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08362_ _01074_ _03580_ _03582_ _03583_ _00297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_19_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07456__A1 _02521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08293_ cpu.uart.receive_div_counter\[4\] _03525_ _03527_ _03520_ _03528_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_73_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07313_ _01005_ _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_62_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07244_ _01707_ _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_6_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07175_ _02648_ _02637_ _02649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05947__I _01451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06126_ cpu.spi.divisor\[3\] _01628_ _01629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06057_ _01455_ _01560_ _01561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09381__A1 _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09816_ net59 _04814_ _04817_ _04765_ _04818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_94_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09747_ cpu.ROM_spi_dat_out\[1\] _04731_ _04761_ _04762_ _04763_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06959_ cpu.startup_cycle\[2\] _02453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05537__A4 _00672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05942__A1 _01326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09133__A1 _04178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09678_ _02450_ _04703_ _04704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_68_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07603__S _02968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08629_ _03777_ _03788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_83_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09436__A2 _04043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_64_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_64_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_91_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10522_ _00460_ clknet_leaf_81_wb_clk_i cpu.last_addr\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10453_ _00392_ clknet_leaf_8_wb_clk_i cpu.timer\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06670__A2 _00894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10384_ _00323_ clknet_leaf_60_wb_clk_i cpu.had_int vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09427__A2 _02626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07312__I _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05290_ _00821_ _00822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08143__I _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07610__A1 _02932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08980_ _04055_ _04065_ _00433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07931_ _03235_ _03240_ _00209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07862_ _00726_ _00681_ _00765_ _01086_ _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_48_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09601_ _00751_ _04356_ _04631_ _04633_ _04634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_39_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06813_ _02167_ _00993_ _02311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07793_ cpu.spi.data_in_buff\[5\] _03108_ _03116_ _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09532_ _03090_ _04520_ _04567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06744_ _00918_ _02238_ _02241_ _02242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09130__A4 _01279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09463_ _04497_ _04500_ _04306_ _04501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06675_ _00637_ _00928_ _02172_ _02173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__07677__A1 _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08318__I _03510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08414_ _03620_ _03621_ _03610_ _00311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09394_ cpu.PC\[5\] _00706_ _04434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05626_ _01131_ _01127_ _00868_ _01132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08345_ _03226_ _03570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_74_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05557_ _01062_ _01063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_58_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08276_ _02834_ _03513_ _02871_ _03514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05488_ _00996_ _00997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_34_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07227_ _02690_ _02677_ _02691_ _02693_ _02694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_61_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08929__A1 cpu.uart.divisor\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07158_ _01429_ _02635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09149__I _01548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06109_ cpu.uart.divisor\[3\] _01612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_14_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07089_ net19 _02405_ _02063_ _02576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_100_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_4_4_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_111_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_111_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05626__B _00868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05915__A1 _01419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07132__I _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10505_ _00443_ clknet_leaf_87_wb_clk_i cpu.ROM_addr_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07840__A1 cpu.timer_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07840__B2 cpu.timer_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10436_ _00375_ clknet_leaf_10_wb_clk_i cpu.timer_top\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_100_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10367_ _00306_ clknet_leaf_91_wb_clk_i cpu.orig_flags\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05049__I3 cpu.regs\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10298_ _00237_ clknet_leaf_66_wb_clk_i cpu.spi.counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06460_ cpu.pwm_top\[7\] _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05411_ _00865_ _00896_ _00922_ _00923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_44_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06331__A1 _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08130_ _03369_ _03402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06391_ _00684_ _01890_ _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05342_ cpu.PORTA_DDR\[0\] net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_70_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08061_ _03309_ _03340_ _03341_ _00239_ _00233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05437__A3 _00947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05273_ cpu.regs\[0\]\[0\] _00801_ _00802_ cpu.regs\[3\]\[0\] _00803_ _00805_ _00806_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07012_ _02505_ _02506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05497__I _01004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08387__A2 _03596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06398__A1 cpu.timer_capture\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08963_ _03768_ _04051_ _00430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07914_ _03220_ _03224_ _03225_ _00207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09336__B2 _04378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08894_ cpu.timer_div\[7\] _03972_ _03992_ _03988_ _03993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_98_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07845_ _01879_ _02714_ _03166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07776_ cpu.spi.counter\[3\] cpu.spi.counter\[2\] cpu.spi.counter\[4\] _03100_ _03104_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__09639__A2 cpu.ROM_addr_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09515_ _03077_ _00924_ _04550_ _04551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06727_ _02209_ _02210_ _02225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_65_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09446_ _04482_ _04483_ _04484_ _00480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06658_ _02152_ _02155_ _02156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07887__I _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05609_ _00675_ _01115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09377_ _04298_ _04411_ _04418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06589_ _02084_ _02085_ _02087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08328_ _03554_ _03547_ _03555_ _03541_ _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08075__A1 _03354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08259_ _03502_ _00275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_105_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07822__A1 cpu.timer_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06389__A1 _01881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10221_ _00160_ clknet_leaf_119_wb_clk_i cpu.regs\[6\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output78_I net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10152_ _00091_ clknet_leaf_2_wb_clk_i cpu.regs\[14\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10083_ _00026_ clknet_leaf_92_wb_clk_i cpu.base_address\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07127__I _02527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_22_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07290__C _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06864__A2 _01997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07813__B2 cpu.timer_div\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09010__C _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10419_ _00358_ clknet_leaf_15_wb_clk_i cpu.pwm_top\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_61_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07041__A2 _02516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05960_ _00863_ _00867_ _01330_ _01465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_05891_ _01202_ _01394_ _01395_ _01396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_49_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07630_ _02996_ _00152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05780__I _00874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07561_ cpu.regs\[10\]\[3\] _02949_ _02955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09300_ _04342_ _04343_ _03853_ _00475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06512_ _02007_ _02009_ _02011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06304__A1 cpu.PORTA_DDR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07492_ _01701_ _02904_ _02909_ _00101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09231_ _02795_ _01035_ _04275_ _04276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_8_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06443_ _01923_ _01940_ _01942_ _01943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09162_ _04042_ _04209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06374_ _01874_ _01875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08113_ _03335_ _03384_ _03388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05325_ _00586_ _00854_ _00855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09093_ _04150_ _04151_ _04152_ _00459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_102_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08044_ cpu.uart.div_counter\[12\] _03330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_05256_ _00699_ _00785_ _00786_ _00791_ _00008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_3_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05187_ cpu.uart.busy cpu.spi.busy _00724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07032__A2 _02516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09995_ _02493_ _04959_ _04960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08946_ _04033_ _04034_ _04035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08877_ _03128_ _03976_ _03979_ _03980_ _00415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_99_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07828_ _03147_ _03148_ cpu.timer\[9\] _03144_ _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_79_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07759_ cpu.PC\[11\] _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05623__C _00863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_106_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09429_ _04465_ _04466_ _04467_ _04468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08048__B2 _01881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08048__A1 _02824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10204_ _00143_ clknet_leaf_119_wb_clk_i cpu.regs\[8\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10135_ _00074_ clknet_leaf_108_wb_clk_i _00004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_89_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10066_ _01950_ cpu.regs\[15\]\[6\] _05011_ _05021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08523__A2 cpu.toggle_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09787__A1 net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05110_ _00647_ _00648_ _00649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_26_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06090_ _01558_ _01593_ _01594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05041_ cpu.regs\[4\]\[4\] cpu.regs\[5\]\[4\] cpu.regs\[6\]\[4\] cpu.regs\[7\]\[4\]
+ _00571_ _00575_ _00584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05708__C _01090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08800_ _03921_ _03922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09780_ cpu.ROM_spi_cycle\[2\] _04785_ _03122_ _04788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06992_ _02473_ _02485_ _02486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08731_ _03863_ _03864_ _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05943_ _01327_ _01445_ _01447_ _01448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08662_ _03801_ _03809_ _03810_ _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08514__A2 cpu.toggle_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07613_ _02983_ _02986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05874_ _01158_ _01379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08593_ _03759_ _03760_ _03761_ _03762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08278__B2 _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07544_ _02943_ cpu.regs\[11\]\[5\] _02933_ _02944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07475_ _01875_ cpu.regs\[14\]\[5\] _02890_ _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_9_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09214_ _00730_ _00784_ _04257_ _04259_ _03594_ _04260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_06426_ _01923_ _01925_ _01926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09145_ _00794_ _04184_ _04192_ _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06357_ _01739_ _00987_ _01755_ _01858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_17_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09076_ cpu.ROM_addr_buff\[0\] _04138_ _04139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07253__A2 _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08450__A1 cpu.orig_PC\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06288_ _01789_ cpu.regs\[9\]\[4\] _01702_ _01790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05103__I2 cpu.regs\[10\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05308_ _00833_ _00838_ _00580_ _00839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08027_ _02856_ cpu.uart.div_counter\[13\] cpu.uart.div_counter\[6\] _01881_ _03312_
+ _03313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_102_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05264__A1 _00793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05239_ _00773_ _00774_ _00775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_13_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09978_ _02049_ _02475_ _02469_ _04943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_89_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_89_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08929_ cpu.uart.divisor\[13\] _04013_ _04019_ _04020_ _04021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08929__C _04020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_18_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_18_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_99_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08505__A2 cpu.toggle_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06516__A1 _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_51_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07140__I _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05558__A2 _01059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10118_ _00061_ clknet_leaf_20_wb_clk_i cpu.timer_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10049_ _05010_ _00557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_59_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_11_Left_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05590_ _00675_ _00681_ _01096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_58_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07260_ _02721_ _02722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06211_ net43 _01510_ _01711_ _01712_ _01515_ _01713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_07191_ cpu.uart.divisor\[5\] _02651_ _02659_ _02662_ _02663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06142_ _01608_ _01172_ _01644_ _01258_ _01645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_41_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05246__A1 _00772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06073_ _01575_ _01576_ _01577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09901_ cpu.PORTB_DDR\[5\] _04876_ _04880_ _04881_ _04882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_1_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05024_ _00566_ _00567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09832_ _04014_ _04829_ _04830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09932__A1 cpu.PORTA_DDR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09763_ _02448_ _04722_ _04775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_67_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06975_ _02468_ _02469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08714_ _03178_ _03849_ _03837_ _03850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_4_9_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09694_ cpu.startup_cycle\[1\] _04718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07225__I _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05926_ _00721_ _01156_ _01093_ _01431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_107_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07171__A1 cpu.uart.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08645_ _01959_ _03778_ _03799_ _02744_ _00364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09160__A2 _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05857_ _01319_ _01358_ _01361_ _01362_ _01363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_77_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08576_ cpu.toggle_ctr\[11\] _03679_ _03748_ _03751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_05788_ _00914_ _01289_ _01293_ _01294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_07527_ _02065_ _01136_ _02932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_37_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07458_ _02887_ _00089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_107_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07389_ _02613_ _02821_ _02627_ _02822_ _00085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06409_ _01878_ _01908_ _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09128_ _01026_ _04177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_118_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09059_ _03997_ _04126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_102_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09923__A1 cpu.PORTA_DDR\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output60_I net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07135__I _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09206__A3 _01548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10598_ _00536_ clknet_leaf_70_wb_clk_i cpu.PORTB_DDR\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05228__A1 _00714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08193__A3 _03451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput90 net90 sram_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06760_ _02245_ _02257_ _02255_ _02258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05951__A2 _00919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05711_ _01216_ _01217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06691_ _02188_ _02171_ _02189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08430_ _03586_ _03633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05642_ _01147_ _01148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_93_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05573_ _01078_ _01048_ _01079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08361_ _03413_ _03583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_34_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08292_ cpu.uart.receive_div_counter\[4\] _03526_ _03527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_62_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07312_ _02748_ _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07243_ cpu.timer\[5\] _02707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07174_ _02647_ _02648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06125_ _01097_ _01628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06056_ _01346_ _01450_ _01560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09815_ _04815_ _04816_ _04817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06719__A1 _00820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06958_ _02451_ _02452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09746_ _02506_ _04745_ _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09677_ cpu.startup_cycle\[4\] _04703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_96_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09133__A2 _04180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05909_ _01413_ _01414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08628_ _03777_ _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07144__A1 _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06889_ _02379_ _02380_ _02386_ _02387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_68_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08559_ _03706_ _03736_ _03701_ _03740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08644__A1 _02722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10521_ _00459_ clknet_leaf_81_wb_clk_i cpu.last_addr\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10452_ _00391_ clknet_leaf_8_wb_clk_i cpu.timer\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10383_ _00322_ clknet_leaf_84_wb_clk_i cpu.orig_PC\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_33_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_33_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_20_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05069__S0 _00600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05873__I _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05933__A2 _00831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08883__A1 cpu.timer_div\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09013__C _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05449__A1 _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05113__I cpu.br_rel_dest\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06949__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07930_ _03237_ _01023_ _03238_ _03239_ _03240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_07861_ _03120_ _00703_ _03181_ _00198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07374__A1 _02810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07792_ _00789_ _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09600_ _04209_ _04622_ _04632_ _04327_ _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_39_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06812_ _00836_ _00927_ _02186_ _02263_ _02310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_09531_ _04544_ _04566_ _04484_ _00483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06743_ _02238_ _02240_ _02241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_104_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06674_ _02168_ _02169_ _02170_ _02171_ _02172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_19_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09462_ _04498_ _04499_ _04500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08413_ cpu.orig_PC\[2\] _03607_ _03621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09393_ _04432_ _04433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05625_ cpu.br_rel_dest\[0\] _01131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08344_ _02846_ _03520_ _03562_ _03569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05556_ _01061_ _01057_ _01062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08275_ _03495_ _03513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05487_ _00995_ _00996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_27_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07226_ _02692_ _02679_ _02693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07157_ _02633_ _02634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_4_1_0_wb_clk_i clknet_0_wb_clk_i clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_06108_ _01610_ _01611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05612__A1 _01052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07088_ _02574_ _02342_ _02575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06039_ _00997_ _01281_ _01542_ _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09354__A2 _04178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_12_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09729_ _04718_ _02043_ _02046_ _04746_ _04747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_97_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05868__I _01373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10504_ _00442_ clknet_leaf_79_wb_clk_i cpu.ROM_addr_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_80_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10435_ _00374_ clknet_leaf_10_wb_clk_i cpu.timer_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05851__B2 _01354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_51_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10366_ _00305_ clknet_leaf_90_wb_clk_i cpu.orig_flags\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10297_ _00236_ clknet_leaf_65_wb_clk_i cpu.spi.counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05410_ _00921_ _00922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08608__A1 _03573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06390_ cpu.uart.divisor\[14\] _01623_ _01890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05341_ cpu.PORTA_DDR\[7\] net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA_clkbuf_leaf_90_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08060_ _03345_ _00239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05272_ _00804_ _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_113_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07011_ _00668_ _02505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_70_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09033__A1 _03623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07595__A1 cpu.regs\[8\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08962_ _01098_ _04038_ _04048_ _04050_ _04051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07913_ cpu.spi.data_out_buff\[7\] _03113_ _03224_ _03225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08893_ _02775_ _03983_ _03992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_110_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07844_ _01879_ cpu.timer\[6\] cpu.timer\[5\] _01802_ _03165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XPHY_EDGE_ROW_3_Left_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07775_ _03097_ _03102_ _03103_ _02628_ _00190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08847__A1 cpu.spi.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06726_ _02222_ _02223_ _02224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09514_ _04526_ _04548_ _04549_ _04550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09445_ _00689_ _04484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06657_ _02153_ _02154_ _02155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05608_ _01110_ _01113_ _01114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_47_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07370__I1 _02078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09376_ _02562_ _00752_ _04416_ _04417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_46_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06588_ _02084_ _02085_ _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08327_ _03554_ _03548_ _03555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05688__I _00683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05539_ _01044_ _01045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08258_ cpu.uart.receive_buff\[4\] _03494_ _03498_ cpu.uart.receive_buff\[3\] _03502_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_62_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Left_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07209_ _02673_ _02678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08189_ _03345_ _03448_ _00259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10220_ _00159_ clknet_leaf_114_wb_clk_i cpu.regs\[6\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10151_ _00090_ clknet_leaf_2_wb_clk_i cpu.regs\[14\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10082_ _00025_ clknet_leaf_69_wb_clk_i net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XPHY_EDGE_ROW_58_Left_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05372__B _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07510__A1 cpu.regs\[12\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_67_Left_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_41_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06077__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09015__A1 _02531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10418_ _00357_ clknet_leaf_14_wb_clk_i cpu.pwm_top\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10349_ _00288_ clknet_leaf_37_wb_clk_i cpu.uart.receive_div_counter\[8\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07318__I _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_76_Left_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05039__S _00581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05890_ cpu.uart.divisor\[1\] _01202_ _01395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06001__A1 cpu.uart.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07560_ _02923_ _02950_ _02954_ _00124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06511_ _02007_ _02009_ _02010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07053__I _02541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08593__B _03761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09230_ cpu.PC\[0\] cpu.br_rel_dest\[0\] _04275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07491_ cpu.regs\[13\]\[3\] _02903_ _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05502__S _00885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06442_ _01471_ _01941_ _01942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09161_ _01429_ _01274_ _02668_ _04207_ _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_06373_ _01873_ _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_28_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08112_ _00793_ _03387_ _00243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09092_ cpu.last_addr\[3\] _04143_ _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06068__A1 _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05324_ cpu.regs\[12\]\[3\] cpu.regs\[13\]\[3\] cpu.regs\[14\]\[3\] cpu.regs\[15\]\[3\]
+ _00846_ _00847_ _00854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08043_ _02847_ _03325_ cpu.uart.div_counter\[13\] _02856_ _03328_ _03329_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_43_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05255_ _00790_ _00791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09006__A1 _01020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_112_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05186_ _00708_ _00722_ _00660_ _00723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_12_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09994_ _04950_ _04958_ _02448_ _04959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08945_ _00749_ _01704_ _00755_ _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__08517__B1 _01419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06791__A2 _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input22_I io_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08876_ _03346_ _03980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_98_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07827_ cpu.timer\[10\] _03148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07758_ _03086_ _03087_ _03088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07740__A1 _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06709_ _02205_ _02206_ _02207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07689_ _03007_ cpu.regs\[4\]\[4\] _03027_ _03034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_109_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09428_ _04465_ _04466_ _04298_ _04467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_81_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09359_ _04375_ _04384_ _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output90_I net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07559__A1 cpu.regs\[10\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10203_ _00142_ clknet_leaf_124_wb_clk_i cpu.regs\[8\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10134_ _00011_ clknet_leaf_86_wb_clk_i cpu.instr_cycle\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06231__A1 cpu.toggle_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10065_ _05020_ _00563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_46_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07731__A1 _00823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09484__A1 _03637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05830__B _01335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09787__A2 _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05040_ _00581_ _00583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_84_Left_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06222__A1 cpu.timer_div\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06991_ _02053_ _02483_ _02057_ _02484_ _02485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_08730_ cpu.timer_capture\[4\] _03858_ _03529_ _03864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05942_ _01326_ _01446_ _01447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08661_ cpu.timer_div_counter\[5\] _03807_ _03810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05873_ _01140_ _01378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07612_ _02984_ _02985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08592_ _00789_ _03761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XPHY_EDGE_ROW_93_Left_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07543_ _01873_ _02943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_118_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07474_ _02898_ _00094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09213_ _00729_ _04258_ _04259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09227__A1 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06425_ _01850_ _01852_ _01924_ _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09144_ _01025_ _04184_ _04191_ _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_44_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06356_ _01841_ _01774_ _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05031__I _00573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09075_ _04137_ _04138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06287_ _01788_ _01789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05307_ cpu.regs\[0\]\[2\] _00836_ _00837_ cpu.regs\[3\]\[2\] _00570_ _00574_ _00838_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_08026_ _02853_ _03310_ cpu.uart.div_counter\[5\] _01804_ _03312_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05238_ _00738_ _00741_ _00774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05103__I3 cpu.regs\[11\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05169_ cpu.br_rel_dest\[5\] _00706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09977_ net78 _04942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08928_ _03987_ _04020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08859_ cpu.spi.divisor\[5\] _03966_ _03968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_58_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_58_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_109_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_14_0_wb_clk_i clknet_0_wb_clk_i clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_10117_ _00060_ clknet_leaf_20_wb_clk_i cpu.timer_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10048_ _03223_ net69 _05009_ _05010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08201__B _03232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09016__C _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07704__A1 _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06210_ net55 _01211_ _01510_ _01712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_73_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09209__A1 _02327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07190_ _02661_ _02662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05494__A2 _00980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06141_ cpu.pwm_top\[3\] _01253_ _01642_ _01643_ _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_41_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06072_ _01316_ _01463_ _01576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09900_ _04846_ _04881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05023_ _00003_ _00566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_22_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09831_ _04813_ _04829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_67_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09762_ _04756_ _04773_ _04774_ _00506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06974_ _02053_ _02467_ _02468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07943__B2 _03247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08713_ _02690_ _02684_ _02675_ _03849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_05925_ _01133_ _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07506__I _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09696__A1 _03247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09693_ _04715_ _04716_ _02462_ _04717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_107_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08644_ _02722_ _03779_ _03799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09160__A3 _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05856_ _01320_ _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05026__I _00568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08765__C _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08575_ _03679_ _03748_ cpu.toggle_ctr\[11\] _03750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_1_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05787_ _00907_ _01292_ _01293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_77_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07526_ _02930_ _02919_ _02931_ _00113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_37_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07457_ _02880_ _02886_ _02887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_107_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07388_ _02610_ _02821_ _02625_ _02822_ _00084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06408_ _01018_ _01426_ _01791_ _01907_ _01908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_8_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09127_ _04166_ _04175_ _04176_ _00469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_leaf_105_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_105_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06339_ net94 _00616_ _01758_ _01840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_118_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08072__I _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09058_ cpu.regs\[3\]\[2\] _03641_ _04117_ _04125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06434__A1 _00656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08009_ _03297_ _03298_ _03299_ _03296_ _00228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_9_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08800__I _03921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output53_I net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10597_ _00535_ clknet_leaf_71_wb_clk_i cpu.PORTB_DDR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05228__A2 _00658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput80 net80 io_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput91 net91 sram_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_05710_ _00649_ _01107_ _01051_ _01216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06690_ _02187_ _02170_ _02188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05641_ _01146_ _01085_ _01095_ _01126_ _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_08360_ cpu.orig_IO_addr_buff\[0\] _03581_ _03582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_53_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05572_ _00676_ _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07311_ _02760_ _00069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_3_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_3_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_34_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08291_ _02841_ _03519_ _03526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_102_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07242_ _02706_ _00054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_33_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07173_ _00974_ _02647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06124_ cpu.uart.dout\[3\] _01522_ _01624_ _01626_ _01101_ _01627_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__05219__A2 _00754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06055_ _01558_ _01559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_112_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09814_ _04813_ _04816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_6_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07236__I _02673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09745_ _02452_ _04719_ _04761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06957_ cpu.startup_cycle\[3\] _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09676_ _04643_ _04701_ _04702_ _04231_ _00492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_69_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05908_ _01123_ _01413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06888_ cpu.PC\[5\] _02381_ _02385_ _02386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_96_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08627_ _03786_ _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09451__I _04408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05839_ _01343_ _01344_ _01345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_96_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08558_ cpu.toggle_ctr\[5\] cpu.toggle_ctr\[4\] cpu.toggle_ctr\[3\] _03733_ _03739_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_92_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08489_ cpu.toggle_top\[7\] _03666_ _03675_ _03671_ _03676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07509_ _01494_ _02921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_37_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10520_ _00458_ clknet_leaf_77_wb_clk_i cpu.last_addr\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_30_Left_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10451_ _00390_ clknet_leaf_25_wb_clk_i cpu.timer\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10382_ _00321_ clknet_leaf_84_wb_clk_i cpu.orig_PC\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_41_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05069__S1 _00601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_73_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_73_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_99_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09361__I _04194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06894__A1 _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09832__A1 _04014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_80_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05449__A2 _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06110__A3 _01243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09964__C _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09899__A1 _04018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07860_ _03122_ _03180_ cpu.needs_timer_interrupt _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07056__I _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07791_ _01709_ _03107_ _03115_ _00194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06811_ _00926_ _02186_ _02262_ _02309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_09530_ _04487_ _04562_ _04563_ _04565_ _04049_ _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__06895__I _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06742_ _00604_ _00928_ _02240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09271__I _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05505__S _00885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09461_ _04485_ _00866_ _04499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_104_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06673_ _00603_ _00954_ _02171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08412_ _02810_ _03619_ _03620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09392_ _02571_ _04410_ _04432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05304__I _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05624_ _00748_ _01033_ _01129_ _01130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_08343_ cpu.uart.receive_div_counter\[14\] _03567_ _03568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05555_ _00647_ _01060_ _01061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_58_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08274_ _03509_ _03512_ _03381_ _00280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_19_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07225_ _00957_ _02692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05486_ _00994_ _00995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07156_ _01199_ _02632_ _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__09051__A2 cpu.regs\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06107_ _01187_ _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07087_ _02036_ _02574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_112_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08350__I _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06038_ _01425_ _01542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_125_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07989_ cpu.uart.receive_buff\[0\] _03283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09728_ _04745_ _04746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09659_ _02537_ _04643_ _02484_ _04689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_8_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_120_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_120_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_53_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10503_ _00441_ clknet_leaf_97_wb_clk_i cpu.base_address\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10434_ _00373_ clknet_leaf_23_wb_clk_i cpu.timer_top\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05851__A2 _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06045__I _01548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10365_ _00304_ clknet_leaf_90_wb_clk_i cpu.orig_IO_addr_buff\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07585__B _02967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05884__I _01216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10296_ _00235_ clknet_leaf_66_wb_clk_i cpu.spi.counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05119__A1 _00656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05340_ cpu.PORTB_DDR\[7\] net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09281__A2 _04178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07292__A1 _02670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05271_ _00001_ _00804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07010_ _02471_ _02500_ _02503_ _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08792__A1 _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09266__I _04309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08961_ _04049_ _04050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07912_ _03105_ _03200_ _03223_ _00745_ _03224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_08892_ _03991_ _00419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_110_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07843_ _01802_ cpu.timer\[5\] cpu.timer\[4\] _01708_ _03163_ _03164_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_07774_ cpu.spi.dout\[0\] _03102_ _03103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06725_ _02184_ _02189_ _02223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09513_ _02376_ _00862_ _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09444_ _02588_ _04262_ _04483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06858__A1 _00638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06656_ _02138_ _02139_ _02154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05607_ _01112_ _01113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_74_Right_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_93_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09375_ _04387_ _04414_ _04415_ _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06587_ _00603_ _01015_ _02085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08326_ cpu.uart.receive_div_counter\[11\] _03554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08345__I _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05538_ _01043_ _01044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08257_ _03501_ _00274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_104_Left_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05469_ cpu.regs\[12\]\[4\] cpu.regs\[13\]\[4\] cpu.regs\[14\]\[4\] cpu.regs\[15\]\[4\]
+ _00871_ _00977_ _00978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_08188_ cpu.uart.counter\[2\] _03443_ _03447_ _03340_ _03448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07208_ _02676_ _02677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07139_ _02596_ _02539_ _02619_ _02511_ _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_30_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_83_Right_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_76_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07586__A2 _02967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10150_ _00089_ clknet_leaf_43_wb_clk_i cpu.uart.receive_counter\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08080__I _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10081_ _00024_ clknet_leaf_100_wb_clk_i cpu.regs\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05209__I _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07625__S _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_113_Left_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07424__I cpu.uart.divisor\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08838__A2 _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_92_Right_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07299__C _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07274__A1 _02732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06077__A2 _00919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10417_ _00356_ clknet_leaf_17_wb_clk_i cpu.pwm_counter\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10348_ _00287_ clknet_leaf_35_wb_clk_i cpu.uart.receive_div_counter\[7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05588__A1 _00721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10279_ _00218_ clknet_leaf_47_wb_clk_i cpu.spi.data_in_buff\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09814__I _04813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05760__A1 _00706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06510_ _01941_ _02008_ _02009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07490_ _01603_ _02904_ _02908_ _00100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06441_ _01915_ _01940_ _01941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_118_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_100_Right_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05789__I _01294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09160_ _00921_ _00945_ _01801_ _04206_ _04207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_16_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06372_ _01833_ _01872_ _01873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08111_ cpu.uart.div_counter\[3\] _03370_ _03386_ _03379_ _03387_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09091_ cpu.ROM_addr_buff\[3\] _04145_ _04151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05323_ _00848_ _00852_ _00581_ _00853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08042_ cpu.uart.div_counter\[4\] cpu.uart.divisor\[4\] _03328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05254_ _00789_ _00790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07017__A1 _00671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05185_ _00714_ _00721_ _00722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_12_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09993_ _04707_ _04953_ _04957_ _04958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05579__A1 _01053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07509__I _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08944_ _04032_ _04033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06240__A2 _01004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08875_ _02692_ _03973_ _03979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09190__A1 _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07244__I _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07826_ cpu.timer_top\[10\] _03147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input15_I io_in[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07757_ _02551_ _02352_ _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06708_ _00588_ _00954_ _02206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07688_ _02992_ _03028_ _03033_ _00173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09427_ _02587_ _02626_ _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06639_ _02081_ _02136_ _02137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09358_ _04347_ _04384_ _04399_ _04373_ _04400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_35_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08309_ _02826_ _03537_ _03540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07256__A1 cpu.timer_capture\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09289_ _00740_ _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_35_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10202_ _00141_ clknet_leaf_126_wb_clk_i cpu.regs\[8\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10133_ _00010_ clknet_leaf_88_wb_clk_i cpu.instr_cycle\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_89_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10064_ _01874_ cpu.regs\[15\]\[5\] _05011_ _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_46_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07103__B _02588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05558__B _01063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07329__I _02668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08747__A1 cpu.timer_capture\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06990_ _02058_ _02484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input7_I io_in[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05981__A1 _01484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05941_ _01327_ _01445_ _01446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08660_ cpu.timer_div_counter\[5\] _03807_ _03809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05872_ _01035_ _01377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_07611_ _02983_ _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08591_ cpu.pwm_counter\[1\] _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07542_ _02942_ _00118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_62_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07473_ _01789_ cpu.regs\[14\]\[4\] _02891_ _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_9_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09212_ _04256_ _04251_ _04255_ _04258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_63_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06424_ _01841_ _01017_ _01924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_84_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09143_ cpu.orig_flags\[2\] _04186_ _04190_ _04191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06355_ _01854_ _01855_ _01335_ _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_29_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05306_ cpu.regs\[2\]\[2\] _00837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09074_ _04136_ _04137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06286_ _01787_ _01788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08025_ cpu.uart.div_counter\[2\] _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05237_ _00710_ _00773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05168_ _00690_ _00705_ _00011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07410__A1 _02827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09976_ _04713_ _04941_ _00553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05099_ cpu.regs\[0\]\[7\] _00638_ cpu.regs\[2\]\[7\] cpu.regs\[3\]\[7\] _00633_
+ _00634_ _00639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08927_ _04018_ _04015_ _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08858_ _02653_ _03965_ _03967_ _00409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09163__A1 _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07809_ cpu.timer_div\[0\] _03127_ cpu.timer_div_counter\[2\] _03128_ _03129_ _03130_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_4_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05724__A1 cpu.timer_div\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08789_ _03911_ _03912_ _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_27_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_27_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_55_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08977__A1 _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10116_ _00059_ clknet_leaf_20_wb_clk_i cpu.timer_top\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10047_ _03238_ _03201_ _03812_ _05009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_59_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08708__I _03835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09457__A2 _01036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07612__I _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06140_ _01118_ _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06071_ _01377_ net91 _01575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09830_ _04813_ _04828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_67_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09761_ cpu.ROM_spi_dat_out\[5\] _04751_ _03761_ _04774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06973_ cpu.mem_cycle\[4\] _02467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08712_ cpu.timer_capture\[2\] _03841_ _03848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09145__A1 _00794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05924_ _01354_ _01429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09692_ cpu.startup_cycle\[1\] cpu.startup_cycle\[0\] _04716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_107_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08643_ _03798_ _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05855_ _00992_ _01359_ _01360_ _01361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08574_ _03729_ _03749_ _00343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_1_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05786_ _01290_ _01291_ _00886_ _01292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07525_ cpu.regs\[12\]\[7\] _02917_ _02931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_37_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07456_ _02521_ _02885_ cpu.uart.receive_counter\[3\] _02886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06131__A1 cpu.timer_div\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07387_ _02607_ _02821_ _02624_ _02822_ _00083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_45_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06407_ _01281_ _01295_ _01906_ _01542_ _01907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_20_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09126_ cpu.last_addr\[13\] _04142_ _04176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08959__A1 _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06338_ _01837_ _01838_ _01839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10066__I0 _01950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_31_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09057_ _04124_ _00451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06269_ _01554_ _01759_ _01771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08008_ cpu.uart.dout\[3\] _03294_ _03299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_103_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09959_ _02472_ _04640_ _02469_ _02470_ _04927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA_output46_I net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06122__A1 cpu.uart.divisor\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_70_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06048__I _01325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10596_ _00534_ clknet_leaf_71_wb_clk_i cpu.PORTB_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput70 net70 io_out[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__08178__A2 _03439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput81 net81 io_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput92 net92 sram_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07607__I _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05936__A1 _00831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_qcpu_99 io_oeb[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_37_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05640_ _01042_ _01146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06361__A1 _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05571_ cpu.IO_addr_buff\[2\] _01077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_4_13_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07310_ cpu.toggle_top\[11\] _02749_ _02759_ _02756_ _02760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08290_ _03510_ _03525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_85_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07861__A1 _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07241_ cpu.timer_capture\[4\] _02701_ _02705_ _02687_ _02706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_61_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10048__I0 _03223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07172_ _02646_ _00044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06123_ _01194_ _01625_ _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05475__I0 _00980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06054_ _01555_ _01557_ _01558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09218__B _03853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_115_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09813_ _01429_ _04815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_6_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05927__A1 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09744_ _04750_ _04760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06956_ cpu.startup_cycle\[5\] _02450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_118_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09675_ _02052_ _04695_ _04702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05907_ _01411_ _01234_ _01382_ _01412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06887_ _02382_ _02383_ _02384_ _02385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_96_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08626_ cpu.pwm_top\[2\] _03778_ _03785_ _03783_ _03786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05838_ _00891_ _00884_ _01344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07252__I _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08557_ _02521_ _03738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_81_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05769_ _00658_ _01030_ _01274_ _01275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08488_ _02775_ _03667_ _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07508_ _02914_ _02918_ _02920_ _00106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07439_ _00788_ _02871_ _02872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10450_ _00389_ clknet_leaf_25_wb_clk_i cpu.timer\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09109_ cpu.ROM_addr_buff\[8\] _04159_ _04164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10381_ _00320_ clknet_leaf_84_wb_clk_i cpu.orig_PC\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06407__A2 _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_92_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05656__B _01158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_42_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_42_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_99_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07162__I _02521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06894__A2 _02391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07843__A1 _01802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07843__B2 _01708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05410__I _00921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09596__A1 cpu.PC\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10579_ _00517_ clknet_leaf_69_wb_clk_i net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_51_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08721__I _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05472__I3 cpu.regs\[7\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07790_ cpu.spi.data_in_buff\[4\] _03108_ _03109_ _03115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06810_ _02306_ _02307_ _02308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_39_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06741_ _00919_ _02238_ _02239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09460_ _02377_ _01348_ _04498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_104_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08411_ _03586_ _03619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06334__A1 _00614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06672_ _00636_ _00893_ _01995_ _00801_ _02170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_80_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09391_ _04406_ _04431_ _04381_ _00478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_19_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05623_ _01035_ _01127_ _01128_ _00863_ _01129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_08342_ _02871_ _03566_ _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05554_ cpu.IO_addr_buff\[0\] _01060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08273_ _02834_ _03511_ _03512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05485_ _00993_ _00994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08117__B _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07224_ _02673_ _02691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07155_ _02631_ _02632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_42_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06106_ cpu.timer_top\[11\] _01609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_07086_ _02302_ _02341_ _02340_ _02322_ _02573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06037_ _01169_ _01537_ _01539_ _01268_ _01540_ _01541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_100_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06151__I _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07988_ _03282_ _00224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05990__I _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_114_Right_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09727_ cpu.startup_cycle\[6\] cpu.startup_cycle\[5\] cpu.startup_cycle\[4\] _04744_
+ _04745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_06939_ _02432_ _02434_ _02435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_97_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09658_ _02049_ _04686_ _04688_ _04231_ _00488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__06325__A1 cpu.toggle_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08609_ cpu.pwm_counter\[6\] _03772_ _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09589_ _04621_ _04622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06876__A2 _01156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10502_ _00440_ clknet_4_10_0_wb_clk_i cpu.base_address\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05230__I _00765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10433_ _00372_ clknet_leaf_28_wb_clk_i cpu.timer_div_counter\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10364_ _00303_ clknet_leaf_56_wb_clk_i cpu.orig_IO_addr_buff\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10295_ _00234_ clknet_leaf_63_wb_clk_i cpu.spi.counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07157__I _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06564__A1 _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07093__S _02567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05270_ _00000_ _00803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_12_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08960_ _02630_ _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07911_ _03221_ _03222_ _03223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08891_ cpu.timer_div\[6\] _03972_ _03990_ _03988_ _03991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_110_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07842_ cpu.timer_top\[4\] _02702_ _02696_ cpu.timer_top\[3\] _03162_ _03163_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07347__A3 _02541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09282__I _00761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07773_ _03101_ _03102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09512_ cpu.PC\[9\] _00862_ _04548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06307__A1 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06724_ _02219_ _02220_ _02221_ _02222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__05315__I _00845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09443_ _04293_ _04478_ _04481_ _04482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06858__A2 _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06655_ _02150_ _02151_ _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05606_ _00674_ _00679_ _01111_ _01112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09374_ cpu.PC\[4\] _00756_ _04415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08325_ _03552_ _03553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06586_ cpu.regs\[1\]\[6\] _02083_ _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05537_ cpu.instr_cycle\[2\] net25 _00661_ _00672_ _01043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_7_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08256_ cpu.uart.receive_buff\[3\] _03494_ _03498_ cpu.uart.receive_buff\[2\] _03501_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_105_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05468_ _00005_ _00977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08187_ cpu.uart.counter\[2\] _03342_ _03447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07207_ _01082_ _02676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_62_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07138_ _00696_ _02539_ _02619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08232__A1 _02657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05399_ _00897_ _00910_ _00911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_76_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06794__A1 _00918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07069_ _02338_ _02339_ _02557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_100_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10080_ _00023_ clknet_leaf_100_wb_clk_i cpu.regs\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_97_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09141__B _03853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10416_ _00355_ clknet_leaf_17_wb_clk_i cpu.pwm_counter\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09367__I _04407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10347_ _00286_ clknet_leaf_33_wb_clk_i cpu.uart.receive_div_counter\[6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10278_ _00217_ clknet_leaf_47_wb_clk_i cpu.spi.data_in_buff\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09023__I0 _00823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08526__A2 cpu.toggle_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09830__I _04813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06440_ _01837_ _01858_ _01924_ _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06371_ net31 _01368_ _01379_ _01871_ _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_29_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08110_ _03335_ _03384_ _03386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09090_ _03346_ _04150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_83_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08462__A1 _02636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05322_ cpu.regs\[0\]\[3\] _00850_ _00851_ cpu.regs\[3\]\[3\] _00846_ _00847_ _00852_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08041_ _02825_ _03324_ cpu.uart.div_counter\[8\] _02827_ _03326_ _03327_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_05253_ _00788_ _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05276__A1 _00002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09277__I _04309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08214__A1 _00922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05184_ _00715_ _00716_ _00720_ _00721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_110_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09992_ _04929_ _04956_ _04957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05579__A2 _01084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08943_ _01953_ _01155_ _00757_ _04032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__08517__A2 _01498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08874_ _03978_ _00414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_98_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05200__A1 _00733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07825_ _03144_ cpu.timer\[9\] cpu.timer\[8\] _03145_ _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07756_ _02351_ _02203_ _02350_ _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_79_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05751__A2 _01204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06707_ cpu.regs\[1\]\[6\] _00893_ _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09426_ _04436_ _04437_ _04464_ _04465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07687_ cpu.regs\[4\]\[3\] _03027_ _03033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07260__I _02721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06638_ _02114_ _02135_ _02136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09357_ _04391_ _04395_ _04398_ _04399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06569_ _01144_ _01164_ _02067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__10538__D _00476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08308_ _02832_ _03534_ _03539_ _03414_ _00287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_62_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09288_ _04294_ _04297_ _04329_ _04331_ _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08239_ _02669_ _03454_ _03489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10201_ _00140_ clknet_leaf_3_wb_clk_i cpu.regs\[8\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output76_I net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10132_ _00009_ clknet_leaf_88_wb_clk_i cpu.instr_cycle\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06767__B2 _00891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10062__S _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10063_ _05019_ _00562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07567__I0 _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06519__A1 _01451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06519__B2 _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08692__A1 _02670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09944__A1 _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05940_ _01437_ _01440_ _01444_ _01445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07183__A1 cpu.uart.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05871_ _01167_ _01374_ _01376_ _00013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08590_ _03759_ _00747_ _00349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07610_ _02932_ _02982_ _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_109_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07541_ _02941_ cpu.regs\[11\]\[4\] _02934_ _02942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_88_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07472_ _01701_ _02892_ _02897_ _00093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08109__C _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09211_ _04251_ _04255_ _04256_ _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_57_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06423_ _01915_ _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08904__I _04000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09142_ _00946_ _04186_ _04190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08435__A1 _02378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06354_ _01780_ _01851_ _01855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05305_ _00835_ _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09073_ _02047_ _04135_ _04136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_21_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06285_ _01492_ _01738_ _01785_ _01786_ _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_31_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08024_ cpu.uart.div_counter\[9\] _03310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_102_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05236_ _00771_ _00772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05167_ cpu.instr_cycle\[3\] _00699_ _00703_ _00704_ _00705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09935__A1 cpu.PORTA_DDR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10093__D _00036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09975_ net76 _04922_ _04924_ _04940_ _04941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_110_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05098_ _00637_ _00638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08926_ _02708_ _04018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08857_ cpu.spi.divisor\[4\] _03966_ _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07808_ cpu.timer_div\[0\] _03127_ _03125_ cpu.timer_div\[1\] _03129_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_79_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08788_ cpu.timer_capture\[14\] _03836_ _03897_ _03912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05280__S0 _00803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07739_ net12 _03054_ _02072_ _03071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_60_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08019__C _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09409_ _01877_ _04444_ _04447_ _04448_ _04449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_23_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_67_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_67_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_50_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08729__A2 _03811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05660__A1 _01137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07165__I cpu.uart.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10115_ _00058_ clknet_leaf_20_wb_clk_i cpu.timer_top\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10046_ _05008_ _00556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_59_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07640__A2 _03002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06070_ _01565_ _01574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09917__A1 cpu.PORTA_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_105_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09760_ cpu.ROM_spi_dat_out\[4\] _04732_ _04767_ _04773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06972_ cpu.mem_cycle\[0\] _02466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09691_ _02506_ _04715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08711_ _03847_ _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05923_ _01427_ _01428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05954__A2 _01452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07156__A1 _01199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08642_ cpu.pwm_top\[6\] _03787_ _03797_ _03795_ _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_107_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05854_ _01150_ _01151_ _01360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08573_ _03717_ _03748_ _03749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05785_ cpu.regs\[8\]\[7\] cpu.regs\[9\]\[7\] cpu.regs\[10\]\[7\] cpu.regs\[11\]\[7\]
+ _00961_ _01286_ _01291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_9_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07524_ _02032_ _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07459__A2 _01153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07455_ cpu.uart.receiving _02884_ _02885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_91_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06406_ _01276_ _01905_ _01906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08408__A1 _02797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07386_ _02595_ _02821_ _02623_ _02822_ _00082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_20_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05890__A1 cpu.uart.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09125_ cpu.ROM_addr_buff\[13\] _04154_ _04175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06337_ _01740_ _01750_ _01742_ _01838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_17_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_118_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09056_ _04123_ cpu.ROM_addr_buff\[9\] _04115_ _04124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06268_ _01554_ _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08007_ _03287_ _03298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05219_ _00659_ _00754_ _00755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_13_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06199_ _01166_ _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_9_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07395__B2 _02827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09958_ cpu.ROM_addr_buff\[12\] _02486_ _04925_ _04926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08909_ _03658_ _04002_ _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06103__B _01380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09889_ cpu.PORTB_DDR\[2\] _04865_ _04872_ _04870_ _04873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_99_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_114_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_114_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_99_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_56_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08809__I _03921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output39_I net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08647__A1 _03121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07870__A2 cpu.spi.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10595_ _00533_ clknet_leaf_71_wb_clk_i cpu.PORTB_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05881__A1 net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06830__B1 _00955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput60 net60 io_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput71 net71 io_out[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput82 net82 io_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput93 net93 sram_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05408__I _00919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05936__A2 _00918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07138__A1 _00696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10029_ _01993_ _04991_ _04992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_53_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05570_ _01075_ _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_53_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07240_ _02702_ _02703_ _02691_ _02704_ _02705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10048__I1 net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09994__B _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07171_ cpu.uart.divisor\[2\] _02634_ _02645_ _02639_ _02646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_26_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06122_ cpu.uart.divisor\[11\] _01623_ _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08810__A1 _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06053_ _01556_ _01557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09812_ _04813_ _04814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_6_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09743_ _04759_ _00502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06955_ cpu.startup_cycle\[6\] _02449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07129__A1 _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09674_ _04135_ _04645_ _04701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05906_ cpu.timer_capture\[9\] _01411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06886_ cpu.PC\[1\] _02384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_68_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08625_ _02754_ _03779_ _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05837_ _00876_ _00881_ _01343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_68_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08556_ _03727_ _03737_ _00337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_81_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05768_ _00706_ _00755_ _01274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07507_ cpu.regs\[12\]\[0\] _02919_ _02920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05699_ _01196_ _01048_ _01204_ _01205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_65_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08487_ _03674_ _00331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07301__A1 cpu.toggle_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07438_ _02870_ net15 _02871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_107_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05863__A1 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07369_ _01601_ _02780_ _02807_ _02808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09108_ _04162_ _04138_ _04163_ _03980_ _00463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_33_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10380_ _00319_ clknet_leaf_85_wb_clk_i cpu.orig_PC\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05615__A1 _01029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09039_ _00606_ _02563_ _04102_ _04111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05656__C _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08868__A1 _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_82_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_82_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_68_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09293__A1 _02078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_11_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_11_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_31_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10578_ _00516_ clknet_leaf_87_wb_clk_i net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09596__A2 _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09319__B _00776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05621__A4 _01126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10191__D _00130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07359__A1 _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06031__A1 cpu.timer_top\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08877__C _03980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06582__A2 _00955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08859__A1 cpu.spi.divisor\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06740_ _02236_ _02237_ _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_78_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06671_ _00636_ _01995_ _02169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08410_ _03617_ _03618_ _03610_ _00310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06334__A2 _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07382__I1 _02108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05622_ _01032_ _01128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09390_ _04346_ _04427_ _04430_ _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08341_ _02868_ _03565_ _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05553_ _00650_ _01058_ _01059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_59_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08272_ _03510_ _03511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_104_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05484_ _00970_ _00966_ _00914_ _00993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07223_ _02689_ _02690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_27_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07154_ _02630_ _00766_ _02631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09587__A2 _02391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06105_ cpu.toggle_top\[3\] _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_14_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07085_ _02571_ _02560_ _02572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_112_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06036_ _00930_ _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06022__A1 cpu.spi.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07987_ cpu.spi.data_in_buff\[7\] _03277_ _03278_ cpu.spi.data_in_buff\[6\] _03282_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09726_ _02463_ _04738_ _04739_ _02454_ _04743_ _04744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_06938_ _02169_ _02357_ _02433_ _02434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09657_ _04645_ _04687_ _04686_ _04688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06869_ _02353_ _02366_ _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08608_ _03573_ _03771_ _03772_ _00354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09588_ cpu.PC\[13\] _04620_ _04621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_38_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08539_ _03232_ _03724_ _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10501_ _00439_ clknet_leaf_97_wb_clk_i cpu.base_address\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05836__A1 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10432_ _00371_ clknet_leaf_28_wb_clk_i cpu.timer_div_counter\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10363_ _00302_ clknet_leaf_90_wb_clk_i cpu.orig_IO_addr_buff\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10294_ _00233_ clknet_leaf_48_wb_clk_i net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07761__A1 _03090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07173__I _00974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05827__A1 _01311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07910_ _03101_ _03199_ _03222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08890_ _02769_ _03983_ _03990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07841_ _03159_ _03160_ _03161_ _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06004__A1 net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07347__A4 _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07772_ _03098_ _03099_ cpu.spi.counter\[4\] _03100_ _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_09511_ _04546_ _04547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06723_ _02215_ _02218_ _02221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07083__I _02076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09442_ _04455_ _04463_ _04480_ _04339_ _04340_ _04481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06654_ _02150_ _02151_ _02152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05605_ _01067_ _01058_ _01111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09373_ cpu.PC\[4\] _00756_ _04414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06585_ _00985_ _02083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08324_ _00688_ _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_86_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05536_ _01039_ _01041_ _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_46_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08255_ _03500_ _00273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07967__B _00788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05467_ _00976_ net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09738__I _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08186_ _03446_ _00258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07206_ cpu.timer\[0\] _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_05398_ cpu.regs\[8\]\[1\] cpu.regs\[9\]\[1\] cpu.regs\[10\]\[1\] cpu.regs\[11\]\[1\]
+ _00899_ _00902_ _00910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07137_ _02613_ _02603_ _02616_ _02618_ _00037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_76_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_18_Left_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07068_ _02264_ _02544_ _02556_ _00030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06019_ _01504_ _01521_ _01522_ _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09709_ _03738_ _04729_ _04730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09496__A1 _00865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_27_Left_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07721__I _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05241__I _00776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10415_ _00354_ clknet_leaf_17_wb_clk_i cpu.pwm_counter\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_36_Left_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09420__A1 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06234__A1 _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10346_ _00285_ clknet_leaf_35_wb_clk_i cpu.uart.receive_div_counter\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10277_ _00216_ clknet_leaf_64_wb_clk_i cpu.spi.data_out_buff\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09023__I1 _02797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_45_Left_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05416__I _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_0_0_wb_clk_i clknet_0_wb_clk_i clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__09239__A1 _00751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07631__I _02031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05363__I3 cpu.regs\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05151__I _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06370_ _01599_ _01870_ _01871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05321_ cpu.regs\[2\]\[3\] _00851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_114_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05252_ _00787_ _00788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08040_ _02840_ cpu.uart.div_counter\[15\] _03325_ cpu.uart.divisor\[14\] _03326_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XPHY_EDGE_ROW_54_Left_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_11_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08214__A2 _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06225__A1 cpu.timer_capture\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05183_ _00718_ _00719_ _00720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_110_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09991_ _04951_ _04955_ _02463_ _04956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08942_ _00760_ _04031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05984__B1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06776__A2 _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08873_ cpu.timer_div\[1\] _03976_ _03977_ _03956_ _03978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_63_Left_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07824_ cpu.timer_top\[8\] _03145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09478__A1 _00802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07755_ _03085_ _00188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08637__I _02771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06706_ _02197_ _02198_ _02177_ _02204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_07686_ _02990_ _03028_ _03032_ _00172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_50_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09425_ _04438_ _04464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06637_ _02134_ _02135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_66_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09356_ _04324_ _04384_ _04396_ _04397_ _04398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06568_ _02065_ _01135_ _02066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08307_ cpu.uart.receive_div_counter\[7\] _03525_ _03538_ _03539_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05519_ _00726_ _01025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XPHY_EDGE_ROW_72_Left_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08453__A2 _03581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09287_ _04330_ _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06499_ net97 _01997_ _01998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08238_ _03488_ _00268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_62_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08169_ _03325_ _03426_ _03390_ _03427_ _03434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_10200_ _00139_ clknet_leaf_3_wb_clk_i cpu.regs\[8\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09953__A2 _00696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07964__A1 _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10131_ _00008_ clknet_leaf_87_wb_clk_i net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA_output69_I net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10062_ _01788_ cpu.regs\[15\]\[4\] _05012_ _05019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07716__A1 _02032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09931__I _03236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05236__I _00771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08444__A2 _03596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07404__B1 _02641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10329_ _00268_ clknet_leaf_54_wb_clk_i cpu.uart.data_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05855__B _01360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07707__A1 cpu.regs\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10052__I _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05870_ cpu.regs\[9\]\[0\] _01375_ _01376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_109_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07540_ _01788_ _02941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07471_ cpu.regs\[14\]\[3\] _02891_ _02897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09210_ _00739_ _04256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06422_ _01325_ _01921_ _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05041__S1 _00575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09141_ _04185_ _04189_ _03853_ _00470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_57_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06353_ _01835_ _01836_ _01854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_114_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09072_ _00694_ _04134_ _04135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08192__I _03450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05249__A2 _00783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05304_ _00834_ _00835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06446__A1 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06997__A2 _00733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08023_ net68 _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06284_ net30 _01368_ _01380_ _01786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_114_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08199__A1 _00728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05235_ _00770_ _00771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_102_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08920__I _04000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05166_ cpu.TIE cpu.needs_timer_interrupt _00704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_4_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07946__A1 _00975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09974_ _04938_ _04939_ _04930_ _04940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05421__A2 _00930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05097_ _00636_ _00637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09699__A1 _03227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08925_ _04017_ _00426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input20_I io_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08856_ _03958_ _03966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07807_ cpu.timer_div\[2\] _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__05185__A1 _00714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05999_ _01502_ _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08787_ _03908_ _03800_ _03833_ _03910_ _03881_ _03911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_07738_ _03064_ _03069_ _03070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05280__S1 _00573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07669_ _03007_ cpu.regs\[5\]\[4\] _03015_ _03022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_94_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09408_ _04309_ _04448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_23_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09339_ _04345_ _04380_ _04381_ _00476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_51_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_109_Right_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05660__A2 _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_36_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_36_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10114_ _00057_ clknet_leaf_29_wb_clk_i cpu.timer_capture\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10045_ _01299_ _04976_ _05007_ _04904_ _05008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08362__A1 _01074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07181__I _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06428__A1 _01479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09836__I _04683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06971_ _02456_ _02461_ _02464_ _02465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_09690_ _04074_ _04714_ _00494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08710_ cpu.timer_capture\[1\] _03843_ _03846_ _03795_ _03847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05922_ _00957_ _01282_ _01426_ _01427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08353__A1 _03573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08641_ _02769_ _03788_ _03797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05853_ _00862_ _01348_ _01359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_83_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08572_ _03732_ _03747_ _03748_ _00342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05784_ cpu.regs\[12\]\[7\] cpu.regs\[13\]\[7\] cpu.regs\[14\]\[7\] cpu.regs\[15\]\[7\]
+ _00961_ _01286_ _01290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07523_ _02929_ _00112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07454_ net15 _02884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06405_ _01168_ _01903_ _01904_ _01266_ _01707_ _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_91_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07385_ _02605_ _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06419__A1 _01437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09124_ _04166_ _04173_ _04174_ _00468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_60_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06336_ _01835_ _01836_ _01837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09055_ cpu.regs\[3\]\[1\] _03637_ _04117_ _04123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06267_ _01655_ _01668_ _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08006_ cpu.uart.receive_buff\[3\] _03297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_102_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05218_ cpu.br_rel_dest\[6\] _00754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06198_ _01700_ _01701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05149_ _00686_ _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09957_ _02469_ _02470_ _04644_ _04925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08908_ _04004_ _00422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09888_ _04823_ _04866_ _04872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08839_ cpu.timer\[15\] _03922_ _03953_ _03954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_56_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05514__I _00895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09844__A1 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10594_ _00532_ clknet_leaf_70_wb_clk_i net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_97_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06830__A1 _02078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06830__B2 _02327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput61 net61 io_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput50 net50 io_oeb[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput72 net72 io_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput94 net94 sram_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput83 net83 sram_addr[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10028_ _01998_ _02000_ _04991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09835__A1 _04018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07170_ _02644_ _02637_ _02645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06121_ _01612_ _01201_ _01621_ _01622_ _01623_ _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__07795__B _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06052_ _01550_ _00944_ _01556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_112_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09811_ _01087_ _04812_ _04813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09742_ cpu.ROM_spi_dat_out\[1\] _04756_ _04758_ _04684_ _04759_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06954_ _02447_ _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07129__A2 _02601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09673_ _04700_ _00491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05905_ _01405_ _01408_ _01409_ _01242_ _01410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_27_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06885_ cpu.PC\[2\] _02383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_96_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08624_ _03784_ _00358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05836_ net90 _00895_ _01341_ _01342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_89_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08555_ cpu.toggle_ctr\[4\] _03736_ _03737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05767_ _01169_ _01260_ _01264_ _01268_ _01272_ _01273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_TAPCELL_ROW_81_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07506_ _02916_ _02919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05698_ _01068_ _01050_ _01204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_65_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08486_ cpu.toggle_top\[6\] _03666_ _03673_ _03671_ _03674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07437_ _02866_ _02870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_13_0_wb_clk_i clknet_0_wb_clk_i clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_91_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07368_ _02547_ _02803_ _02806_ _02567_ _02807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_33_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09107_ cpu.ROM_addr_buff\[7\] _04154_ _04163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06319_ cpu.timer_capture\[5\] _01181_ _01817_ _01819_ _01240_ _01820_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_60_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09476__I _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07299_ _01261_ _02749_ _02751_ _02744_ _00066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06812__A1 _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09038_ _04110_ _00446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_60_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output51_I net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10646_ net49 net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06075__I _01465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_51_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_51_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10577_ _00515_ clknet_leaf_17_wb_clk_i net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_11_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08290__I _03510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07603__I0 _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05419__I _00929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06031__A2 _01175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_39_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06670_ _02167_ _00894_ _02168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_59_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05621_ _01042_ _01085_ _01095_ _01126_ _01127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_86_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09808__A1 _03738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08340_ cpu.uart.receive_div_counter\[14\] _03562_ _03565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05552_ _01057_ _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08465__I _00921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08271_ _02870_ _02884_ _03510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_74_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07295__A1 _01204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08492__B1 _01261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05483_ _00991_ _00992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_117_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07222_ cpu.timer\[2\] _02689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07153_ _01091_ _02630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06104_ cpu.TIE _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__09296__I _04194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09587__A3 _04408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07084_ _02380_ _02571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06035_ _01538_ _01263_ _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07986_ _03281_ _00223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09725_ _04741_ _04742_ _04743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06937_ _02356_ _02357_ _02169_ _02433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09656_ _04644_ _02597_ _04687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08607_ cpu.pwm_counter\[5\] _03769_ _03767_ _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06868_ _02363_ _02365_ _02366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09587_ _04597_ _02391_ _04408_ _04620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05533__A1 _01036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06799_ _02294_ _02296_ _02297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05819_ _01323_ _01324_ _01325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_65_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08538_ _03652_ _03723_ _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__08308__C _03414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08469_ _03661_ _00326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10500_ _00438_ clknet_leaf_97_wb_clk_i cpu.base_address\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05836__A2 _00895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10431_ _00370_ clknet_leaf_26_wb_clk_i cpu.timer_div_counter\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10362_ _00301_ clknet_leaf_90_wb_clk_i cpu.orig_IO_addr_buff\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10293_ _00232_ clknet_leaf_44_wb_clk_i cpu.uart.dout\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08710__A1 cpu.timer_capture\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05524__A1 _00714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07122__C _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05577__C _01082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08777__A1 cpu.timer_capture\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06533__I _02031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07565__S _02948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07201__A1 _02670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06004__A2 _00675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07840_ cpu.timer_top\[3\] _02696_ _02689_ cpu.timer_top\[2\] _03161_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_07771_ cpu.spi.counter\[0\] cpu.spi.counter\[1\] _03100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_75_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09510_ _03079_ _04349_ _04545_ _04546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06722_ _02205_ _02206_ _02220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_40_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09441_ _02418_ _04375_ _04479_ _04480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06653_ _02117_ _02118_ _02151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05604_ _01109_ _01110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_87_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09372_ _04278_ _04413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06584_ _00590_ _01996_ _02082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08323_ _03522_ _03551_ _00290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05535_ _00748_ _01040_ _01041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08254_ cpu.uart.receive_buff\[2\] _03494_ _03498_ cpu.uart.receive_buff\[1\] _03500_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05466_ _00949_ _00959_ _00975_ _00976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_62_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08185_ cpu.uart.counter\[1\] _03444_ _03445_ _02773_ _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07205_ _02673_ _02674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05397_ _00904_ _00908_ _00909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07136_ _02617_ _02618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_76_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07067_ _02544_ _02555_ _02556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06018_ _00684_ _01522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05059__I _00575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09708_ _04727_ _04711_ _04724_ _04729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07969_ _00788_ _03223_ _03271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_97_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05754__A1 _01170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09639_ cpu.last_addr\[1\] cpu.ROM_addr_buff\[1\] cpu.last_addr\[0\] _04671_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_87_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_41_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10414_ _00353_ clknet_leaf_17_wb_clk_i cpu.pwm_counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10345_ _00284_ clknet_leaf_34_wb_clk_i cpu.uart.receive_div_counter\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10276_ _00215_ clknet_leaf_58_wb_clk_i cpu.spi.data_out_buff\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_70_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05993__A1 _01161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09239__A2 _00761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06170__A1 _01454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_124_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08998__A1 _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05320_ _00849_ _00850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05251_ _00685_ _00787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_9_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05182_ cpu.base_address\[2\] _00719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__09411__A2 _04043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_7_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09990_ _02461_ _04954_ _04955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08941_ _04029_ _01449_ _04030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_86_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08872_ _03658_ _03973_ _03977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05607__I _01112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07823_ cpu.timer_top\[9\] _03144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07725__A2 _03057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07754_ _03084_ _00837_ _03052_ _03085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06705_ _02201_ _02202_ _02203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07685_ cpu.regs\[4\]\[2\] _03029_ _03032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09424_ _04462_ _04463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06636_ _02128_ _02133_ _02134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05342__I cpu.PORTA_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09355_ _04326_ _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06567_ _01130_ _02065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_117_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09749__I _04683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08306_ _03495_ _03537_ _03538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05518_ _01024_ net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09286_ _00739_ _03456_ _04330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06498_ _01996_ _01997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_90_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08237_ cpu.uart.data_buff\[7\] _03475_ _03487_ _03462_ _03488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_62_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05449_ _00925_ _00945_ _00958_ _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_43_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08168_ cpu.uart.div_counter\[14\] _03432_ _03433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08205__A3 _03451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_108_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_108_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08099_ _03376_ _03339_ _03377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07119_ _01304_ _02602_ _02604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_100_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10130_ _00073_ clknet_leaf_12_wb_clk_i cpu.toggle_top\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10061_ _01700_ _05013_ _05018_ _00561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08913__A1 _02754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07716__A2 _03041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05252__I _00787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07179__I _01005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10328_ _00267_ clknet_leaf_57_wb_clk_i cpu.uart.data_buff\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10259_ _00198_ clknet_leaf_60_wb_clk_i cpu.needs_timer_interrupt vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_0_Left_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08380__A2 _03596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05162__I net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07470_ _01603_ _02892_ _02896_ _00092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06421_ _01848_ _01920_ _01921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09140_ _00730_ _04177_ _04183_ _04188_ _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_57_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_6_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_6_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06352_ _01850_ _01852_ _01853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09071_ cpu.mem_cycle\[1\] _02050_ _04134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_72_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06283_ _01031_ _01784_ _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_05303_ cpu.regs\[1\]\[2\] _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_115_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08022_ _03307_ _03289_ _03308_ _03306_ _00232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_114_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05234_ _00710_ _00769_ _00712_ _00770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_12_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05165_ _00702_ net18 _00698_ _00703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_40_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09973_ cpu.ROM_addr_buff\[2\] _04927_ _02502_ cpu.ROM_addr_buff\[10\] _04939_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_73_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05096_ cpu.regs\[1\]\[7\] _00636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08924_ _02824_ _04013_ _04016_ _04006_ _04017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05501__S0 _00887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05337__I cpu.PORTA_DDR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08855_ _03958_ _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07806_ cpu.timer_div_counter\[0\] _03127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__06382__A1 cpu.PORTA_DDR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08786_ _03908_ _03909_ _03910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05185__A2 _00721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input13_I io_in[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05998_ _01197_ _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_79_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07552__I _02948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07737_ _02547_ _03065_ _03068_ _03069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_84_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07668_ _02992_ _03016_ _03021_ _00165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07882__A1 _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09407_ _04316_ _04432_ _04445_ _04446_ _04447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06619_ _02115_ _02116_ _02117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07599_ _02941_ cpu.regs\[8\]\[4\] _02969_ _02976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09338_ _00689_ _04381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_51_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07634__A1 _02071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09269_ _04268_ _04313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output81_I net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10113_ _00056_ clknet_leaf_29_wb_clk_i cpu.timer_capture\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09139__A1 _02647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05948__A1 _00991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_76_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_76_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10044_ _04378_ _04985_ _04990_ _05006_ _04976_ _05007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_59_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_3_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06676__A2 _00929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07130__C _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05651__A3 _00685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08050__A1 cpu.uart.divisor\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07637__I _02999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06970_ _02452_ _02462_ _02463_ _02464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input5_I io_in[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05921_ _01425_ _01426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08640_ _03796_ _00362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05852_ _00868_ _01330_ _01358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_83_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06364__A1 _01454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08571_ _03680_ _03715_ _03744_ _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_05783_ _01287_ _01288_ _00886_ _01289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06116__A1 net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07522_ _01951_ cpu.regs\[12\]\[6\] _02916_ _02929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07453_ _02880_ _02883_ _00088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06404_ cpu.toggle_top\[14\] _01262_ _01904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09123_ cpu.last_addr\[12\] _04142_ _04174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07384_ _02621_ _02821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06335_ _00615_ _01017_ _01836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08931__I _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09054_ _04122_ _00450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06266_ _01748_ _01767_ _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_32_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08005_ _03293_ _03288_ _03295_ _03296_ _00227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_103_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05217_ _00655_ _00658_ _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06451__I _01950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06197_ _01699_ _01700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08041__B2 _02827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05148_ _00685_ _00686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09956_ _04923_ _04921_ _04924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05079_ cpu.regs\[1\]\[6\] _00620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09887_ _04871_ _00534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08907_ cpu.uart.divisor\[8\] _04001_ _04003_ _03988_ _04004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08838_ _03923_ _02669_ _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_56_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08769_ _03894_ _03800_ _03866_ _03895_ _03881_ _03896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_56_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_123_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_123_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_118_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10593_ _00531_ clknet_leaf_68_wb_clk_i net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_97_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06830__A2 _00895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput51 net51 io_oeb[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput40 net40 io_oeb[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput62 net62 io_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput73 net73 io_out[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput84 net84 sram_addr[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput95 net95 sram_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_37_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09532__A1 _03090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10027_ _04292_ _04989_ _04990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06310__B _01200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05705__I _01210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_90_Left_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09847__I _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06120_ _01197_ _01623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08751__I _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06051_ _01550_ _00944_ _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_117_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_99_Right_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_94_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09810_ _01069_ _02746_ _04812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_10_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09741_ _04715_ _04707_ _04755_ _04757_ _04758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06953_ _02046_ _02447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_94_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05904_ cpu.timer_capture\[1\] _01236_ _01409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09523__A1 _04281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09672_ _03120_ _04699_ _04700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08198__I _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06884_ cpu.PC\[3\] _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08623_ cpu.pwm_top\[1\] _03778_ _03782_ _03783_ _03784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05835_ _01340_ _01341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08926__I _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08554_ cpu.toggle_ctr\[3\] _03733_ _03736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05766_ _01271_ _01272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_81_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07505_ _02917_ _02918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05697_ net6 _01203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08485_ _02769_ _03667_ _03673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07436_ _02868_ _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_92_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07367_ _02534_ _02334_ _02805_ _02576_ _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_33_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09106_ cpu.last_addr\[7\] _04162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06318_ _01180_ _01818_ _01819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09037_ _04109_ cpu.ROM_addr_buff\[4\] _04104_ _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07298_ _01023_ _02750_ _02751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07277__I _02735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06249_ _01744_ _01750_ _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09062__I0 cpu.regs\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09939_ _04909_ _00548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_99_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output44_I net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06500__A1 _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10645_ net49 net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_51_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10576_ _00514_ clknet_leaf_67_wb_clk_i net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_51_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06305__B _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05606__A3 _01111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_91_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_91_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07915__I _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_20_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_20_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06319__A1 cpu.timer_capture\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05435__I _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05790__A2 _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_30_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05620_ _01102_ _01106_ _01119_ _01125_ _01126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_80_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_19_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05551_ cpu.IO_addr_buff\[3\] cpu.IO_addr_buff\[2\] _01057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_59_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08270_ _02835_ _02869_ _03509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05170__I _00706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05482_ _00717_ _00991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07221_ _02688_ _00051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07152_ cpu.uart.divisor\[0\] _02629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08244__A1 _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06103_ _01605_ _01378_ _01380_ _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_112_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07083_ _02076_ _02570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_112_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06034_ cpu.toggle_top\[10\] _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_10_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07985_ cpu.spi.data_in_buff\[6\] _03277_ _03278_ cpu.spi.data_in_buff\[5\] _03281_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09724_ _02451_ _02462_ _04706_ _04742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06936_ _02430_ _02431_ _02432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05081__I1 _00621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09655_ _04642_ _04686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06867_ _02082_ _02097_ _02364_ _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_69_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08606_ _03769_ _03767_ cpu.pwm_counter\[5\] _03771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05818_ _01313_ _01324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09586_ _03649_ _04261_ _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06798_ _02290_ _02295_ _02296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_65_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05749_ _01171_ _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08537_ _03722_ _03723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_108_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08468_ cpu.toggle_top\[1\] _03654_ _03659_ _03660_ _03661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_49_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08483__A1 cpu.toggle_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07419_ cpu.uart.receive_div_counter\[6\] cpu.uart.divisor\[6\] _02852_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_18_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10430_ _00369_ clknet_leaf_27_wb_clk_i cpu.timer_div_counter\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08399_ _03606_ _03608_ _03610_ _00307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08391__I cpu.Z vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06904__I _02068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10361_ _00300_ clknet_leaf_104_wb_clk_i cpu.orig_IO_addr_buff\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10292_ _00231_ clknet_leaf_44_wb_clk_i cpu.uart.dout\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05221__A1 cpu.br_rel_dest\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05255__I _00790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07671__S _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05524__A2 _01029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_114_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10559_ _00497_ clknet_leaf_76_wb_clk_i cpu.startup_cycle\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_59_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10033__A1 _01992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07770_ cpu.spi.counter\[2\] _03099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06721_ _02215_ _02218_ _02219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09440_ _04335_ _04463_ _04479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08476__I _03653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06652_ _02147_ _02148_ _02149_ _02150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05603_ _01108_ _01109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_93_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09371_ _04411_ _04412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06583_ _00972_ _02079_ _02080_ _02081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_08322_ _02862_ _03547_ _03550_ _03541_ _03551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05534_ _00756_ _01040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08253_ _03499_ _00272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07204_ _01076_ _01099_ _01235_ _02631_ _02673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_74_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05465_ _00974_ _00975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_62_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08184_ _03441_ cpu.uart.counter\[1\] _03339_ _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_61_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05396_ _00905_ _00906_ _00907_ _00908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07135_ _00779_ _02617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07066_ _02545_ _02546_ _02554_ _02555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06017_ _01505_ _01520_ _01198_ _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_76_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07968_ _03269_ _03270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09707_ _04711_ _04724_ _04727_ _04728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06919_ _00621_ _02416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07899_ _03206_ _03213_ _03214_ _00203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09638_ _04140_ _04669_ _04670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05803__I _01157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09569_ _04298_ _04598_ _04603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08456__A1 _03354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10413_ _00352_ clknet_leaf_104_wb_clk_i cpu.pwm_counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10344_ _00283_ clknet_leaf_38_wb_clk_i cpu.uart.receive_div_counter\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10275_ _00214_ clknet_4_12_0_wb_clk_i cpu.spi.data_out_buff\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07195__A1 _02665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05745__A2 _01175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05250_ net18 _00699_ _00732_ _00786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05181_ _00717_ _00718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_110_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08940_ _04028_ _04029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08871_ _03971_ _03976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07822_ cpu.timer_top\[12\] _03141_ _03142_ cpu.timer_top\[11\] _03143_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05292__S0 _00568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07753_ _01601_ _02073_ _03083_ _03084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08686__A1 _02653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07684_ _02988_ _03028_ _03031_ _00171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06704_ _02140_ _02163_ _02202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07489__A2 _02905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07043__C _02522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09423_ _03614_ _02387_ _04461_ _02587_ _04462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_06635_ _02131_ _02132_ _02133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09354_ cpu.orig_PC\[4\] _04178_ _04396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08305_ _02832_ _03534_ _03537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_19_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06566_ _02062_ _02063_ _02064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05517_ _01020_ _01023_ _01024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_62_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09285_ _04311_ _04323_ _04328_ _04329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06497_ _01995_ _01996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08236_ _02664_ _03476_ _03486_ _03487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05448_ _00952_ _00957_ _00933_ _00958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07661__A2 _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08167_ _03402_ _03431_ _03432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07118_ _02602_ _02603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05379_ _00890_ _00886_ _00891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_30_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08098_ _03342_ _03343_ _03376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05424__A1 _00870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07049_ _02484_ _02537_ _02538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_11_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10060_ cpu.regs\[15\]\[3\] _05012_ _05018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09714__B _00689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08677__A1 _02732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05035__S0 _00572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08601__A1 _03573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10327_ _00266_ clknet_leaf_58_wb_clk_i cpu.uart.data_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10258_ _00197_ clknet_leaf_48_wb_clk_i cpu.spi.dout\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07168__A1 _02641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10189_ _00128_ clknet_leaf_120_wb_clk_i cpu.regs\[10\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_109_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06420_ _01437_ _01911_ _01919_ _01920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06351_ _01780_ _01851_ _01852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_29_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09070_ _04133_ _00455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_84_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06282_ _01739_ _01548_ _01768_ _01783_ _01784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_05302_ cpu.regs\[4\]\[2\] cpu.regs\[5\]\[2\] cpu.regs\[6\]\[2\] cpu.regs\[7\]\[2\]
+ _00570_ _00574_ _00833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_112_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08021_ cpu.uart.dout\[7\] _03287_ _03308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_71_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05233_ _00709_ _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05164_ _00701_ _00702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09972_ _04114_ _02501_ _04925_ _04938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05095_ cpu.regs\[4\]\[7\] cpu.regs\[5\]\[7\] cpu.regs\[6\]\[7\] cpu.regs\[7\]\[7\]
+ _00633_ _00634_ _00635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08923_ _04014_ _04015_ _04016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05501__S1 _00900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_110_Left_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07038__C _02522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08854_ _02648_ _03959_ _03964_ _00408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06906__A1 _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06906__B2 _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05997_ cpu.uart.dout\[2\] _00012_ _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07805_ cpu.timer_div_counter\[5\] _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08785_ _03904_ _03899_ _03909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_46_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07736_ _03066_ _03067_ _03068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07331__A1 cpu.toggle_top\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07667_ cpu.regs\[5\]\[3\] _03015_ _03021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08664__I _02660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09406_ _04269_ _04446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06618_ cpu.regs\[1\]\[3\] _01014_ _02116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07598_ _02925_ _02970_ _02975_ _00141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09084__A1 cpu.ROM_addr_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06549_ _02045_ _02046_ _02047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_63_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09337_ _04346_ _04374_ _04379_ _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_51_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09268_ _00762_ _04312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08219_ cpu.uart.data_buff\[3\] _03460_ _03473_ _03467_ _03474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08831__A1 cpu.timer_capture\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09199_ _02782_ _04244_ _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07398__A1 cpu.uart.divisor\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06912__I _02063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07398__B2 _02824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output74_I net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10112_ _00055_ clknet_leaf_29_wb_clk_i cpu.timer_capture\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05948__A2 _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10043_ _01552_ _04996_ _05001_ _05005_ _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_59_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_45_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_45_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_97_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07873__A2 cpu.spi.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05651__A4 _01091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05920_ _01133_ _01094_ _01425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05851_ _01346_ _01350_ _01353_ _01354_ _01356_ _01357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_83_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08570_ _03715_ _03744_ _03680_ _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10012__C _03347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07521_ _02928_ _00111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05782_ cpu.regs\[0\]\[7\] cpu.regs\[1\]\[7\] cpu.regs\[2\]\[7\] cpu.regs\[3\]\[7\]
+ _00898_ _01286_ _01288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_88_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07452_ _02873_ _02882_ cpu.uart.receive_counter\[2\] _02883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06403_ cpu.toggle_top\[6\] _01643_ _01902_ _01257_ _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_45_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07383_ _02820_ _00081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09122_ cpu.ROM_addr_buff\[12\] _04154_ _04173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06334_ _00614_ _01706_ _01835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_29_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09053_ _04121_ cpu.ROM_addr_buff\[8\] _04115_ _04122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06265_ _01360_ _01751_ _01754_ _01756_ _01766_ _01767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_32_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08004_ _02617_ _03296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_102_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05216_ _00708_ _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_13_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06196_ _01606_ _01653_ _01698_ _01492_ _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_05147_ _00651_ _00685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_40_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09955_ _02465_ _04923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_110_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05078_ cpu.regs\[4\]\[6\] cpu.regs\[5\]\[6\] cpu.regs\[6\]\[6\] cpu.regs\[7\]\[6\]
+ _00617_ _00618_ _00619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09886_ cpu.PORTB_DDR\[1\] _04865_ _04869_ _04870_ _04871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08906_ _02636_ _04002_ _04003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08837_ _03952_ _00403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_56_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08768_ _03894_ _03890_ _03895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08699_ _03831_ _03837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07304__A1 _02754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_0_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07719_ _02574_ _02409_ _02072_ _03051_ _03052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_94_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05811__I cpu.br_rel_dest\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10592_ _00530_ clknet_leaf_68_wb_clk_i net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_106_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05258__I _00792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput52 net52 io_oeb[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput41 net41 io_oeb[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput63 net63 io_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput74 net74 io_out[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_101_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput85 net85 sram_addr[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput96 net96 sram_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10026_ _00865_ _04985_ _04988_ _04196_ _04989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_clkbuf_leaf_20_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09599__A2 _04033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06050_ _01553_ _01554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_117_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09863__I _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09740_ cpu.ROM_spi_dat_out\[0\] _04731_ _04757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06952_ _02446_ _00024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
.ends

