magic
tech gf180mcuD
magscale 1 10
timestamp 1753967993
<< metal1 >>
rect 1344 20410 22784 20444
rect 1344 20358 6534 20410
rect 6586 20358 6638 20410
rect 6690 20358 6742 20410
rect 6794 20358 11854 20410
rect 11906 20358 11958 20410
rect 12010 20358 12062 20410
rect 12114 20358 17174 20410
rect 17226 20358 17278 20410
rect 17330 20358 17382 20410
rect 17434 20358 22494 20410
rect 22546 20358 22598 20410
rect 22650 20358 22702 20410
rect 22754 20358 22784 20410
rect 1344 20324 22784 20358
rect 2158 20130 2210 20142
rect 2158 20066 2210 20078
rect 4510 20130 4562 20142
rect 4510 20066 4562 20078
rect 6750 20130 6802 20142
rect 6750 20066 6802 20078
rect 9550 20130 9602 20142
rect 9550 20066 9602 20078
rect 11230 20130 11282 20142
rect 11230 20066 11282 20078
rect 13358 20130 13410 20142
rect 13358 20066 13410 20078
rect 15710 20130 15762 20142
rect 15710 20066 15762 20078
rect 17950 20130 18002 20142
rect 17950 20066 18002 20078
rect 20078 20130 20130 20142
rect 20078 20066 20130 20078
rect 20974 20130 21026 20142
rect 20974 20066 21026 20078
rect 22094 20130 22146 20142
rect 22094 20066 22146 20078
rect 2494 20018 2546 20030
rect 2494 19954 2546 19966
rect 4174 20018 4226 20030
rect 4174 19954 4226 19966
rect 6414 20018 6466 20030
rect 6414 19954 6466 19966
rect 9214 20018 9266 20030
rect 9214 19954 9266 19966
rect 10894 20018 10946 20030
rect 10894 19954 10946 19966
rect 13694 20018 13746 20030
rect 13694 19954 13746 19966
rect 15374 20018 15426 20030
rect 15374 19954 15426 19966
rect 17614 20018 17666 20030
rect 17614 19954 17666 19966
rect 19742 20018 19794 20030
rect 19742 19954 19794 19966
rect 20638 20018 20690 20030
rect 20638 19954 20690 19966
rect 21758 20018 21810 20030
rect 21758 19954 21810 19966
rect 1344 19626 22624 19660
rect 1344 19574 3874 19626
rect 3926 19574 3978 19626
rect 4030 19574 4082 19626
rect 4134 19574 9194 19626
rect 9246 19574 9298 19626
rect 9350 19574 9402 19626
rect 9454 19574 14514 19626
rect 14566 19574 14618 19626
rect 14670 19574 14722 19626
rect 14774 19574 19834 19626
rect 19886 19574 19938 19626
rect 19990 19574 20042 19626
rect 20094 19574 22624 19626
rect 1344 19540 22624 19574
rect 3054 19458 3106 19470
rect 3054 19394 3106 19406
rect 3726 19458 3778 19470
rect 3726 19394 3778 19406
rect 4510 19458 4562 19470
rect 4510 19394 4562 19406
rect 5854 19458 5906 19470
rect 5854 19394 5906 19406
rect 10894 19458 10946 19470
rect 10894 19394 10946 19406
rect 15150 19458 15202 19470
rect 14242 19350 14254 19402
rect 14306 19350 14318 19402
rect 15150 19394 15202 19406
rect 16382 19458 16434 19470
rect 16382 19394 16434 19406
rect 18622 19458 18674 19470
rect 18622 19394 18674 19406
rect 21534 19458 21586 19470
rect 21534 19394 21586 19406
rect 3390 19234 3442 19246
rect 3390 19170 3442 19182
rect 4062 19234 4114 19246
rect 4062 19170 4114 19182
rect 4174 19234 4226 19246
rect 5518 19234 5570 19246
rect 5170 19182 5182 19234
rect 5234 19182 5246 19234
rect 4174 19170 4226 19182
rect 5518 19170 5570 19182
rect 7982 19234 8034 19246
rect 9102 19234 9154 19246
rect 8642 19182 8654 19234
rect 8706 19182 8718 19234
rect 7982 19170 8034 19182
rect 9102 19170 9154 19182
rect 11230 19234 11282 19246
rect 14814 19234 14866 19246
rect 14130 19182 14142 19234
rect 14194 19182 14206 19234
rect 14466 19182 14478 19234
rect 14530 19182 14542 19234
rect 11230 19170 11282 19182
rect 14814 19170 14866 19182
rect 16046 19234 16098 19246
rect 16046 19170 16098 19182
rect 18286 19234 18338 19246
rect 18286 19170 18338 19182
rect 19070 19234 19122 19246
rect 20078 19234 20130 19246
rect 19730 19182 19742 19234
rect 19794 19182 19806 19234
rect 19070 19170 19122 19182
rect 20078 19170 20130 19182
rect 21198 19234 21250 19246
rect 21198 19170 21250 19182
rect 5014 19066 5066 19078
rect 8530 19014 8542 19066
rect 8594 19014 8606 19066
rect 5014 19002 5066 19014
rect 9438 19010 9490 19022
rect 9438 18946 9490 18958
rect 15766 19010 15818 19022
rect 19506 19014 19518 19066
rect 19570 19014 19582 19066
rect 15766 18946 15818 18958
rect 20414 19010 20466 19022
rect 20414 18946 20466 18958
rect 1344 18842 22784 18876
rect 1344 18790 6534 18842
rect 6586 18790 6638 18842
rect 6690 18790 6742 18842
rect 6794 18790 11854 18842
rect 11906 18790 11958 18842
rect 12010 18790 12062 18842
rect 12114 18790 17174 18842
rect 17226 18790 17278 18842
rect 17330 18790 17382 18842
rect 17434 18790 22494 18842
rect 22546 18790 22598 18842
rect 22650 18790 22702 18842
rect 22754 18790 22784 18842
rect 1344 18756 22784 18790
rect 11006 18674 11058 18686
rect 8866 18566 8878 18618
rect 8930 18566 8942 18618
rect 11006 18610 11058 18622
rect 15038 18674 15090 18686
rect 15038 18610 15090 18622
rect 14410 18510 14422 18562
rect 14474 18510 14486 18562
rect 20122 18510 20134 18562
rect 20186 18510 20198 18562
rect 7410 18398 7422 18450
rect 7474 18398 7486 18450
rect 7634 18413 7646 18465
rect 7698 18413 7710 18465
rect 8530 18454 8542 18506
rect 8594 18454 8606 18506
rect 8766 18450 8818 18462
rect 8082 18398 8094 18450
rect 8146 18398 8158 18450
rect 9650 18413 9662 18465
rect 9714 18413 9726 18465
rect 10670 18450 10722 18462
rect 9986 18398 9998 18450
rect 10050 18398 10062 18450
rect 8766 18386 8818 18398
rect 10670 18386 10722 18398
rect 14030 18450 14082 18462
rect 14030 18386 14082 18398
rect 14142 18450 14194 18462
rect 14142 18386 14194 18398
rect 14702 18450 14754 18462
rect 14702 18386 14754 18398
rect 17838 18450 17890 18462
rect 17838 18386 17890 18398
rect 18174 18450 18226 18462
rect 18174 18386 18226 18398
rect 19294 18450 19346 18462
rect 19294 18386 19346 18398
rect 19630 18450 19682 18462
rect 19630 18386 19682 18398
rect 19854 18450 19906 18462
rect 20862 18450 20914 18462
rect 20570 18398 20582 18450
rect 20634 18398 20646 18450
rect 19854 18386 19906 18398
rect 20862 18386 20914 18398
rect 20974 18450 21026 18462
rect 20974 18386 21026 18398
rect 21590 18450 21642 18462
rect 21590 18386 21642 18398
rect 22318 18450 22370 18462
rect 22318 18386 22370 18398
rect 3558 18338 3610 18350
rect 18958 18338 19010 18350
rect 7746 18286 7758 18338
rect 7810 18286 7822 18338
rect 9538 18286 9550 18338
rect 9602 18286 9614 18338
rect 3558 18274 3610 18286
rect 18958 18274 19010 18286
rect 21982 18226 22034 18238
rect 21982 18162 22034 18174
rect 1344 18058 22624 18092
rect 1344 18006 3874 18058
rect 3926 18006 3978 18058
rect 4030 18006 4082 18058
rect 4134 18006 9194 18058
rect 9246 18006 9298 18058
rect 9350 18006 9402 18058
rect 9454 18006 14514 18058
rect 14566 18006 14618 18058
rect 14670 18006 14722 18058
rect 14774 18006 19834 18058
rect 19886 18006 19938 18058
rect 19990 18006 20042 18058
rect 20094 18006 22624 18058
rect 1344 17972 22624 18006
rect 8318 17890 8370 17902
rect 3502 17834 3554 17846
rect 8318 17826 8370 17838
rect 9382 17834 9434 17846
rect 13850 17838 13862 17890
rect 13914 17838 13926 17890
rect 14634 17838 14646 17890
rect 14698 17838 14710 17890
rect 3502 17770 3554 17782
rect 4510 17778 4562 17790
rect 9382 17770 9434 17782
rect 4510 17714 4562 17726
rect 8710 17666 8762 17678
rect 8990 17666 9042 17678
rect 13358 17666 13410 17678
rect 2702 17576 2714 17628
rect 2766 17576 2778 17628
rect 3378 17614 3390 17666
rect 3442 17614 3454 17666
rect 3950 17628 4002 17640
rect 4274 17614 4286 17666
rect 4338 17614 4350 17666
rect 3950 17564 4002 17576
rect 4678 17610 4730 17622
rect 8866 17614 8878 17666
rect 8930 17614 8942 17666
rect 9538 17614 9550 17666
rect 9602 17614 9614 17666
rect 8710 17602 8762 17614
rect 8990 17602 9042 17614
rect 13358 17602 13410 17614
rect 13582 17666 13634 17678
rect 13582 17602 13634 17614
rect 14254 17666 14306 17678
rect 14254 17602 14306 17614
rect 14366 17666 14418 17678
rect 14366 17602 14418 17614
rect 4678 17546 4730 17558
rect 11510 17442 11562 17454
rect 11510 17378 11562 17390
rect 12966 17442 13018 17454
rect 12966 17378 13018 17390
rect 1344 17274 22784 17308
rect 1344 17222 6534 17274
rect 6586 17222 6638 17274
rect 6690 17222 6742 17274
rect 6794 17222 11854 17274
rect 11906 17222 11958 17274
rect 12010 17222 12062 17274
rect 12114 17222 17174 17274
rect 17226 17222 17278 17274
rect 17330 17222 17382 17274
rect 17434 17222 22494 17274
rect 22546 17222 22598 17274
rect 22650 17222 22702 17274
rect 22754 17222 22784 17274
rect 1344 17188 22784 17222
rect 8486 17106 8538 17118
rect 8486 17042 8538 17054
rect 13134 16994 13186 17006
rect 10826 16942 10838 16994
rect 10890 16942 10902 16994
rect 3166 16882 3218 16894
rect 3726 16882 3778 16894
rect 3434 16830 3446 16882
rect 3498 16830 3510 16882
rect 3166 16818 3218 16830
rect 3726 16818 3778 16830
rect 3950 16882 4002 16894
rect 3950 16818 4002 16830
rect 4174 16882 4226 16894
rect 11118 16882 11170 16894
rect 4834 16830 4846 16882
rect 4898 16830 4910 16882
rect 7634 16830 7646 16882
rect 7698 16830 7710 16882
rect 7970 16830 7982 16882
rect 8034 16830 8046 16882
rect 4174 16818 4226 16830
rect 11118 16818 11170 16830
rect 11342 16882 11394 16894
rect 12002 16863 12014 16915
rect 12066 16863 12078 16915
rect 12226 16886 12238 16938
rect 12290 16886 12302 16938
rect 13134 16930 13186 16942
rect 21590 16994 21642 17006
rect 21590 16930 21642 16942
rect 12674 16863 12686 16915
rect 12738 16863 12750 16915
rect 12984 16863 12996 16915
rect 13048 16863 13060 16915
rect 18286 16882 18338 16894
rect 11342 16818 11394 16830
rect 18286 16818 18338 16830
rect 21982 16882 22034 16894
rect 21982 16818 22034 16830
rect 22318 16882 22370 16894
rect 22318 16818 22370 16830
rect 7534 16714 7586 16726
rect 2830 16658 2882 16670
rect 4946 16662 4958 16714
rect 5010 16662 5022 16714
rect 7534 16650 7586 16662
rect 18622 16658 18674 16670
rect 2830 16594 2882 16606
rect 18622 16594 18674 16606
rect 1344 16490 22624 16524
rect 1344 16438 3874 16490
rect 3926 16438 3978 16490
rect 4030 16438 4082 16490
rect 4134 16438 9194 16490
rect 9246 16438 9298 16490
rect 9350 16438 9402 16490
rect 9454 16438 14514 16490
rect 14566 16438 14618 16490
rect 14670 16438 14722 16490
rect 14774 16438 19834 16490
rect 19886 16438 19938 16490
rect 19990 16438 20042 16490
rect 20094 16438 22624 16490
rect 1344 16404 22624 16438
rect 4286 16266 4338 16278
rect 18218 16270 18230 16322
rect 18282 16270 18294 16322
rect 19338 16270 19350 16322
rect 19402 16270 19414 16322
rect 3154 16214 3166 16266
rect 3218 16214 3230 16266
rect 4286 16202 4338 16214
rect 11622 16210 11674 16222
rect 11622 16146 11674 16158
rect 3950 16098 4002 16110
rect 14926 16098 14978 16110
rect 3378 16046 3390 16098
rect 3442 16046 3454 16098
rect 4386 16046 4398 16098
rect 4450 16046 4462 16098
rect 4610 16046 4622 16098
rect 4674 16046 4686 16098
rect 14242 16046 14254 16098
rect 14306 16046 14318 16098
rect 3950 16034 4002 16046
rect 14690 15990 14702 16042
rect 14754 15990 14766 16042
rect 14926 16034 14978 16046
rect 15374 16098 15426 16110
rect 15374 16034 15426 16046
rect 18510 16098 18562 16110
rect 18510 16034 18562 16046
rect 18734 16098 18786 16110
rect 18734 16034 18786 16046
rect 18846 16098 18898 16110
rect 18846 16034 18898 16046
rect 19070 16098 19122 16110
rect 19070 16034 19122 16046
rect 15026 15878 15038 15930
rect 15090 15878 15102 15930
rect 15710 15874 15762 15886
rect 15710 15810 15762 15822
rect 1344 15706 22784 15740
rect 1344 15654 6534 15706
rect 6586 15654 6638 15706
rect 6690 15654 6742 15706
rect 6794 15654 11854 15706
rect 11906 15654 11958 15706
rect 12010 15654 12062 15706
rect 12114 15654 17174 15706
rect 17226 15654 17278 15706
rect 17330 15654 17382 15706
rect 17434 15654 22494 15706
rect 22546 15654 22598 15706
rect 22650 15654 22702 15706
rect 22754 15654 22784 15706
rect 1344 15620 22784 15654
rect 3602 15430 3614 15482
rect 3666 15430 3678 15482
rect 12674 15430 12686 15482
rect 12738 15430 12750 15482
rect 19170 15430 19182 15482
rect 19234 15430 19246 15482
rect 20402 15430 20414 15482
rect 20466 15430 20478 15482
rect 3490 15262 3502 15314
rect 3554 15262 3566 15314
rect 3826 15306 3838 15358
rect 3890 15306 3902 15358
rect 12574 15353 12626 15365
rect 12226 15262 12238 15314
rect 12290 15262 12302 15314
rect 12574 15289 12626 15301
rect 12798 15314 12850 15326
rect 14914 15277 14926 15329
rect 14978 15277 14990 15329
rect 15250 15262 15262 15314
rect 15314 15262 15326 15314
rect 18274 15262 18286 15314
rect 18338 15262 18350 15314
rect 18498 15306 18510 15358
rect 18562 15306 18574 15358
rect 19058 15262 19070 15314
rect 19122 15262 19134 15314
rect 19394 15277 19406 15329
rect 19458 15277 19470 15329
rect 20526 15314 20578 15326
rect 20906 15318 20918 15370
rect 20970 15318 20982 15370
rect 21186 15262 21198 15314
rect 21250 15262 21262 15314
rect 12798 15250 12850 15262
rect 20526 15250 20578 15262
rect 14802 15150 14814 15202
rect 14866 15150 14878 15202
rect 18610 15150 18622 15202
rect 18674 15150 18686 15202
rect 1344 14922 22624 14956
rect 1344 14870 3874 14922
rect 3926 14870 3978 14922
rect 4030 14870 4082 14922
rect 4134 14870 9194 14922
rect 9246 14870 9298 14922
rect 9350 14870 9402 14922
rect 9454 14870 14514 14922
rect 14566 14870 14618 14922
rect 14670 14870 14722 14922
rect 14774 14870 19834 14922
rect 19886 14870 19938 14922
rect 19990 14870 20042 14922
rect 20094 14870 22624 14922
rect 1344 14836 22624 14870
rect 4666 14702 4678 14754
rect 4730 14702 4742 14754
rect 5798 14642 5850 14654
rect 5798 14578 5850 14590
rect 4958 14530 5010 14542
rect 4958 14466 5010 14478
rect 5182 14530 5234 14542
rect 5182 14466 5234 14478
rect 8654 14530 8706 14542
rect 8654 14466 8706 14478
rect 13806 14530 13858 14542
rect 13806 14466 13858 14478
rect 14030 14530 14082 14542
rect 14030 14466 14082 14478
rect 21198 14530 21250 14542
rect 21198 14466 21250 14478
rect 13514 14366 13526 14418
rect 13578 14366 13590 14418
rect 8318 14306 8370 14318
rect 21534 14306 21586 14318
rect 8978 14254 8990 14306
rect 9042 14303 9054 14306
rect 9762 14303 9774 14306
rect 9042 14257 9774 14303
rect 9042 14254 9054 14257
rect 9762 14254 9774 14257
rect 9826 14254 9838 14306
rect 8318 14242 8370 14254
rect 21534 14242 21586 14254
rect 1344 14138 22784 14172
rect 1344 14086 6534 14138
rect 6586 14086 6638 14138
rect 6690 14086 6742 14138
rect 6794 14086 11854 14138
rect 11906 14086 11958 14138
rect 12010 14086 12062 14138
rect 12114 14086 17174 14138
rect 17226 14086 17278 14138
rect 17330 14086 17382 14138
rect 17434 14086 22494 14138
rect 22546 14086 22598 14138
rect 22650 14086 22702 14138
rect 22754 14086 22784 14138
rect 1344 14052 22784 14086
rect 5686 13970 5738 13982
rect 5686 13906 5738 13918
rect 9774 13970 9826 13982
rect 4174 13858 4226 13870
rect 8866 13862 8878 13914
rect 8930 13862 8942 13914
rect 9774 13906 9826 13918
rect 11778 13862 11790 13914
rect 11842 13862 11854 13914
rect 20514 13862 20526 13914
rect 20578 13862 20590 13914
rect 4174 13794 4226 13806
rect 4510 13746 4562 13758
rect 4510 13682 4562 13694
rect 4622 13746 4674 13758
rect 4622 13682 4674 13694
rect 4846 13746 4898 13758
rect 7410 13709 7422 13761
rect 7474 13709 7486 13761
rect 7746 13694 7758 13746
rect 7810 13694 7822 13746
rect 8082 13694 8094 13746
rect 8146 13694 8158 13746
rect 8418 13721 8430 13773
rect 8482 13721 8494 13773
rect 8766 13746 8818 13758
rect 4846 13682 4898 13694
rect 8766 13682 8818 13694
rect 9438 13746 9490 13758
rect 12002 13750 12014 13802
rect 12066 13750 12078 13802
rect 21460 13783 21512 13795
rect 12238 13746 12290 13758
rect 11666 13694 11678 13746
rect 11730 13694 11742 13746
rect 9438 13682 9490 13694
rect 12238 13682 12290 13694
rect 13806 13746 13858 13758
rect 13806 13682 13858 13694
rect 14030 13746 14082 13758
rect 14030 13682 14082 13694
rect 17278 13746 17330 13758
rect 19730 13694 19742 13746
rect 19794 13694 19806 13746
rect 20066 13721 20078 13773
rect 20130 13721 20142 13773
rect 20414 13746 20466 13758
rect 21758 13746 21810 13758
rect 21460 13719 21512 13731
rect 21634 13694 21646 13746
rect 21698 13694 21710 13746
rect 17278 13682 17330 13694
rect 20414 13682 20466 13694
rect 21758 13682 21810 13694
rect 21086 13634 21138 13646
rect 7298 13582 7310 13634
rect 7362 13582 7374 13634
rect 21086 13570 21138 13582
rect 17614 13522 17666 13534
rect 5114 13470 5126 13522
rect 5178 13470 5190 13522
rect 13514 13470 13526 13522
rect 13578 13470 13590 13522
rect 17614 13458 17666 13470
rect 1344 13354 22624 13388
rect 1344 13302 3874 13354
rect 3926 13302 3978 13354
rect 4030 13302 4082 13354
rect 4134 13302 9194 13354
rect 9246 13302 9298 13354
rect 9350 13302 9402 13354
rect 9454 13302 14514 13354
rect 14566 13302 14618 13354
rect 14670 13302 14722 13354
rect 14774 13302 19834 13354
rect 19886 13302 19938 13354
rect 19990 13302 20042 13354
rect 20094 13302 22624 13354
rect 1344 13268 22624 13302
rect 21982 13186 22034 13198
rect 21982 13122 22034 13134
rect 20806 13074 20858 13086
rect 7410 13022 7422 13074
rect 7474 13022 7486 13074
rect 8866 13022 8878 13074
rect 8930 13022 8942 13074
rect 12338 13022 12350 13074
rect 12402 13022 12414 13074
rect 14242 13022 14254 13074
rect 14306 13022 14318 13074
rect 18050 13022 18062 13074
rect 18114 13022 18126 13074
rect 20806 13010 20858 13022
rect 21478 13074 21530 13086
rect 21478 13010 21530 13022
rect 5182 12962 5234 12974
rect 13806 12962 13858 12974
rect 5182 12898 5234 12910
rect 7522 12866 7534 12918
rect 7586 12866 7598 12918
rect 7858 12910 7870 12962
rect 7922 12910 7934 12962
rect 8530 12910 8542 12962
rect 8594 12910 8606 12962
rect 8754 12866 8766 12918
rect 8818 12866 8830 12918
rect 12002 12910 12014 12962
rect 12066 12910 12078 12962
rect 12226 12895 12238 12947
rect 12290 12895 12302 12947
rect 13806 12898 13858 12910
rect 13918 12962 13970 12974
rect 17054 12962 17106 12974
rect 22318 12962 22370 12974
rect 13918 12898 13970 12910
rect 14354 12895 14366 12947
rect 14418 12895 14430 12947
rect 14690 12910 14702 12962
rect 14754 12910 14766 12962
rect 16370 12910 16382 12962
rect 16434 12910 16446 12962
rect 16830 12923 16882 12935
rect 17602 12910 17614 12962
rect 17666 12910 17678 12962
rect 17054 12898 17106 12910
rect 16830 12859 16882 12871
rect 17938 12866 17950 12918
rect 18002 12866 18014 12918
rect 22318 12898 22370 12910
rect 13514 12798 13526 12850
rect 13578 12798 13590 12850
rect 4846 12738 4898 12750
rect 17154 12742 17166 12794
rect 17218 12742 17230 12794
rect 4846 12674 4898 12686
rect 1344 12570 22784 12604
rect 1344 12518 6534 12570
rect 6586 12518 6638 12570
rect 6690 12518 6742 12570
rect 6794 12518 11854 12570
rect 11906 12518 11958 12570
rect 12010 12518 12062 12570
rect 12114 12518 17174 12570
rect 17226 12518 17278 12570
rect 17330 12518 17382 12570
rect 17434 12518 22494 12570
rect 22546 12518 22598 12570
rect 22650 12518 22702 12570
rect 22754 12518 22784 12570
rect 1344 12484 22784 12518
rect 3502 12402 3554 12414
rect 3502 12338 3554 12350
rect 11566 12402 11618 12414
rect 11566 12338 11618 12350
rect 15318 12402 15370 12414
rect 9998 12290 10050 12302
rect 14018 12294 14030 12346
rect 14082 12294 14094 12346
rect 15318 12338 15370 12350
rect 9998 12226 10050 12238
rect 3166 12178 3218 12190
rect 8642 12141 8654 12193
rect 8706 12141 8718 12193
rect 9886 12178 9938 12190
rect 8866 12126 8878 12178
rect 8930 12126 8942 12178
rect 3166 12114 3218 12126
rect 9886 12114 9938 12126
rect 10166 12178 10218 12190
rect 10166 12114 10218 12126
rect 10334 12178 10386 12190
rect 10334 12114 10386 12126
rect 11902 12178 11954 12190
rect 11902 12114 11954 12126
rect 12014 12178 12066 12190
rect 12014 12114 12066 12126
rect 12238 12178 12290 12190
rect 13234 12126 13246 12178
rect 13298 12126 13310 12178
rect 13570 12153 13582 12205
rect 13634 12153 13646 12205
rect 13918 12178 13970 12190
rect 18062 12178 18114 12190
rect 18622 12178 18674 12190
rect 15138 12126 15150 12178
rect 15202 12126 15214 12178
rect 18330 12126 18342 12178
rect 18394 12126 18406 12178
rect 12238 12114 12290 12126
rect 13918 12114 13970 12126
rect 18062 12114 18114 12126
rect 18622 12114 18674 12126
rect 18734 12178 18786 12190
rect 19338 12182 19350 12234
rect 19402 12182 19414 12234
rect 19058 12126 19070 12178
rect 19122 12126 19134 12178
rect 19842 12126 19854 12178
rect 19906 12126 19918 12178
rect 20178 12170 20190 12222
rect 20242 12170 20254 12222
rect 18734 12114 18786 12126
rect 8530 12014 8542 12066
rect 8594 12014 8606 12066
rect 19506 12014 19518 12066
rect 19570 12014 19582 12066
rect 20290 12014 20302 12066
rect 20354 12014 20366 12066
rect 20738 12014 20750 12066
rect 20802 12063 20814 12066
rect 21410 12063 21422 12066
rect 20802 12017 21422 12063
rect 20802 12014 20814 12017
rect 21410 12014 21422 12017
rect 21474 12014 21486 12066
rect 9606 11954 9658 11966
rect 17726 11954 17778 11966
rect 4386 11902 4398 11954
rect 4450 11951 4462 11954
rect 4834 11951 4846 11954
rect 4450 11905 4846 11951
rect 4450 11902 4462 11905
rect 4834 11902 4846 11905
rect 4898 11902 4910 11954
rect 12506 11902 12518 11954
rect 12570 11902 12582 11954
rect 9606 11890 9658 11902
rect 17726 11890 17778 11902
rect 1344 11786 22624 11820
rect 1344 11734 3874 11786
rect 3926 11734 3978 11786
rect 4030 11734 4082 11786
rect 4134 11734 9194 11786
rect 9246 11734 9298 11786
rect 9350 11734 9402 11786
rect 9454 11734 14514 11786
rect 14566 11734 14618 11786
rect 14670 11734 14722 11786
rect 14774 11734 19834 11786
rect 19886 11734 19938 11786
rect 19990 11734 20042 11786
rect 20094 11734 22624 11786
rect 1344 11700 22624 11734
rect 2924 11618 2976 11630
rect 19114 11566 19126 11618
rect 19178 11566 19190 11618
rect 2924 11554 2976 11566
rect 3670 11450 3722 11462
rect 3166 11394 3218 11406
rect 3670 11386 3722 11398
rect 4846 11394 4898 11406
rect 4274 11342 4286 11394
rect 4338 11342 4350 11394
rect 3166 11330 3218 11342
rect 4498 11315 4510 11367
rect 4562 11315 4574 11367
rect 4846 11330 4898 11342
rect 18622 11394 18674 11406
rect 18622 11330 18674 11342
rect 18846 11394 18898 11406
rect 18846 11330 18898 11342
rect 3838 11282 3890 11294
rect 3838 11218 3890 11230
rect 4274 11174 4286 11226
rect 4338 11174 4350 11226
rect 1344 11002 22784 11036
rect 1344 10950 6534 11002
rect 6586 10950 6638 11002
rect 6690 10950 6742 11002
rect 6794 10950 11854 11002
rect 11906 10950 11958 11002
rect 12010 10950 12062 11002
rect 12114 10950 17174 11002
rect 17226 10950 17278 11002
rect 17330 10950 17382 11002
rect 17434 10950 22494 11002
rect 22546 10950 22598 11002
rect 22650 10950 22702 11002
rect 22754 10950 22784 11002
rect 1344 10916 22784 10950
rect 17950 10834 18002 10846
rect 17950 10770 18002 10782
rect 3950 10722 4002 10734
rect 3546 10614 3558 10666
rect 3610 10614 3622 10666
rect 3950 10658 4002 10670
rect 4118 10666 4170 10678
rect 3714 10558 3726 10610
rect 3778 10558 3790 10610
rect 4118 10602 4170 10614
rect 18286 10610 18338 10622
rect 18286 10546 18338 10558
rect 22318 10610 22370 10622
rect 22318 10546 22370 10558
rect 21590 10498 21642 10510
rect 21590 10434 21642 10446
rect 21982 10386 22034 10398
rect 21982 10322 22034 10334
rect 1344 10218 22624 10252
rect 1344 10166 3874 10218
rect 3926 10166 3978 10218
rect 4030 10166 4082 10218
rect 4134 10166 9194 10218
rect 9246 10166 9298 10218
rect 9350 10166 9402 10218
rect 9454 10166 14514 10218
rect 14566 10166 14618 10218
rect 14670 10166 14722 10218
rect 14774 10166 19834 10218
rect 19886 10166 19938 10218
rect 19990 10166 20042 10218
rect 20094 10166 22624 10218
rect 1344 10132 22624 10166
rect 18174 10050 18226 10062
rect 18174 9986 18226 9998
rect 21422 10050 21474 10062
rect 21422 9986 21474 9998
rect 6302 9938 6354 9950
rect 4230 9882 4282 9894
rect 14018 9886 14030 9938
rect 14082 9886 14094 9938
rect 6302 9874 6354 9886
rect 4230 9818 4282 9830
rect 8766 9826 8818 9838
rect 17838 9826 17890 9838
rect 20526 9826 20578 9838
rect 4610 9774 4622 9826
rect 4674 9774 4686 9826
rect 4958 9770 5010 9782
rect 4398 9714 4450 9726
rect 4958 9706 5010 9718
rect 5742 9770 5794 9782
rect 6066 9774 6078 9826
rect 6130 9774 6142 9826
rect 5742 9706 5794 9718
rect 6470 9770 6522 9782
rect 8194 9774 8206 9826
rect 8258 9774 8270 9826
rect 9426 9774 9438 9826
rect 9490 9774 9502 9826
rect 13570 9774 13582 9826
rect 13634 9774 13646 9826
rect 8766 9762 8818 9774
rect 13906 9759 13918 9811
rect 13970 9759 13982 9811
rect 19058 9774 19070 9826
rect 19122 9774 19134 9826
rect 17838 9762 17890 9774
rect 20526 9762 20578 9774
rect 20862 9826 20914 9838
rect 20862 9762 20914 9774
rect 21814 9826 21866 9838
rect 22094 9826 22146 9838
rect 21970 9774 21982 9826
rect 22034 9774 22046 9826
rect 21814 9762 21866 9774
rect 22094 9762 22146 9774
rect 6470 9706 6522 9718
rect 6918 9714 6970 9726
rect 4398 9650 4450 9662
rect 6918 9650 6970 9662
rect 19462 9714 19514 9726
rect 8374 9602 8426 9614
rect 9538 9606 9550 9658
rect 9602 9606 9614 9658
rect 19462 9650 19514 9662
rect 8374 9538 8426 9550
rect 18902 9602 18954 9614
rect 18902 9538 18954 9550
rect 1344 9434 22784 9468
rect 1344 9382 6534 9434
rect 6586 9382 6638 9434
rect 6690 9382 6742 9434
rect 6794 9382 11854 9434
rect 11906 9382 11958 9434
rect 12010 9382 12062 9434
rect 12114 9382 17174 9434
rect 17226 9382 17278 9434
rect 17330 9382 17382 9434
rect 17434 9382 22494 9434
rect 22546 9382 22598 9434
rect 22650 9382 22702 9434
rect 22754 9382 22784 9434
rect 1344 9348 22784 9382
rect 20638 9266 20690 9278
rect 9550 9154 9602 9166
rect 9550 9090 9602 9102
rect 13526 9154 13578 9166
rect 18498 9158 18510 9210
rect 18562 9158 18574 9210
rect 20638 9202 20690 9214
rect 13526 9090 13578 9102
rect 14366 9098 14418 9110
rect 4722 8990 4734 9042
rect 4786 8990 4798 9042
rect 5058 8990 5070 9042
rect 5122 8990 5134 9042
rect 7410 8990 7422 9042
rect 7474 8990 7486 9042
rect 7746 8990 7758 9042
rect 7810 8990 7822 9042
rect 8418 9018 8430 9070
rect 8482 9018 8494 9070
rect 10222 9042 10274 9054
rect 8642 8990 8654 9042
rect 8706 8990 8718 9042
rect 9046 8986 9098 8998
rect 5686 8930 5738 8942
rect 5182 8874 5234 8886
rect 8878 8930 8930 8942
rect 5686 8866 5738 8878
rect 7870 8874 7922 8886
rect 5182 8810 5234 8822
rect 9046 8922 9098 8934
rect 9718 8986 9770 8998
rect 10222 8978 10274 8990
rect 10782 9042 10834 9054
rect 10782 8978 10834 8990
rect 11006 9042 11058 9054
rect 12338 8990 12350 9042
rect 12402 8990 12414 9042
rect 13014 9028 13026 9080
rect 13078 9028 13090 9080
rect 13806 9070 13858 9082
rect 13806 9006 13858 9018
rect 14030 9070 14082 9082
rect 14030 9006 14082 9018
rect 14254 9070 14306 9082
rect 14960 9080 15012 9092
rect 14366 9034 14418 9046
rect 14702 9042 14754 9054
rect 14254 9006 14306 9018
rect 14802 8990 14814 9042
rect 14866 8990 14878 9042
rect 18174 9081 18226 9093
rect 14960 9016 15012 9028
rect 17950 9042 18002 9054
rect 18958 9042 19010 9054
rect 19406 9042 19458 9054
rect 18174 9017 18226 9029
rect 18610 8990 18622 9042
rect 18674 8990 18686 9042
rect 11006 8978 11058 8990
rect 14702 8978 14754 8990
rect 17950 8978 18002 8990
rect 18958 8978 19010 8990
rect 19126 8986 19178 8998
rect 19282 8990 19294 9042
rect 19346 8990 19358 9042
rect 9718 8922 9770 8934
rect 19406 8978 19458 8990
rect 19686 9042 19738 9054
rect 19686 8978 19738 8990
rect 20302 9042 20354 9054
rect 20302 8978 20354 8990
rect 11274 8878 11286 8930
rect 11338 8878 11350 8930
rect 19126 8922 19178 8934
rect 8878 8866 8930 8878
rect 12238 8874 12290 8886
rect 7870 8810 7922 8822
rect 10464 8818 10516 8830
rect 12238 8810 12290 8822
rect 15374 8818 15426 8830
rect 10464 8754 10516 8766
rect 15374 8754 15426 8766
rect 1344 8650 22624 8684
rect 1344 8598 3874 8650
rect 3926 8598 3978 8650
rect 4030 8598 4082 8650
rect 4134 8598 9194 8650
rect 9246 8598 9298 8650
rect 9350 8598 9402 8650
rect 9454 8598 14514 8650
rect 14566 8598 14618 8650
rect 14670 8598 14722 8650
rect 14774 8598 19834 8650
rect 19886 8598 19938 8650
rect 19990 8598 20042 8650
rect 20094 8598 22624 8650
rect 1344 8564 22624 8598
rect 3950 8482 4002 8494
rect 3950 8418 4002 8430
rect 9830 8482 9882 8494
rect 10452 8430 10464 8482
rect 10516 8479 10528 8482
rect 10994 8479 11006 8482
rect 10516 8433 11006 8479
rect 10516 8430 10528 8433
rect 10994 8430 11006 8433
rect 11058 8430 11070 8482
rect 13850 8430 13862 8482
rect 13914 8430 13926 8482
rect 9830 8418 9882 8430
rect 5126 8370 5178 8382
rect 5126 8306 5178 8318
rect 5798 8370 5850 8382
rect 5798 8306 5850 8318
rect 8206 8370 8258 8382
rect 8206 8306 8258 8318
rect 18230 8314 18282 8326
rect 4622 8258 4674 8270
rect 3490 8206 3502 8258
rect 3554 8206 3566 8258
rect 4498 8206 4510 8258
rect 4562 8206 4574 8258
rect 4330 8150 4342 8202
rect 4394 8150 4406 8202
rect 4622 8194 4674 8206
rect 8542 8258 8594 8270
rect 8542 8194 8594 8206
rect 9102 8258 9154 8270
rect 9550 8258 9602 8270
rect 9426 8206 9438 8258
rect 9490 8206 9502 8258
rect 9102 8194 9154 8206
rect 9258 8150 9270 8202
rect 9322 8150 9334 8202
rect 9550 8194 9602 8206
rect 13358 8258 13410 8270
rect 13358 8194 13410 8206
rect 13582 8258 13634 8270
rect 13582 8194 13634 8206
rect 17502 8220 17554 8232
rect 17826 8206 17838 8258
rect 17890 8206 17902 8258
rect 18230 8250 18282 8262
rect 18454 8258 18506 8270
rect 21982 8258 22034 8270
rect 18834 8206 18846 8258
rect 18898 8206 18910 8258
rect 18454 8194 18506 8206
rect 17502 8156 17554 8168
rect 18062 8146 18114 8158
rect 18062 8082 18114 8094
rect 18622 8146 18674 8158
rect 19058 8150 19070 8202
rect 19122 8150 19134 8202
rect 21982 8194 22034 8206
rect 22318 8258 22370 8270
rect 22318 8194 22370 8206
rect 18622 8082 18674 8094
rect 21590 8146 21642 8158
rect 21590 8082 21642 8094
rect 3334 8034 3386 8046
rect 3334 7970 3386 7982
rect 1344 7866 22784 7900
rect 1344 7814 6534 7866
rect 6586 7814 6638 7866
rect 6690 7814 6742 7866
rect 6794 7814 11854 7866
rect 11906 7814 11958 7866
rect 12010 7814 12062 7866
rect 12114 7814 17174 7866
rect 17226 7814 17278 7866
rect 17330 7814 17382 7866
rect 17434 7814 22494 7866
rect 22546 7814 22598 7866
rect 22650 7814 22702 7866
rect 22754 7814 22784 7866
rect 1344 7780 22784 7814
rect 4678 7698 4730 7710
rect 4678 7634 4730 7646
rect 17894 7698 17946 7710
rect 17894 7634 17946 7646
rect 18342 7698 18394 7710
rect 18342 7634 18394 7646
rect 4174 7586 4226 7598
rect 3894 7530 3946 7542
rect 3378 7452 3390 7504
rect 3442 7452 3454 7504
rect 3602 7461 3614 7513
rect 3666 7461 3678 7513
rect 4174 7522 4226 7534
rect 20246 7530 20298 7542
rect 3894 7466 3946 7478
rect 5238 7474 5290 7486
rect 4498 7422 4510 7474
rect 4562 7422 4574 7474
rect 18050 7422 18062 7474
rect 18114 7422 18126 7474
rect 18498 7422 18510 7474
rect 18562 7422 18574 7474
rect 20246 7466 20298 7478
rect 20974 7530 21026 7542
rect 20626 7422 20638 7474
rect 20690 7422 20702 7474
rect 20974 7466 21026 7478
rect 5238 7410 5290 7422
rect 20414 7362 20466 7374
rect 20414 7298 20466 7310
rect 1344 7082 22624 7116
rect 1344 7030 3874 7082
rect 3926 7030 3978 7082
rect 4030 7030 4082 7082
rect 4134 7030 9194 7082
rect 9246 7030 9298 7082
rect 9350 7030 9402 7082
rect 9454 7030 14514 7082
rect 14566 7030 14618 7082
rect 14670 7030 14722 7082
rect 14774 7030 19834 7082
rect 19886 7030 19938 7082
rect 19990 7030 20042 7082
rect 20094 7030 22624 7082
rect 1344 6996 22624 7030
rect 7590 6746 7642 6758
rect 7590 6682 7642 6694
rect 7758 6690 7810 6702
rect 7970 6638 7982 6690
rect 8034 6638 8046 6690
rect 7758 6626 7810 6638
rect 8194 6610 8206 6662
rect 8258 6610 8270 6662
rect 1344 6298 22784 6332
rect 1344 6246 6534 6298
rect 6586 6246 6638 6298
rect 6690 6246 6742 6298
rect 6794 6246 11854 6298
rect 11906 6246 11958 6298
rect 12010 6246 12062 6298
rect 12114 6246 17174 6298
rect 17226 6246 17278 6298
rect 17330 6246 17382 6298
rect 17434 6246 22494 6298
rect 22546 6246 22598 6298
rect 22650 6246 22702 6298
rect 22754 6246 22784 6298
rect 1344 6212 22784 6246
rect 15038 6130 15090 6142
rect 3614 6018 3666 6030
rect 3614 5954 3666 5966
rect 8206 6018 8258 6030
rect 11330 6022 11342 6074
rect 11394 6022 11406 6074
rect 15038 6066 15090 6078
rect 20414 6130 20466 6142
rect 20414 6066 20466 6078
rect 14186 5966 14198 6018
rect 14250 5966 14262 6018
rect 3845 5910 3857 5962
rect 3909 5910 3921 5962
rect 8206 5954 8258 5966
rect 4734 5906 4786 5918
rect 4734 5842 4786 5854
rect 6806 5906 6858 5918
rect 7086 5906 7138 5918
rect 6962 5854 6974 5906
rect 7026 5854 7038 5906
rect 6806 5842 6858 5854
rect 7086 5842 7138 5854
rect 8094 5906 8146 5918
rect 8362 5910 8374 5962
rect 8426 5910 8438 5962
rect 8094 5842 8146 5854
rect 8542 5906 8594 5918
rect 11218 5854 11230 5906
rect 11282 5854 11294 5906
rect 11554 5869 11566 5921
rect 11618 5869 11630 5921
rect 14478 5906 14530 5918
rect 11890 5854 11902 5906
rect 11954 5854 11966 5906
rect 8542 5842 8594 5854
rect 14478 5842 14530 5854
rect 14590 5906 14642 5918
rect 14590 5842 14642 5854
rect 15374 5906 15426 5918
rect 15374 5842 15426 5854
rect 19406 5906 19458 5918
rect 19406 5842 19458 5854
rect 19518 5906 19570 5918
rect 19518 5842 19570 5854
rect 20078 5906 20130 5918
rect 20078 5842 20130 5854
rect 6414 5682 6466 5694
rect 6414 5618 6466 5630
rect 7814 5682 7866 5694
rect 7814 5618 7866 5630
rect 12070 5682 12122 5694
rect 19786 5630 19798 5682
rect 19850 5630 19862 5682
rect 12070 5618 12122 5630
rect 1344 5514 22624 5548
rect 1344 5462 3874 5514
rect 3926 5462 3978 5514
rect 4030 5462 4082 5514
rect 4134 5462 9194 5514
rect 9246 5462 9298 5514
rect 9350 5462 9402 5514
rect 9454 5462 14514 5514
rect 14566 5462 14618 5514
rect 14670 5462 14722 5514
rect 14774 5462 19834 5514
rect 19886 5462 19938 5514
rect 19990 5462 20042 5514
rect 20094 5462 22624 5514
rect 1344 5428 22624 5462
rect 8318 5346 8370 5358
rect 8318 5282 8370 5294
rect 8878 5346 8930 5358
rect 8878 5282 8930 5294
rect 13526 5346 13578 5358
rect 13526 5282 13578 5294
rect 20526 5346 20578 5358
rect 9606 5234 9658 5246
rect 7366 5178 7418 5190
rect 3502 5122 3554 5134
rect 3502 5058 3554 5070
rect 4622 5122 4674 5134
rect 6514 5126 6526 5178
rect 6578 5126 6590 5178
rect 7198 5122 7250 5134
rect 4366 5014 4378 5066
rect 4430 5014 4442 5066
rect 4622 5058 4674 5070
rect 6738 5042 6750 5094
rect 6802 5042 6814 5094
rect 9606 5170 9658 5182
rect 12014 5234 12066 5246
rect 15598 5234 15650 5246
rect 12674 5182 12686 5234
rect 12738 5182 12750 5234
rect 12014 5170 12066 5182
rect 15598 5170 15650 5182
rect 17166 5234 17218 5246
rect 18610 5238 18622 5290
rect 18674 5238 18686 5290
rect 20526 5282 20578 5294
rect 17166 5170 17218 5182
rect 21982 5234 22034 5246
rect 21982 5170 22034 5182
rect 7366 5114 7418 5126
rect 7646 5122 7698 5134
rect 7926 5122 7978 5134
rect 7198 5058 7250 5070
rect 7746 5070 7758 5122
rect 7810 5070 7822 5122
rect 7646 5058 7698 5070
rect 7926 5058 7978 5070
rect 9214 5122 9266 5134
rect 13806 5122 13858 5134
rect 10658 5070 10670 5122
rect 10722 5070 10734 5122
rect 10994 5070 11006 5122
rect 11058 5070 11070 5122
rect 11554 5070 11566 5122
rect 11618 5070 11630 5122
rect 11778 5070 11790 5122
rect 11842 5070 11854 5122
rect 12226 5070 12238 5122
rect 12290 5070 12302 5122
rect 9214 5058 9266 5070
rect 12562 5055 12574 5107
rect 12626 5055 12638 5107
rect 13682 5070 13694 5122
rect 13746 5070 13758 5122
rect 13806 5058 13858 5070
rect 14030 5122 14082 5134
rect 14030 5058 14082 5070
rect 15262 5122 15314 5134
rect 16830 5122 16882 5134
rect 20862 5122 20914 5134
rect 15262 5058 15314 5070
rect 15486 5083 15538 5095
rect 15922 5070 15934 5122
rect 15986 5070 15998 5122
rect 17714 5070 17726 5122
rect 17778 5070 17790 5122
rect 16830 5058 16882 5070
rect 18050 5055 18062 5107
rect 18114 5055 18126 5107
rect 18498 5070 18510 5122
rect 18562 5070 18574 5122
rect 18834 5070 18846 5122
rect 18898 5070 18910 5122
rect 19282 5070 19294 5122
rect 19346 5070 19358 5122
rect 19574 5092 19626 5104
rect 15486 5019 15538 5031
rect 20862 5058 20914 5070
rect 21590 5122 21642 5134
rect 21590 5058 21642 5070
rect 22318 5122 22370 5134
rect 22318 5058 22370 5070
rect 19574 5028 19626 5040
rect 14298 4958 14310 5010
rect 14362 4958 14374 5010
rect 19630 4954 19682 4966
rect 17826 4902 17838 4954
rect 17890 4902 17902 4954
rect 19630 4890 19682 4902
rect 1344 4730 22784 4764
rect 1344 4678 6534 4730
rect 6586 4678 6638 4730
rect 6690 4678 6742 4730
rect 6794 4678 11854 4730
rect 11906 4678 11958 4730
rect 12010 4678 12062 4730
rect 12114 4678 17174 4730
rect 17226 4678 17278 4730
rect 17330 4678 17382 4730
rect 17434 4678 22494 4730
rect 22546 4678 22598 4730
rect 22650 4678 22702 4730
rect 22754 4678 22784 4730
rect 1344 4644 22784 4678
rect 4790 4562 4842 4574
rect 4790 4498 4842 4510
rect 7758 4562 7810 4574
rect 7758 4498 7810 4510
rect 8710 4562 8762 4574
rect 8710 4498 8762 4510
rect 13638 4562 13690 4574
rect 13638 4498 13690 4510
rect 14142 4562 14194 4574
rect 14142 4498 14194 4510
rect 17446 4562 17498 4574
rect 17446 4498 17498 4510
rect 19406 4562 19458 4574
rect 19406 4498 19458 4510
rect 4174 4450 4226 4462
rect 3054 4338 3106 4350
rect 3918 4342 3930 4394
rect 3982 4342 3994 4394
rect 4174 4386 4226 4398
rect 12014 4450 12066 4462
rect 12014 4386 12066 4398
rect 12574 4394 12626 4406
rect 20010 4398 20022 4450
rect 20074 4398 20086 4450
rect 3054 4274 3106 4286
rect 8094 4338 8146 4350
rect 8094 4274 8146 4286
rect 11622 4338 11674 4350
rect 11622 4274 11674 4286
rect 11846 4338 11898 4350
rect 12226 4286 12238 4338
rect 12290 4286 12302 4338
rect 12574 4330 12626 4342
rect 14478 4338 14530 4350
rect 19742 4338 19794 4350
rect 17602 4286 17614 4338
rect 17666 4286 17678 4338
rect 11846 4274 11898 4286
rect 14478 4274 14530 4286
rect 19742 4274 19794 4286
rect 20302 4338 20354 4350
rect 20302 4274 20354 4286
rect 20526 4338 20578 4350
rect 20850 4286 20862 4338
rect 20914 4286 20926 4338
rect 21186 4286 21198 4338
rect 21250 4286 21262 4338
rect 20526 4274 20578 4286
rect 21702 4226 21754 4238
rect 20750 4170 20802 4182
rect 21702 4162 21754 4174
rect 22150 4226 22202 4238
rect 22150 4162 22202 4174
rect 20750 4106 20802 4118
rect 1344 3946 22624 3980
rect 1344 3894 3874 3946
rect 3926 3894 3978 3946
rect 4030 3894 4082 3946
rect 4134 3894 9194 3946
rect 9246 3894 9298 3946
rect 9350 3894 9402 3946
rect 9454 3894 14514 3946
rect 14566 3894 14618 3946
rect 14670 3894 14722 3946
rect 14774 3894 19834 3946
rect 19886 3894 19938 3946
rect 19990 3894 20042 3946
rect 20094 3894 22624 3946
rect 1344 3860 22624 3894
rect 1344 3162 22784 3196
rect 1344 3110 6534 3162
rect 6586 3110 6638 3162
rect 6690 3110 6742 3162
rect 6794 3110 11854 3162
rect 11906 3110 11958 3162
rect 12010 3110 12062 3162
rect 12114 3110 17174 3162
rect 17226 3110 17278 3162
rect 17330 3110 17382 3162
rect 17434 3110 22494 3162
rect 22546 3110 22598 3162
rect 22650 3110 22702 3162
rect 22754 3110 22784 3162
rect 1344 3076 22784 3110
<< via1 >>
rect 6534 20358 6586 20410
rect 6638 20358 6690 20410
rect 6742 20358 6794 20410
rect 11854 20358 11906 20410
rect 11958 20358 12010 20410
rect 12062 20358 12114 20410
rect 17174 20358 17226 20410
rect 17278 20358 17330 20410
rect 17382 20358 17434 20410
rect 22494 20358 22546 20410
rect 22598 20358 22650 20410
rect 22702 20358 22754 20410
rect 2158 20078 2210 20130
rect 4510 20078 4562 20130
rect 6750 20078 6802 20130
rect 9550 20078 9602 20130
rect 11230 20078 11282 20130
rect 13358 20078 13410 20130
rect 15710 20078 15762 20130
rect 17950 20078 18002 20130
rect 20078 20078 20130 20130
rect 20974 20078 21026 20130
rect 22094 20078 22146 20130
rect 2494 19966 2546 20018
rect 4174 19966 4226 20018
rect 6414 19966 6466 20018
rect 9214 19966 9266 20018
rect 10894 19966 10946 20018
rect 13694 19966 13746 20018
rect 15374 19966 15426 20018
rect 17614 19966 17666 20018
rect 19742 19966 19794 20018
rect 20638 19966 20690 20018
rect 21758 19966 21810 20018
rect 3874 19574 3926 19626
rect 3978 19574 4030 19626
rect 4082 19574 4134 19626
rect 9194 19574 9246 19626
rect 9298 19574 9350 19626
rect 9402 19574 9454 19626
rect 14514 19574 14566 19626
rect 14618 19574 14670 19626
rect 14722 19574 14774 19626
rect 19834 19574 19886 19626
rect 19938 19574 19990 19626
rect 20042 19574 20094 19626
rect 3054 19406 3106 19458
rect 3726 19406 3778 19458
rect 4510 19406 4562 19458
rect 5854 19406 5906 19458
rect 10894 19406 10946 19458
rect 15150 19406 15202 19458
rect 14254 19350 14306 19402
rect 16382 19406 16434 19458
rect 18622 19406 18674 19458
rect 21534 19406 21586 19458
rect 3390 19182 3442 19234
rect 4062 19182 4114 19234
rect 4174 19182 4226 19234
rect 5182 19182 5234 19234
rect 5518 19182 5570 19234
rect 7982 19182 8034 19234
rect 8654 19182 8706 19234
rect 9102 19182 9154 19234
rect 11230 19182 11282 19234
rect 14142 19182 14194 19234
rect 14478 19182 14530 19234
rect 14814 19182 14866 19234
rect 16046 19182 16098 19234
rect 18286 19182 18338 19234
rect 19070 19182 19122 19234
rect 19742 19182 19794 19234
rect 20078 19182 20130 19234
rect 21198 19182 21250 19234
rect 5014 19014 5066 19066
rect 8542 19014 8594 19066
rect 9438 18958 9490 19010
rect 19518 19014 19570 19066
rect 15766 18958 15818 19010
rect 20414 18958 20466 19010
rect 6534 18790 6586 18842
rect 6638 18790 6690 18842
rect 6742 18790 6794 18842
rect 11854 18790 11906 18842
rect 11958 18790 12010 18842
rect 12062 18790 12114 18842
rect 17174 18790 17226 18842
rect 17278 18790 17330 18842
rect 17382 18790 17434 18842
rect 22494 18790 22546 18842
rect 22598 18790 22650 18842
rect 22702 18790 22754 18842
rect 11006 18622 11058 18674
rect 8878 18566 8930 18618
rect 15038 18622 15090 18674
rect 14422 18510 14474 18562
rect 20134 18510 20186 18562
rect 7422 18398 7474 18450
rect 7646 18413 7698 18465
rect 8542 18454 8594 18506
rect 8094 18398 8146 18450
rect 8766 18398 8818 18450
rect 9662 18413 9714 18465
rect 9998 18398 10050 18450
rect 10670 18398 10722 18450
rect 14030 18398 14082 18450
rect 14142 18398 14194 18450
rect 14702 18398 14754 18450
rect 17838 18398 17890 18450
rect 18174 18398 18226 18450
rect 19294 18398 19346 18450
rect 19630 18398 19682 18450
rect 19854 18398 19906 18450
rect 20582 18398 20634 18450
rect 20862 18398 20914 18450
rect 20974 18398 21026 18450
rect 21590 18398 21642 18450
rect 22318 18398 22370 18450
rect 3558 18286 3610 18338
rect 7758 18286 7810 18338
rect 9550 18286 9602 18338
rect 18958 18286 19010 18338
rect 21982 18174 22034 18226
rect 3874 18006 3926 18058
rect 3978 18006 4030 18058
rect 4082 18006 4134 18058
rect 9194 18006 9246 18058
rect 9298 18006 9350 18058
rect 9402 18006 9454 18058
rect 14514 18006 14566 18058
rect 14618 18006 14670 18058
rect 14722 18006 14774 18058
rect 19834 18006 19886 18058
rect 19938 18006 19990 18058
rect 20042 18006 20094 18058
rect 3502 17782 3554 17834
rect 8318 17838 8370 17890
rect 13862 17838 13914 17890
rect 14646 17838 14698 17890
rect 4510 17726 4562 17778
rect 9382 17782 9434 17834
rect 2714 17576 2766 17628
rect 3390 17614 3442 17666
rect 3950 17576 4002 17628
rect 4286 17614 4338 17666
rect 4678 17558 4730 17610
rect 8710 17614 8762 17666
rect 8878 17614 8930 17666
rect 8990 17614 9042 17666
rect 9550 17614 9602 17666
rect 13358 17614 13410 17666
rect 13582 17614 13634 17666
rect 14254 17614 14306 17666
rect 14366 17614 14418 17666
rect 11510 17390 11562 17442
rect 12966 17390 13018 17442
rect 6534 17222 6586 17274
rect 6638 17222 6690 17274
rect 6742 17222 6794 17274
rect 11854 17222 11906 17274
rect 11958 17222 12010 17274
rect 12062 17222 12114 17274
rect 17174 17222 17226 17274
rect 17278 17222 17330 17274
rect 17382 17222 17434 17274
rect 22494 17222 22546 17274
rect 22598 17222 22650 17274
rect 22702 17222 22754 17274
rect 8486 17054 8538 17106
rect 10838 16942 10890 16994
rect 13134 16942 13186 16994
rect 3166 16830 3218 16882
rect 3446 16830 3498 16882
rect 3726 16830 3778 16882
rect 3950 16830 4002 16882
rect 4174 16830 4226 16882
rect 4846 16830 4898 16882
rect 7646 16830 7698 16882
rect 7982 16830 8034 16882
rect 11118 16830 11170 16882
rect 11342 16830 11394 16882
rect 12014 16863 12066 16915
rect 12238 16886 12290 16938
rect 21590 16942 21642 16994
rect 12686 16863 12738 16915
rect 12996 16863 13048 16915
rect 18286 16830 18338 16882
rect 21982 16830 22034 16882
rect 22318 16830 22370 16882
rect 4958 16662 5010 16714
rect 7534 16662 7586 16714
rect 2830 16606 2882 16658
rect 18622 16606 18674 16658
rect 3874 16438 3926 16490
rect 3978 16438 4030 16490
rect 4082 16438 4134 16490
rect 9194 16438 9246 16490
rect 9298 16438 9350 16490
rect 9402 16438 9454 16490
rect 14514 16438 14566 16490
rect 14618 16438 14670 16490
rect 14722 16438 14774 16490
rect 19834 16438 19886 16490
rect 19938 16438 19990 16490
rect 20042 16438 20094 16490
rect 18230 16270 18282 16322
rect 19350 16270 19402 16322
rect 3166 16214 3218 16266
rect 4286 16214 4338 16266
rect 11622 16158 11674 16210
rect 3390 16046 3442 16098
rect 3950 16046 4002 16098
rect 4398 16046 4450 16098
rect 4622 16046 4674 16098
rect 14254 16046 14306 16098
rect 14926 16046 14978 16098
rect 14702 15990 14754 16042
rect 15374 16046 15426 16098
rect 18510 16046 18562 16098
rect 18734 16046 18786 16098
rect 18846 16046 18898 16098
rect 19070 16046 19122 16098
rect 15038 15878 15090 15930
rect 15710 15822 15762 15874
rect 6534 15654 6586 15706
rect 6638 15654 6690 15706
rect 6742 15654 6794 15706
rect 11854 15654 11906 15706
rect 11958 15654 12010 15706
rect 12062 15654 12114 15706
rect 17174 15654 17226 15706
rect 17278 15654 17330 15706
rect 17382 15654 17434 15706
rect 22494 15654 22546 15706
rect 22598 15654 22650 15706
rect 22702 15654 22754 15706
rect 3614 15430 3666 15482
rect 12686 15430 12738 15482
rect 19182 15430 19234 15482
rect 20414 15430 20466 15482
rect 3502 15262 3554 15314
rect 3838 15306 3890 15358
rect 12238 15262 12290 15314
rect 12574 15301 12626 15353
rect 12798 15262 12850 15314
rect 14926 15277 14978 15329
rect 15262 15262 15314 15314
rect 18286 15262 18338 15314
rect 18510 15306 18562 15358
rect 19070 15262 19122 15314
rect 19406 15277 19458 15329
rect 20918 15318 20970 15370
rect 20526 15262 20578 15314
rect 21198 15262 21250 15314
rect 14814 15150 14866 15202
rect 18622 15150 18674 15202
rect 3874 14870 3926 14922
rect 3978 14870 4030 14922
rect 4082 14870 4134 14922
rect 9194 14870 9246 14922
rect 9298 14870 9350 14922
rect 9402 14870 9454 14922
rect 14514 14870 14566 14922
rect 14618 14870 14670 14922
rect 14722 14870 14774 14922
rect 19834 14870 19886 14922
rect 19938 14870 19990 14922
rect 20042 14870 20094 14922
rect 4678 14702 4730 14754
rect 5798 14590 5850 14642
rect 4958 14478 5010 14530
rect 5182 14478 5234 14530
rect 8654 14478 8706 14530
rect 13806 14478 13858 14530
rect 14030 14478 14082 14530
rect 21198 14478 21250 14530
rect 13526 14366 13578 14418
rect 8318 14254 8370 14306
rect 8990 14254 9042 14306
rect 9774 14254 9826 14306
rect 21534 14254 21586 14306
rect 6534 14086 6586 14138
rect 6638 14086 6690 14138
rect 6742 14086 6794 14138
rect 11854 14086 11906 14138
rect 11958 14086 12010 14138
rect 12062 14086 12114 14138
rect 17174 14086 17226 14138
rect 17278 14086 17330 14138
rect 17382 14086 17434 14138
rect 22494 14086 22546 14138
rect 22598 14086 22650 14138
rect 22702 14086 22754 14138
rect 5686 13918 5738 13970
rect 9774 13918 9826 13970
rect 8878 13862 8930 13914
rect 11790 13862 11842 13914
rect 20526 13862 20578 13914
rect 4174 13806 4226 13858
rect 4510 13694 4562 13746
rect 4622 13694 4674 13746
rect 4846 13694 4898 13746
rect 7422 13709 7474 13761
rect 7758 13694 7810 13746
rect 8094 13694 8146 13746
rect 8430 13721 8482 13773
rect 8766 13694 8818 13746
rect 12014 13750 12066 13802
rect 9438 13694 9490 13746
rect 11678 13694 11730 13746
rect 12238 13694 12290 13746
rect 13806 13694 13858 13746
rect 14030 13694 14082 13746
rect 17278 13694 17330 13746
rect 19742 13694 19794 13746
rect 20078 13721 20130 13773
rect 20414 13694 20466 13746
rect 21460 13731 21512 13783
rect 21646 13694 21698 13746
rect 21758 13694 21810 13746
rect 7310 13582 7362 13634
rect 21086 13582 21138 13634
rect 5126 13470 5178 13522
rect 13526 13470 13578 13522
rect 17614 13470 17666 13522
rect 3874 13302 3926 13354
rect 3978 13302 4030 13354
rect 4082 13302 4134 13354
rect 9194 13302 9246 13354
rect 9298 13302 9350 13354
rect 9402 13302 9454 13354
rect 14514 13302 14566 13354
rect 14618 13302 14670 13354
rect 14722 13302 14774 13354
rect 19834 13302 19886 13354
rect 19938 13302 19990 13354
rect 20042 13302 20094 13354
rect 21982 13134 22034 13186
rect 7422 13022 7474 13074
rect 8878 13022 8930 13074
rect 12350 13022 12402 13074
rect 14254 13022 14306 13074
rect 18062 13022 18114 13074
rect 20806 13022 20858 13074
rect 21478 13022 21530 13074
rect 5182 12910 5234 12962
rect 7534 12866 7586 12918
rect 7870 12910 7922 12962
rect 8542 12910 8594 12962
rect 8766 12866 8818 12918
rect 12014 12910 12066 12962
rect 12238 12895 12290 12947
rect 13806 12910 13858 12962
rect 13918 12910 13970 12962
rect 14366 12895 14418 12947
rect 14702 12910 14754 12962
rect 16382 12910 16434 12962
rect 16830 12871 16882 12923
rect 17054 12910 17106 12962
rect 17614 12910 17666 12962
rect 17950 12866 18002 12918
rect 22318 12910 22370 12962
rect 13526 12798 13578 12850
rect 17166 12742 17218 12794
rect 4846 12686 4898 12738
rect 6534 12518 6586 12570
rect 6638 12518 6690 12570
rect 6742 12518 6794 12570
rect 11854 12518 11906 12570
rect 11958 12518 12010 12570
rect 12062 12518 12114 12570
rect 17174 12518 17226 12570
rect 17278 12518 17330 12570
rect 17382 12518 17434 12570
rect 22494 12518 22546 12570
rect 22598 12518 22650 12570
rect 22702 12518 22754 12570
rect 3502 12350 3554 12402
rect 11566 12350 11618 12402
rect 15318 12350 15370 12402
rect 14030 12294 14082 12346
rect 9998 12238 10050 12290
rect 3166 12126 3218 12178
rect 8654 12141 8706 12193
rect 8878 12126 8930 12178
rect 9886 12126 9938 12178
rect 10166 12126 10218 12178
rect 10334 12126 10386 12178
rect 11902 12126 11954 12178
rect 12014 12126 12066 12178
rect 12238 12126 12290 12178
rect 13246 12126 13298 12178
rect 13582 12153 13634 12205
rect 13918 12126 13970 12178
rect 15150 12126 15202 12178
rect 18062 12126 18114 12178
rect 18342 12126 18394 12178
rect 18622 12126 18674 12178
rect 19350 12182 19402 12234
rect 18734 12126 18786 12178
rect 19070 12126 19122 12178
rect 19854 12126 19906 12178
rect 20190 12170 20242 12222
rect 8542 12014 8594 12066
rect 19518 12014 19570 12066
rect 20302 12014 20354 12066
rect 20750 12014 20802 12066
rect 21422 12014 21474 12066
rect 4398 11902 4450 11954
rect 4846 11902 4898 11954
rect 9606 11902 9658 11954
rect 12518 11902 12570 11954
rect 17726 11902 17778 11954
rect 3874 11734 3926 11786
rect 3978 11734 4030 11786
rect 4082 11734 4134 11786
rect 9194 11734 9246 11786
rect 9298 11734 9350 11786
rect 9402 11734 9454 11786
rect 14514 11734 14566 11786
rect 14618 11734 14670 11786
rect 14722 11734 14774 11786
rect 19834 11734 19886 11786
rect 19938 11734 19990 11786
rect 20042 11734 20094 11786
rect 2924 11566 2976 11618
rect 19126 11566 19178 11618
rect 3166 11342 3218 11394
rect 3670 11398 3722 11450
rect 4286 11342 4338 11394
rect 4510 11315 4562 11367
rect 4846 11342 4898 11394
rect 18622 11342 18674 11394
rect 18846 11342 18898 11394
rect 3838 11230 3890 11282
rect 4286 11174 4338 11226
rect 6534 10950 6586 11002
rect 6638 10950 6690 11002
rect 6742 10950 6794 11002
rect 11854 10950 11906 11002
rect 11958 10950 12010 11002
rect 12062 10950 12114 11002
rect 17174 10950 17226 11002
rect 17278 10950 17330 11002
rect 17382 10950 17434 11002
rect 22494 10950 22546 11002
rect 22598 10950 22650 11002
rect 22702 10950 22754 11002
rect 17950 10782 18002 10834
rect 3950 10670 4002 10722
rect 3558 10614 3610 10666
rect 4118 10614 4170 10666
rect 3726 10558 3778 10610
rect 18286 10558 18338 10610
rect 22318 10558 22370 10610
rect 21590 10446 21642 10498
rect 21982 10334 22034 10386
rect 3874 10166 3926 10218
rect 3978 10166 4030 10218
rect 4082 10166 4134 10218
rect 9194 10166 9246 10218
rect 9298 10166 9350 10218
rect 9402 10166 9454 10218
rect 14514 10166 14566 10218
rect 14618 10166 14670 10218
rect 14722 10166 14774 10218
rect 19834 10166 19886 10218
rect 19938 10166 19990 10218
rect 20042 10166 20094 10218
rect 18174 9998 18226 10050
rect 21422 9998 21474 10050
rect 4230 9830 4282 9882
rect 6302 9886 6354 9938
rect 14030 9886 14082 9938
rect 4622 9774 4674 9826
rect 4398 9662 4450 9714
rect 4958 9718 5010 9770
rect 6078 9774 6130 9826
rect 5742 9718 5794 9770
rect 8206 9774 8258 9826
rect 8766 9774 8818 9826
rect 9438 9774 9490 9826
rect 13582 9774 13634 9826
rect 6470 9718 6522 9770
rect 13918 9759 13970 9811
rect 17838 9774 17890 9826
rect 19070 9774 19122 9826
rect 20526 9774 20578 9826
rect 20862 9774 20914 9826
rect 21814 9774 21866 9826
rect 21982 9774 22034 9826
rect 22094 9774 22146 9826
rect 6918 9662 6970 9714
rect 19462 9662 19514 9714
rect 9550 9606 9602 9658
rect 8374 9550 8426 9602
rect 18902 9550 18954 9602
rect 6534 9382 6586 9434
rect 6638 9382 6690 9434
rect 6742 9382 6794 9434
rect 11854 9382 11906 9434
rect 11958 9382 12010 9434
rect 12062 9382 12114 9434
rect 17174 9382 17226 9434
rect 17278 9382 17330 9434
rect 17382 9382 17434 9434
rect 22494 9382 22546 9434
rect 22598 9382 22650 9434
rect 22702 9382 22754 9434
rect 20638 9214 20690 9266
rect 9550 9102 9602 9154
rect 18510 9158 18562 9210
rect 13526 9102 13578 9154
rect 4734 8990 4786 9042
rect 5070 8990 5122 9042
rect 7422 8990 7474 9042
rect 7758 8990 7810 9042
rect 8430 9018 8482 9070
rect 8654 8990 8706 9042
rect 5182 8822 5234 8874
rect 5686 8878 5738 8930
rect 7870 8822 7922 8874
rect 8878 8878 8930 8930
rect 9046 8934 9098 8986
rect 9718 8934 9770 8986
rect 10222 8990 10274 9042
rect 10782 8990 10834 9042
rect 11006 8990 11058 9042
rect 12350 8990 12402 9042
rect 13026 9028 13078 9080
rect 13806 9018 13858 9070
rect 14030 9018 14082 9070
rect 14254 9018 14306 9070
rect 14366 9046 14418 9098
rect 14702 8990 14754 9042
rect 14814 8990 14866 9042
rect 14960 9028 15012 9080
rect 17950 8990 18002 9042
rect 18174 9029 18226 9081
rect 18622 8990 18674 9042
rect 18958 8990 19010 9042
rect 19294 8990 19346 9042
rect 19406 8990 19458 9042
rect 19126 8934 19178 8986
rect 19686 8990 19738 9042
rect 20302 8990 20354 9042
rect 11286 8878 11338 8930
rect 10464 8766 10516 8818
rect 12238 8822 12290 8874
rect 15374 8766 15426 8818
rect 3874 8598 3926 8650
rect 3978 8598 4030 8650
rect 4082 8598 4134 8650
rect 9194 8598 9246 8650
rect 9298 8598 9350 8650
rect 9402 8598 9454 8650
rect 14514 8598 14566 8650
rect 14618 8598 14670 8650
rect 14722 8598 14774 8650
rect 19834 8598 19886 8650
rect 19938 8598 19990 8650
rect 20042 8598 20094 8650
rect 3950 8430 4002 8482
rect 9830 8430 9882 8482
rect 10464 8430 10516 8482
rect 11006 8430 11058 8482
rect 13862 8430 13914 8482
rect 5126 8318 5178 8370
rect 5798 8318 5850 8370
rect 8206 8318 8258 8370
rect 3502 8206 3554 8258
rect 4510 8206 4562 8258
rect 4622 8206 4674 8258
rect 4342 8150 4394 8202
rect 8542 8206 8594 8258
rect 9102 8206 9154 8258
rect 9438 8206 9490 8258
rect 9550 8206 9602 8258
rect 9270 8150 9322 8202
rect 13358 8206 13410 8258
rect 18230 8262 18282 8314
rect 13582 8206 13634 8258
rect 17502 8168 17554 8220
rect 17838 8206 17890 8258
rect 18454 8206 18506 8258
rect 18846 8206 18898 8258
rect 21982 8206 22034 8258
rect 18062 8094 18114 8146
rect 19070 8150 19122 8202
rect 22318 8206 22370 8258
rect 18622 8094 18674 8146
rect 21590 8094 21642 8146
rect 3334 7982 3386 8034
rect 6534 7814 6586 7866
rect 6638 7814 6690 7866
rect 6742 7814 6794 7866
rect 11854 7814 11906 7866
rect 11958 7814 12010 7866
rect 12062 7814 12114 7866
rect 17174 7814 17226 7866
rect 17278 7814 17330 7866
rect 17382 7814 17434 7866
rect 22494 7814 22546 7866
rect 22598 7814 22650 7866
rect 22702 7814 22754 7866
rect 4678 7646 4730 7698
rect 17894 7646 17946 7698
rect 18342 7646 18394 7698
rect 3390 7452 3442 7504
rect 3614 7461 3666 7513
rect 3894 7478 3946 7530
rect 4174 7534 4226 7586
rect 20246 7478 20298 7530
rect 4510 7422 4562 7474
rect 5238 7422 5290 7474
rect 18062 7422 18114 7474
rect 18510 7422 18562 7474
rect 20974 7478 21026 7530
rect 20638 7422 20690 7474
rect 20414 7310 20466 7362
rect 3874 7030 3926 7082
rect 3978 7030 4030 7082
rect 4082 7030 4134 7082
rect 9194 7030 9246 7082
rect 9298 7030 9350 7082
rect 9402 7030 9454 7082
rect 14514 7030 14566 7082
rect 14618 7030 14670 7082
rect 14722 7030 14774 7082
rect 19834 7030 19886 7082
rect 19938 7030 19990 7082
rect 20042 7030 20094 7082
rect 7590 6694 7642 6746
rect 7758 6638 7810 6690
rect 7982 6638 8034 6690
rect 8206 6610 8258 6662
rect 6534 6246 6586 6298
rect 6638 6246 6690 6298
rect 6742 6246 6794 6298
rect 11854 6246 11906 6298
rect 11958 6246 12010 6298
rect 12062 6246 12114 6298
rect 17174 6246 17226 6298
rect 17278 6246 17330 6298
rect 17382 6246 17434 6298
rect 22494 6246 22546 6298
rect 22598 6246 22650 6298
rect 22702 6246 22754 6298
rect 15038 6078 15090 6130
rect 3614 5966 3666 6018
rect 11342 6022 11394 6074
rect 20414 6078 20466 6130
rect 8206 5966 8258 6018
rect 14198 5966 14250 6018
rect 3857 5910 3909 5962
rect 4734 5854 4786 5906
rect 6806 5854 6858 5906
rect 6974 5854 7026 5906
rect 7086 5854 7138 5906
rect 8374 5910 8426 5962
rect 8094 5854 8146 5906
rect 8542 5854 8594 5906
rect 11230 5854 11282 5906
rect 11566 5869 11618 5921
rect 11902 5854 11954 5906
rect 14478 5854 14530 5906
rect 14590 5854 14642 5906
rect 15374 5854 15426 5906
rect 19406 5854 19458 5906
rect 19518 5854 19570 5906
rect 20078 5854 20130 5906
rect 6414 5630 6466 5682
rect 7814 5630 7866 5682
rect 12070 5630 12122 5682
rect 19798 5630 19850 5682
rect 3874 5462 3926 5514
rect 3978 5462 4030 5514
rect 4082 5462 4134 5514
rect 9194 5462 9246 5514
rect 9298 5462 9350 5514
rect 9402 5462 9454 5514
rect 14514 5462 14566 5514
rect 14618 5462 14670 5514
rect 14722 5462 14774 5514
rect 19834 5462 19886 5514
rect 19938 5462 19990 5514
rect 20042 5462 20094 5514
rect 8318 5294 8370 5346
rect 8878 5294 8930 5346
rect 13526 5294 13578 5346
rect 20526 5294 20578 5346
rect 3502 5070 3554 5122
rect 6526 5126 6578 5178
rect 4622 5070 4674 5122
rect 4378 5014 4430 5066
rect 6750 5042 6802 5094
rect 7198 5070 7250 5122
rect 7366 5126 7418 5178
rect 9606 5182 9658 5234
rect 12014 5182 12066 5234
rect 12686 5182 12738 5234
rect 15598 5182 15650 5234
rect 18622 5238 18674 5290
rect 17166 5182 17218 5234
rect 21982 5182 22034 5234
rect 7646 5070 7698 5122
rect 7758 5070 7810 5122
rect 7926 5070 7978 5122
rect 9214 5070 9266 5122
rect 10670 5070 10722 5122
rect 11006 5070 11058 5122
rect 11566 5070 11618 5122
rect 11790 5070 11842 5122
rect 12238 5070 12290 5122
rect 12574 5055 12626 5107
rect 13694 5070 13746 5122
rect 13806 5070 13858 5122
rect 14030 5070 14082 5122
rect 15262 5070 15314 5122
rect 15486 5031 15538 5083
rect 15934 5070 15986 5122
rect 16830 5070 16882 5122
rect 17726 5070 17778 5122
rect 18062 5055 18114 5107
rect 18510 5070 18562 5122
rect 18846 5070 18898 5122
rect 19294 5070 19346 5122
rect 19574 5040 19626 5092
rect 20862 5070 20914 5122
rect 21590 5070 21642 5122
rect 22318 5070 22370 5122
rect 14310 4958 14362 5010
rect 17838 4902 17890 4954
rect 19630 4902 19682 4954
rect 6534 4678 6586 4730
rect 6638 4678 6690 4730
rect 6742 4678 6794 4730
rect 11854 4678 11906 4730
rect 11958 4678 12010 4730
rect 12062 4678 12114 4730
rect 17174 4678 17226 4730
rect 17278 4678 17330 4730
rect 17382 4678 17434 4730
rect 22494 4678 22546 4730
rect 22598 4678 22650 4730
rect 22702 4678 22754 4730
rect 4790 4510 4842 4562
rect 7758 4510 7810 4562
rect 8710 4510 8762 4562
rect 13638 4510 13690 4562
rect 14142 4510 14194 4562
rect 17446 4510 17498 4562
rect 19406 4510 19458 4562
rect 4174 4398 4226 4450
rect 3930 4342 3982 4394
rect 12014 4398 12066 4450
rect 20022 4398 20074 4450
rect 3054 4286 3106 4338
rect 8094 4286 8146 4338
rect 11622 4286 11674 4338
rect 12574 4342 12626 4394
rect 11846 4286 11898 4338
rect 12238 4286 12290 4338
rect 14478 4286 14530 4338
rect 17614 4286 17666 4338
rect 19742 4286 19794 4338
rect 20302 4286 20354 4338
rect 20526 4286 20578 4338
rect 20862 4286 20914 4338
rect 21198 4286 21250 4338
rect 20750 4118 20802 4170
rect 21702 4174 21754 4226
rect 22150 4174 22202 4226
rect 3874 3894 3926 3946
rect 3978 3894 4030 3946
rect 4082 3894 4134 3946
rect 9194 3894 9246 3946
rect 9298 3894 9350 3946
rect 9402 3894 9454 3946
rect 14514 3894 14566 3946
rect 14618 3894 14670 3946
rect 14722 3894 14774 3946
rect 19834 3894 19886 3946
rect 19938 3894 19990 3946
rect 20042 3894 20094 3946
rect 6534 3110 6586 3162
rect 6638 3110 6690 3162
rect 6742 3110 6794 3162
rect 11854 3110 11906 3162
rect 11958 3110 12010 3162
rect 12062 3110 12114 3162
rect 17174 3110 17226 3162
rect 17278 3110 17330 3162
rect 17382 3110 17434 3162
rect 22494 3110 22546 3162
rect 22598 3110 22650 3162
rect 22702 3110 22754 3162
<< metal2 >>
rect 1792 23200 1904 24000
rect 4032 23200 4144 24000
rect 6272 23200 6384 24000
rect 8512 23200 8624 24000
rect 8876 23212 9604 23268
rect 1820 20188 1876 23200
rect 4060 20188 4116 23200
rect 6300 20188 6356 23200
rect 8540 23044 8596 23200
rect 8876 23044 8932 23212
rect 8540 22988 8932 23044
rect 6532 20412 6796 20422
rect 6588 20356 6636 20412
rect 6692 20356 6740 20412
rect 6532 20346 6796 20356
rect 1820 20132 2212 20188
rect 4060 20132 4564 20188
rect 6300 20132 6804 20188
rect 2156 20130 2212 20132
rect 2156 20078 2158 20130
rect 2210 20078 2212 20130
rect 2156 20066 2212 20078
rect 4508 20130 4564 20132
rect 4508 20078 4510 20130
rect 4562 20078 4564 20130
rect 4508 20066 4564 20078
rect 6748 20130 6804 20132
rect 6748 20078 6750 20130
rect 6802 20078 6804 20130
rect 6748 20066 6804 20078
rect 9548 20130 9604 23212
rect 10752 23200 10864 24000
rect 12992 23200 13104 24000
rect 15232 23200 15344 24000
rect 17472 23200 17584 24000
rect 19712 23200 19824 24000
rect 21952 23200 22064 24000
rect 10780 20188 10836 23200
rect 11852 20412 12116 20422
rect 11908 20356 11956 20412
rect 12012 20356 12060 20412
rect 11852 20346 12116 20356
rect 13020 20188 13076 23200
rect 15260 20188 15316 23200
rect 17172 20412 17436 20422
rect 17228 20356 17276 20412
rect 17332 20356 17380 20412
rect 17172 20346 17436 20356
rect 17500 20188 17556 23200
rect 19740 20188 19796 23200
rect 20076 22036 20132 22046
rect 10780 20132 11284 20188
rect 13020 20132 13412 20188
rect 15260 20132 15764 20188
rect 17500 20132 18004 20188
rect 19740 20132 19908 20188
rect 9548 20078 9550 20130
rect 9602 20078 9604 20130
rect 9548 20066 9604 20078
rect 11228 20130 11284 20132
rect 11228 20078 11230 20130
rect 11282 20078 11284 20130
rect 11228 20066 11284 20078
rect 13356 20130 13412 20132
rect 13356 20078 13358 20130
rect 13410 20078 13412 20130
rect 13356 20066 13412 20078
rect 15708 20130 15764 20132
rect 15708 20078 15710 20130
rect 15762 20078 15764 20130
rect 15708 20066 15764 20078
rect 17948 20130 18004 20132
rect 17948 20078 17950 20130
rect 18002 20078 18004 20130
rect 17948 20066 18004 20078
rect 19852 20066 19908 20076
rect 20076 20130 20132 21980
rect 20076 20078 20078 20130
rect 20130 20078 20132 20130
rect 20076 20066 20132 20078
rect 20972 20132 21028 20142
rect 21980 20132 22036 23200
rect 22492 20412 22756 20422
rect 22548 20356 22596 20412
rect 22652 20356 22700 20412
rect 22492 20346 22756 20356
rect 22092 20132 22148 20142
rect 21980 20130 22148 20132
rect 21980 20078 22094 20130
rect 22146 20078 22148 20130
rect 21980 20076 22148 20078
rect 20972 20038 21028 20076
rect 22092 20066 22148 20076
rect 2492 20020 2548 20030
rect 4172 20020 4228 20030
rect 2492 20018 3108 20020
rect 2492 19966 2494 20018
rect 2546 19966 3108 20018
rect 2492 19964 3108 19966
rect 2492 19954 2548 19964
rect 3052 19458 3108 19964
rect 3052 19406 3054 19458
rect 3106 19406 3108 19458
rect 3052 19394 3108 19406
rect 3724 20018 4228 20020
rect 3724 19966 4174 20018
rect 4226 19966 4228 20018
rect 3724 19964 4228 19966
rect 3724 19458 3780 19964
rect 4172 19954 4228 19964
rect 5852 20020 5908 20030
rect 3872 19628 4136 19638
rect 3928 19572 3976 19628
rect 4032 19572 4080 19628
rect 3872 19562 4136 19572
rect 3724 19406 3726 19458
rect 3778 19406 3780 19458
rect 3724 19394 3780 19406
rect 4508 19460 4564 19470
rect 4508 19366 4564 19404
rect 5852 19458 5908 19964
rect 5852 19406 5854 19458
rect 5906 19406 5908 19458
rect 5852 19394 5908 19406
rect 6412 20018 6468 20030
rect 6412 19966 6414 20018
rect 6466 19966 6468 20018
rect 6412 19460 6468 19966
rect 9212 20020 9268 20030
rect 9212 19926 9268 19964
rect 10892 20018 10948 20030
rect 10892 19966 10894 20018
rect 10946 19966 10948 20018
rect 9192 19628 9456 19638
rect 9248 19572 9296 19628
rect 9352 19572 9400 19628
rect 9192 19562 9456 19572
rect 6412 19394 6468 19404
rect 10892 19458 10948 19966
rect 10892 19406 10894 19458
rect 10946 19406 10948 19458
rect 10892 19394 10948 19406
rect 13692 20018 13748 20030
rect 15372 20020 15428 20030
rect 13692 19966 13694 20018
rect 13746 19966 13748 20018
rect 3388 19236 3444 19246
rect 4060 19236 4116 19246
rect 3388 19234 3556 19236
rect 3388 19182 3390 19234
rect 3442 19182 3556 19234
rect 3388 19180 3556 19182
rect 3388 19170 3444 19180
rect 3388 18564 3444 18574
rect 3388 17666 3444 18508
rect 3500 18350 3556 19180
rect 4060 19142 4116 19180
rect 4172 19234 4228 19246
rect 4172 19182 4174 19234
rect 4226 19182 4228 19234
rect 3500 18338 3612 18350
rect 3500 18286 3558 18338
rect 3610 18286 3612 18338
rect 3500 18284 3612 18286
rect 3556 18004 3612 18284
rect 4172 18228 4228 19182
rect 5012 19236 5068 19246
rect 5012 19066 5068 19180
rect 5180 19236 5236 19246
rect 5180 19142 5236 19180
rect 5516 19234 5572 19246
rect 7980 19236 8036 19246
rect 5516 19182 5518 19234
rect 5570 19182 5572 19234
rect 5012 19014 5014 19066
rect 5066 19014 5068 19066
rect 5012 19002 5068 19014
rect 3556 17938 3612 17948
rect 3724 18172 4228 18228
rect 4508 18564 4564 18574
rect 3500 17834 3556 17846
rect 3500 17782 3502 17834
rect 3554 17782 3556 17834
rect 3500 17780 3556 17782
rect 3500 17714 3556 17724
rect 2712 17628 2768 17640
rect 2712 17576 2714 17628
rect 2766 17576 2768 17628
rect 3388 17614 3390 17666
rect 3442 17614 3444 17666
rect 3388 17602 3444 17614
rect 2712 17108 2768 17576
rect 3724 17108 3780 18172
rect 3872 18060 4136 18070
rect 3928 18004 3976 18060
rect 4032 18004 4080 18060
rect 3872 17994 4136 18004
rect 4508 17892 4564 18508
rect 5516 18564 5572 19182
rect 7420 19234 8372 19236
rect 7420 19182 7982 19234
rect 8034 19182 8372 19234
rect 7420 19180 8372 19182
rect 6532 18844 6796 18854
rect 6588 18788 6636 18844
rect 6692 18788 6740 18844
rect 6532 18778 6796 18788
rect 5516 18498 5572 18508
rect 7420 18450 7476 19180
rect 7980 19170 8036 19180
rect 7420 18398 7422 18450
rect 7474 18398 7476 18450
rect 7420 18386 7476 18398
rect 7644 18564 7700 18574
rect 7644 18465 7700 18508
rect 7644 18413 7646 18465
rect 7698 18413 7700 18465
rect 4172 17836 4564 17892
rect 3948 17780 4004 17790
rect 3948 17628 4004 17724
rect 3948 17576 3950 17628
rect 4002 17576 4004 17628
rect 3948 17564 4004 17576
rect 2712 17052 3108 17108
rect 2828 16658 2884 16670
rect 2828 16606 2830 16658
rect 2882 16606 2884 16658
rect 2828 15428 2884 16606
rect 3052 16324 3108 17052
rect 3612 17052 3780 17108
rect 3164 16884 3220 16894
rect 3444 16884 3500 16894
rect 3164 16882 3500 16884
rect 3164 16830 3166 16882
rect 3218 16830 3446 16882
rect 3498 16830 3500 16882
rect 3164 16828 3500 16830
rect 3164 16818 3220 16828
rect 3444 16818 3500 16828
rect 3612 16324 3668 17052
rect 3724 16884 3780 16894
rect 3724 16790 3780 16828
rect 3948 16882 4004 16894
rect 3948 16830 3950 16882
rect 4002 16830 4004 16882
rect 3948 16660 4004 16830
rect 4172 16882 4228 17836
rect 4508 17778 4564 17836
rect 7644 17780 7700 18413
rect 8092 18450 8148 18462
rect 8092 18398 8094 18450
rect 8146 18398 8148 18450
rect 7756 18340 7812 18350
rect 7756 18246 7812 18284
rect 4508 17726 4510 17778
rect 4562 17726 4564 17778
rect 4508 17714 4564 17726
rect 7532 17724 7700 17780
rect 4172 16830 4174 16882
rect 4226 16830 4228 16882
rect 4172 16818 4228 16830
rect 4284 17666 4340 17678
rect 4284 17614 4286 17666
rect 4338 17614 4340 17666
rect 4844 17668 4900 17678
rect 4284 16660 4340 17614
rect 4676 17610 4732 17622
rect 3948 16604 4340 16660
rect 3872 16492 4136 16502
rect 3928 16436 3976 16492
rect 4032 16436 4080 16492
rect 3872 16426 4136 16436
rect 3052 16268 3220 16324
rect 3612 16268 3780 16324
rect 2828 15362 2884 15372
rect 3164 16266 3220 16268
rect 3164 16214 3166 16266
rect 3218 16214 3220 16266
rect 3164 15316 3220 16214
rect 3388 16100 3444 16110
rect 3612 16100 3668 16110
rect 3388 16098 3612 16100
rect 3388 16046 3390 16098
rect 3442 16046 3612 16098
rect 3388 16044 3612 16046
rect 3388 16034 3444 16044
rect 3612 15482 3668 16044
rect 3612 15430 3614 15482
rect 3666 15430 3668 15482
rect 3612 15418 3668 15430
rect 3500 15316 3556 15326
rect 3164 15314 3556 15316
rect 3164 15262 3502 15314
rect 3554 15262 3556 15314
rect 3164 15260 3556 15262
rect 3500 15250 3556 15260
rect 3724 15148 3780 16268
rect 4284 16266 4340 16604
rect 4284 16214 4286 16266
rect 4338 16214 4340 16266
rect 4284 16202 4340 16214
rect 4508 17556 4564 17566
rect 4508 17108 4564 17500
rect 4676 17558 4678 17610
rect 4730 17558 4732 17610
rect 4676 17108 4732 17558
rect 4676 17052 4788 17108
rect 3948 16098 4004 16110
rect 3948 16046 3950 16098
rect 4002 16046 4004 16098
rect 3836 15428 3892 15438
rect 3836 15358 3892 15372
rect 3836 15306 3838 15358
rect 3890 15306 3892 15358
rect 3836 15294 3892 15306
rect 3948 15316 4004 16046
rect 4396 16100 4452 16110
rect 4396 16006 4452 16044
rect 3948 15250 4004 15260
rect 4508 15148 4564 17052
rect 4620 16098 4676 16110
rect 4620 16046 4622 16098
rect 4674 16046 4676 16098
rect 4620 15326 4676 16046
rect 4732 16100 4788 17052
rect 4844 16884 4900 17612
rect 6532 17276 6796 17286
rect 6588 17220 6636 17276
rect 6692 17220 6740 17276
rect 6532 17210 6796 17220
rect 4844 16790 4900 16828
rect 4732 16034 4788 16044
rect 4956 16714 5012 16726
rect 4956 16662 4958 16714
rect 5010 16662 5012 16714
rect 4620 15316 4732 15326
rect 4620 15260 4676 15316
rect 3500 15092 3780 15148
rect 4396 15092 4564 15148
rect 3500 12404 3556 15092
rect 3872 14924 4136 14934
rect 3928 14868 3976 14924
rect 4032 14868 4080 14924
rect 3872 14858 4136 14868
rect 4172 13860 4228 13870
rect 4172 13766 4228 13804
rect 3872 13356 4136 13366
rect 3928 13300 3976 13356
rect 4032 13300 4080 13356
rect 3872 13290 4136 13300
rect 4284 13076 4340 13086
rect 3500 12402 3668 12404
rect 3500 12350 3502 12402
rect 3554 12350 3668 12402
rect 3500 12348 3668 12350
rect 3500 12338 3556 12348
rect 3164 12180 3220 12190
rect 2922 12178 3220 12180
rect 2922 12126 3166 12178
rect 3218 12126 3220 12178
rect 2922 12124 3220 12126
rect 2922 11618 2978 12124
rect 3164 12114 3220 12124
rect 3612 11732 3668 12348
rect 3872 11788 4136 11798
rect 3928 11732 3976 11788
rect 4032 11732 4080 11788
rect 3612 11676 3724 11732
rect 3872 11722 4136 11732
rect 2922 11566 2924 11618
rect 2976 11566 2978 11618
rect 2922 11554 2978 11566
rect 3668 11450 3724 11676
rect 3164 11396 3220 11406
rect 3164 11302 3220 11340
rect 3668 11398 3670 11450
rect 3722 11398 3724 11450
rect 3668 10836 3724 11398
rect 3948 11396 4004 11406
rect 3388 10780 3724 10836
rect 3836 11282 3892 11294
rect 3836 11230 3838 11282
rect 3890 11230 3892 11282
rect 3388 8260 3444 10780
rect 3556 10666 3612 10678
rect 3556 10614 3558 10666
rect 3610 10614 3612 10666
rect 3556 10612 3612 10614
rect 3724 10612 3780 10622
rect 3836 10612 3892 11230
rect 3948 10722 4004 11340
rect 4284 11394 4340 13020
rect 4396 12852 4452 15092
rect 4676 14754 4732 15260
rect 4956 15148 5012 16662
rect 7532 16714 7588 17724
rect 7980 16996 8036 17006
rect 7532 16662 7534 16714
rect 7586 16662 7588 16714
rect 7532 16650 7588 16662
rect 7644 16882 7700 16894
rect 7644 16830 7646 16882
rect 7698 16830 7700 16882
rect 7532 16100 7588 16110
rect 6532 15708 6796 15718
rect 6588 15652 6636 15708
rect 6692 15652 6740 15708
rect 6532 15642 6796 15652
rect 7532 15148 7588 16044
rect 4676 14702 4678 14754
rect 4730 14702 4732 14754
rect 4676 14690 4732 14702
rect 4844 15092 5012 15148
rect 7196 15092 7588 15148
rect 4620 14308 4676 14318
rect 4508 13746 4564 13758
rect 4508 13694 4510 13746
rect 4562 13694 4564 13746
rect 4508 13076 4564 13694
rect 4620 13746 4676 14252
rect 4844 13972 4900 15092
rect 5180 14644 5236 14654
rect 4620 13694 4622 13746
rect 4674 13694 4676 13746
rect 4620 13682 4676 13694
rect 4732 13916 4900 13972
rect 4956 14530 5012 14542
rect 4956 14478 4958 14530
rect 5010 14478 5012 14530
rect 4508 13010 4564 13020
rect 4396 12796 4676 12852
rect 4284 11342 4286 11394
rect 4338 11342 4340 11394
rect 4284 11330 4340 11342
rect 4396 11954 4452 11966
rect 4396 11902 4398 11954
rect 4450 11902 4452 11954
rect 4284 11226 4340 11238
rect 4284 11174 4286 11226
rect 4338 11174 4340 11226
rect 4284 10948 4340 11174
rect 3948 10670 3950 10722
rect 4002 10670 4004 10722
rect 3948 10658 4004 10670
rect 4116 10892 4340 10948
rect 4116 10666 4172 10892
rect 3556 10556 3668 10612
rect 3612 8484 3668 10556
rect 3724 10610 3892 10612
rect 3724 10558 3726 10610
rect 3778 10558 3892 10610
rect 4116 10614 4118 10666
rect 4170 10614 4172 10666
rect 4116 10602 4172 10614
rect 3724 10556 3892 10558
rect 3724 9940 3780 10556
rect 3872 10220 4136 10230
rect 3928 10164 3976 10220
rect 4032 10164 4080 10220
rect 3872 10154 4136 10164
rect 4396 9940 4452 11902
rect 4508 11396 4564 11406
rect 4508 11315 4510 11340
rect 4562 11315 4564 11340
rect 4508 11302 4564 11315
rect 4620 10052 4676 12796
rect 3724 9874 3780 9884
rect 4228 9884 4452 9940
rect 4508 9996 4676 10052
rect 4228 9882 4340 9884
rect 4228 9830 4230 9882
rect 4282 9830 4340 9882
rect 4228 9818 4340 9830
rect 3872 8652 4136 8662
rect 3928 8596 3976 8652
rect 4032 8596 4080 8652
rect 3872 8586 4136 8596
rect 3948 8484 4004 8494
rect 3612 8482 4004 8484
rect 3612 8430 3950 8482
rect 4002 8430 4004 8482
rect 3612 8428 4004 8430
rect 3948 8418 4004 8428
rect 4284 8372 4340 9818
rect 4396 9716 4452 9726
rect 4396 9622 4452 9660
rect 4508 8596 4564 9996
rect 4620 9826 4676 9838
rect 4620 9774 4622 9826
rect 4674 9774 4676 9826
rect 4620 9044 4676 9774
rect 4732 9828 4788 13916
rect 4844 13748 4900 13758
rect 4844 13654 4900 13692
rect 4844 12738 4900 12750
rect 4844 12686 4846 12738
rect 4898 12686 4900 12738
rect 4844 11954 4900 12686
rect 4844 11902 4846 11954
rect 4898 11902 4900 11954
rect 4844 11890 4900 11902
rect 4844 11394 4900 11406
rect 4844 11342 4846 11394
rect 4898 11342 4900 11394
rect 4844 9940 4900 11342
rect 4844 9874 4900 9884
rect 4732 9268 4788 9772
rect 4956 9770 5012 14478
rect 5180 14530 5236 14588
rect 5796 14644 5852 14654
rect 5796 14550 5852 14588
rect 5180 14478 5182 14530
rect 5234 14478 5236 14530
rect 5180 14466 5236 14478
rect 5684 14308 5740 14318
rect 5684 13972 5740 14252
rect 6532 14140 6796 14150
rect 6588 14084 6636 14140
rect 6692 14084 6740 14140
rect 6532 14074 6796 14084
rect 5684 13970 5908 13972
rect 5684 13918 5686 13970
rect 5738 13918 5908 13970
rect 5684 13916 5908 13918
rect 5684 13906 5740 13916
rect 5124 13522 5180 13534
rect 5124 13470 5126 13522
rect 5178 13470 5180 13522
rect 5124 12974 5180 13470
rect 5124 12962 5236 12974
rect 5124 12910 5182 12962
rect 5234 12910 5236 12962
rect 5124 12908 5236 12910
rect 5180 12898 5236 12908
rect 4956 9718 4958 9770
rect 5010 9718 5012 9770
rect 4956 9268 5012 9718
rect 5740 9770 5796 9782
rect 5740 9718 5742 9770
rect 5794 9718 5796 9770
rect 5740 9268 5796 9718
rect 4732 9212 4900 9268
rect 4732 9044 4788 9054
rect 4620 9042 4788 9044
rect 4620 8990 4734 9042
rect 4786 8990 4788 9042
rect 4620 8988 4788 8990
rect 4732 8932 4788 8988
rect 4732 8866 4788 8876
rect 4508 8540 4788 8596
rect 4060 8316 4340 8372
rect 4508 8372 4564 8382
rect 3500 8260 3556 8270
rect 3388 8258 3556 8260
rect 3388 8206 3502 8258
rect 3554 8206 3556 8258
rect 3388 8204 3556 8206
rect 3500 8194 3556 8204
rect 3332 8036 3388 8046
rect 3332 8034 3444 8036
rect 3332 7982 3334 8034
rect 3386 7982 3444 8034
rect 3332 7970 3444 7982
rect 3388 7504 3444 7970
rect 3892 7700 3948 7710
rect 3892 7530 3948 7644
rect 3388 7452 3390 7504
rect 3442 7452 3444 7504
rect 3388 5460 3444 7452
rect 3612 7513 3668 7525
rect 3612 7461 3614 7513
rect 3666 7461 3668 7513
rect 3892 7478 3894 7530
rect 3946 7478 3948 7530
rect 3892 7466 3948 7478
rect 3612 6018 3668 7461
rect 4060 7252 4116 8316
rect 4508 8258 4564 8316
rect 4340 8202 4396 8214
rect 4340 8150 4342 8202
rect 4394 8150 4396 8202
rect 4508 8206 4510 8258
rect 4562 8206 4564 8258
rect 4508 8194 4564 8206
rect 4620 8260 4676 8270
rect 4620 8166 4676 8204
rect 4340 7700 4396 8150
rect 4732 7924 4788 8540
rect 4172 7644 4396 7700
rect 4508 7868 4788 7924
rect 4172 7586 4228 7644
rect 4172 7534 4174 7586
rect 4226 7534 4228 7586
rect 4172 7522 4228 7534
rect 4508 7476 4564 7868
rect 4676 7700 4732 7710
rect 4676 7606 4732 7644
rect 4508 7382 4564 7420
rect 3724 7196 4116 7252
rect 3724 6580 3780 7196
rect 3872 7084 4136 7094
rect 3928 7028 3976 7084
rect 4032 7028 4080 7084
rect 3872 7018 4136 7028
rect 3724 6524 3911 6580
rect 3612 5966 3614 6018
rect 3666 5966 3668 6018
rect 3612 5572 3668 5966
rect 3855 5962 3911 6524
rect 3855 5910 3857 5962
rect 3909 5910 3911 5962
rect 3855 5908 3911 5910
rect 3855 5832 3911 5852
rect 4732 5908 4788 5918
rect 4844 5908 4900 9212
rect 4956 9202 5012 9212
rect 5180 9212 5796 9268
rect 5068 9042 5124 9054
rect 5068 8990 5070 9042
rect 5122 8990 5124 9042
rect 5068 8382 5124 8990
rect 5180 8874 5236 9212
rect 5180 8822 5182 8874
rect 5234 8822 5236 8874
rect 5180 8810 5236 8822
rect 5684 8930 5740 8942
rect 5684 8878 5686 8930
rect 5738 8878 5740 8930
rect 5068 8372 5180 8382
rect 5068 8316 5124 8372
rect 5124 8278 5180 8316
rect 5684 8372 5740 8878
rect 5852 8382 5908 13916
rect 7196 13860 7252 15092
rect 7644 14084 7700 16830
rect 7980 16882 8036 16940
rect 7980 16830 7982 16882
rect 8034 16830 8036 16882
rect 7980 14644 8036 16830
rect 8092 16100 8148 18398
rect 8316 17890 8372 19180
rect 8652 19234 8708 19246
rect 9100 19236 9156 19246
rect 11228 19236 11284 19246
rect 8652 19182 8654 19234
rect 8706 19182 8708 19234
rect 8316 17838 8318 17890
rect 8370 17838 8372 17890
rect 8316 17826 8372 17838
rect 8540 19066 8596 19078
rect 8540 19014 8542 19066
rect 8594 19014 8596 19066
rect 8540 18506 8596 19014
rect 8540 18454 8542 18506
rect 8594 18454 8596 18506
rect 8652 18564 8708 19182
rect 8876 19234 9156 19236
rect 8876 19182 9102 19234
rect 9154 19182 9156 19234
rect 8876 19180 9156 19182
rect 8876 18618 8932 19180
rect 9100 19170 9156 19180
rect 11004 19234 11284 19236
rect 11004 19182 11230 19234
rect 11282 19182 11284 19234
rect 11004 19180 11284 19182
rect 8876 18566 8878 18618
rect 8930 18566 8932 18618
rect 8876 18554 8932 18566
rect 9436 19010 9492 19022
rect 9436 18958 9438 19010
rect 9490 18958 9492 19010
rect 9436 18564 9492 18958
rect 11004 18674 11060 19180
rect 11228 19170 11284 19180
rect 11852 18844 12116 18854
rect 11908 18788 11956 18844
rect 12012 18788 12060 18844
rect 11852 18778 12116 18788
rect 11004 18622 11006 18674
rect 11058 18622 11060 18674
rect 11004 18610 11060 18622
rect 8652 18498 8708 18508
rect 9436 18498 9492 18508
rect 9660 18465 9716 18477
rect 8540 17668 8596 18454
rect 8764 18450 8820 18462
rect 8764 18398 8766 18450
rect 8818 18398 8820 18450
rect 8764 18340 8820 18398
rect 9660 18413 9662 18465
rect 9714 18413 9716 18465
rect 9548 18340 9604 18350
rect 8764 18338 9604 18340
rect 8764 18286 9550 18338
rect 9602 18286 9604 18338
rect 8764 18284 9604 18286
rect 9548 18274 9604 18284
rect 9660 18340 9716 18413
rect 9996 18452 10052 18462
rect 9996 18358 10052 18396
rect 10668 18452 10724 18462
rect 10668 18450 10836 18452
rect 10668 18398 10670 18450
rect 10722 18398 10836 18450
rect 10668 18396 10836 18398
rect 10668 18386 10724 18396
rect 9192 18060 9456 18070
rect 9248 18004 9296 18060
rect 9352 18004 9400 18060
rect 9192 17994 9456 18004
rect 9380 17834 9436 17846
rect 9380 17782 9382 17834
rect 9434 17782 9436 17834
rect 8708 17668 8764 17678
rect 8540 17666 8764 17668
rect 8540 17614 8710 17666
rect 8762 17614 8764 17666
rect 8540 17612 8764 17614
rect 8708 17602 8764 17612
rect 8876 17668 8932 17678
rect 8484 17444 8540 17454
rect 8484 17106 8540 17388
rect 8484 17054 8486 17106
rect 8538 17054 8540 17106
rect 8484 16996 8540 17054
rect 8484 16930 8540 16940
rect 8876 16996 8932 17612
rect 8988 17668 9044 17678
rect 9380 17668 9436 17782
rect 8988 17666 9436 17668
rect 8988 17614 8990 17666
rect 9042 17614 9436 17666
rect 8988 17612 9436 17614
rect 9548 17668 9604 17678
rect 9660 17668 9716 18284
rect 9548 17666 9716 17668
rect 9548 17614 9550 17666
rect 9602 17614 9716 17666
rect 9548 17612 9716 17614
rect 8988 17602 9044 17612
rect 9548 17602 9604 17612
rect 10780 17006 10836 18396
rect 13692 18340 13748 19966
rect 15148 20018 15428 20020
rect 15148 19966 15374 20018
rect 15426 19966 15428 20018
rect 15148 19964 15428 19966
rect 14512 19628 14776 19638
rect 14568 19572 14616 19628
rect 14672 19572 14720 19628
rect 14512 19562 14776 19572
rect 15148 19458 15204 19964
rect 15372 19954 15428 19964
rect 17612 20018 17668 20030
rect 19740 20020 19796 20030
rect 17612 19966 17614 20018
rect 17666 19966 17668 20018
rect 14252 19402 14308 19414
rect 14252 19350 14254 19402
rect 14306 19350 14308 19402
rect 15148 19406 15150 19458
rect 15202 19406 15204 19458
rect 15148 19394 15204 19406
rect 16380 19460 16436 19470
rect 16380 19366 16436 19404
rect 17612 19460 17668 19966
rect 19628 20018 19796 20020
rect 19628 19966 19742 20018
rect 19794 19966 19796 20018
rect 19628 19964 19796 19966
rect 17612 19394 17668 19404
rect 18620 19460 18676 19470
rect 18620 19366 18676 19404
rect 14140 19234 14196 19246
rect 14140 19182 14142 19234
rect 14194 19182 14196 19234
rect 14140 19012 14196 19182
rect 14252 19236 14308 19350
rect 14252 19170 14308 19180
rect 14476 19234 14532 19246
rect 14476 19182 14478 19234
rect 14530 19182 14532 19234
rect 14140 18946 14196 18956
rect 14476 18574 14532 19182
rect 14812 19236 14868 19246
rect 14812 19234 15092 19236
rect 14812 19182 14814 19234
rect 14866 19182 15092 19234
rect 14812 19180 15092 19182
rect 14812 19170 14868 19180
rect 14420 18562 14532 18574
rect 14420 18510 14422 18562
rect 14474 18510 14532 18562
rect 14420 18508 14532 18510
rect 14924 19012 14980 19022
rect 14420 18498 14476 18508
rect 14028 18452 14084 18462
rect 14028 18358 14084 18396
rect 14140 18452 14196 18462
rect 14140 18450 14308 18452
rect 14140 18398 14142 18450
rect 14194 18398 14308 18450
rect 14140 18396 14308 18398
rect 14140 18386 14196 18396
rect 13692 18274 13748 18284
rect 13860 18228 13916 18238
rect 13860 17890 13916 18172
rect 14252 18004 14308 18396
rect 14700 18450 14756 18462
rect 14700 18398 14702 18450
rect 14754 18398 14756 18450
rect 14700 18228 14756 18398
rect 14700 18162 14756 18172
rect 14512 18060 14776 18070
rect 14568 18004 14616 18060
rect 14672 18004 14720 18060
rect 14252 17948 14420 18004
rect 14512 17994 14776 18004
rect 13860 17838 13862 17890
rect 13914 17838 13916 17890
rect 13860 17826 13916 17838
rect 14364 17892 14420 17948
rect 14644 17892 14700 17902
rect 14364 17890 14700 17892
rect 14364 17838 14646 17890
rect 14698 17838 14700 17890
rect 14364 17836 14700 17838
rect 14644 17826 14700 17836
rect 12684 17668 12740 17678
rect 11508 17442 11564 17454
rect 11508 17390 11510 17442
rect 11562 17390 11564 17442
rect 11508 17108 11564 17390
rect 11852 17276 12116 17286
rect 11908 17220 11956 17276
rect 12012 17220 12060 17276
rect 11852 17210 12116 17220
rect 11116 17052 11564 17108
rect 11676 17108 11732 17118
rect 10780 16994 10892 17006
rect 10780 16942 10838 16994
rect 10890 16942 10892 16994
rect 10780 16940 10892 16942
rect 8876 16930 8932 16940
rect 10836 16930 10892 16940
rect 11116 16882 11172 17052
rect 11116 16830 11118 16882
rect 11170 16830 11172 16882
rect 9192 16492 9456 16502
rect 9248 16436 9296 16492
rect 9352 16436 9400 16492
rect 9192 16426 9456 16436
rect 8092 16034 8148 16044
rect 9192 14924 9456 14934
rect 9248 14868 9296 14924
rect 9352 14868 9400 14924
rect 9192 14858 9456 14868
rect 7980 14578 8036 14588
rect 8652 14532 8708 14542
rect 8540 14530 9044 14532
rect 8540 14478 8654 14530
rect 8706 14478 9044 14530
rect 8540 14476 9044 14478
rect 7196 13794 7252 13804
rect 7308 14028 7700 14084
rect 8316 14306 8372 14318
rect 8316 14254 8318 14306
rect 8370 14254 8372 14306
rect 7308 13748 7364 14028
rect 8092 13860 8148 13870
rect 7308 13634 7364 13692
rect 7308 13582 7310 13634
rect 7362 13582 7364 13634
rect 7308 13570 7364 13582
rect 7420 13761 7476 13773
rect 7420 13709 7422 13761
rect 7474 13709 7476 13761
rect 7420 13524 7476 13709
rect 7756 13748 7812 13758
rect 7756 13746 7924 13748
rect 7756 13694 7758 13746
rect 7810 13694 7924 13746
rect 7756 13692 7924 13694
rect 7756 13682 7812 13692
rect 7420 13458 7476 13468
rect 7868 13188 7924 13692
rect 8092 13746 8148 13804
rect 8092 13694 8094 13746
rect 8146 13694 8148 13746
rect 8092 13682 8148 13694
rect 7420 13074 7476 13086
rect 7420 13022 7422 13074
rect 7474 13022 7476 13074
rect 6532 12572 6796 12582
rect 6588 12516 6636 12572
rect 6692 12516 6740 12572
rect 6532 12506 6796 12516
rect 6532 11004 6796 11014
rect 6588 10948 6636 11004
rect 6692 10948 6740 11004
rect 6532 10938 6796 10948
rect 6300 9940 6356 9950
rect 6300 9846 6356 9884
rect 6076 9826 6132 9838
rect 6076 9774 6078 9826
rect 6130 9774 6132 9826
rect 6076 9716 6132 9774
rect 6076 9044 6132 9660
rect 6468 9770 6524 9782
rect 6468 9718 6470 9770
rect 6522 9718 6524 9770
rect 6468 9716 6524 9718
rect 6468 9650 6524 9660
rect 6916 9716 6972 9726
rect 6916 9622 6972 9660
rect 6532 9436 6796 9446
rect 6588 9380 6636 9436
rect 6692 9380 6740 9436
rect 6532 9370 6796 9380
rect 6076 8978 6132 8988
rect 6972 9268 7028 9278
rect 7420 9268 7476 13022
rect 7868 12962 7924 13132
rect 8316 13188 8372 14254
rect 8316 13122 8372 13132
rect 8428 13773 8484 13785
rect 8428 13721 8430 13773
rect 8482 13721 8484 13773
rect 7532 12918 7588 12930
rect 7532 12866 7534 12918
rect 7586 12866 7588 12918
rect 7868 12910 7870 12962
rect 7922 12910 7924 12962
rect 7868 12898 7924 12910
rect 7532 12180 7588 12866
rect 8428 12404 8484 13721
rect 8540 12962 8596 14476
rect 8652 14466 8708 14476
rect 8988 14306 9044 14476
rect 8988 14254 8990 14306
rect 9042 14254 9044 14306
rect 8988 14242 9044 14254
rect 9772 14306 9828 14318
rect 9772 14254 9774 14306
rect 9826 14254 9828 14306
rect 9772 13970 9828 14254
rect 11116 13972 11172 16830
rect 11340 16884 11396 16894
rect 11340 16790 11396 16828
rect 11676 16222 11732 17052
rect 12236 17108 12292 17118
rect 12236 16938 12292 17052
rect 12012 16915 12068 16927
rect 12012 16884 12014 16915
rect 12066 16884 12068 16915
rect 12236 16886 12238 16938
rect 12290 16886 12292 16938
rect 12236 16874 12292 16886
rect 12684 16915 12740 17612
rect 13356 17666 13412 17678
rect 13356 17614 13358 17666
rect 13410 17614 13412 17666
rect 12964 17444 13020 17454
rect 13356 17444 13412 17614
rect 13580 17668 13636 17678
rect 13580 17574 13636 17612
rect 14252 17666 14308 17678
rect 14252 17614 14254 17666
rect 14306 17614 14308 17666
rect 12964 17442 13412 17444
rect 12964 17390 12966 17442
rect 13018 17390 13412 17442
rect 12964 17388 13412 17390
rect 12964 17378 13020 17388
rect 13132 16996 13188 17006
rect 12012 16818 12068 16828
rect 12684 16863 12686 16915
rect 12738 16863 12740 16915
rect 12994 16915 13050 16927
rect 11620 16210 11732 16222
rect 11620 16158 11622 16210
rect 11674 16158 11732 16210
rect 11620 16156 11732 16158
rect 11620 16146 11676 16156
rect 11852 15708 12116 15718
rect 11908 15652 11956 15708
rect 12012 15652 12060 15708
rect 11852 15642 12116 15652
rect 12684 15482 12740 16863
rect 12796 16884 12852 16894
rect 12796 16212 12852 16828
rect 12994 16863 12996 16915
rect 13048 16863 13050 16915
rect 13132 16902 13188 16940
rect 12994 16324 13050 16863
rect 12994 16268 13188 16324
rect 12796 16156 12964 16212
rect 12684 15430 12686 15482
rect 12738 15430 12740 15482
rect 12684 15418 12740 15430
rect 12572 15353 12628 15365
rect 12236 15314 12292 15326
rect 12236 15262 12238 15314
rect 12290 15262 12292 15314
rect 11852 14140 12116 14150
rect 11908 14084 11956 14140
rect 12012 14084 12060 14140
rect 11852 14074 12116 14084
rect 8876 13914 8932 13926
rect 8876 13862 8878 13914
rect 8930 13862 8932 13914
rect 9772 13918 9774 13970
rect 9826 13918 9828 13970
rect 9772 13906 9828 13918
rect 10892 13916 11116 13972
rect 8764 13748 8820 13758
rect 8876 13748 8932 13862
rect 9436 13748 9492 13758
rect 8876 13746 9492 13748
rect 8876 13694 9438 13746
rect 9490 13694 9492 13746
rect 8876 13692 9492 13694
rect 8764 13654 8820 13692
rect 9436 13682 9492 13692
rect 9996 13524 10052 13534
rect 9192 13356 9456 13366
rect 9248 13300 9296 13356
rect 9352 13300 9400 13356
rect 9192 13290 9456 13300
rect 8540 12910 8542 12962
rect 8594 12910 8596 12962
rect 8876 13074 8932 13086
rect 8876 13022 8878 13074
rect 8930 13022 8932 13074
rect 8540 12898 8596 12910
rect 8764 12918 8820 12930
rect 8428 12338 8484 12348
rect 8764 12866 8766 12918
rect 8818 12866 8820 12918
rect 8764 12292 8820 12866
rect 8876 12740 8932 13022
rect 9884 12852 9940 12862
rect 8876 12674 8932 12684
rect 9772 12740 9828 12750
rect 8764 12226 8820 12236
rect 8876 12404 8932 12414
rect 7532 12114 7588 12124
rect 8652 12193 8708 12218
rect 8652 12180 8654 12193
rect 8706 12180 8708 12193
rect 8652 12114 8708 12124
rect 8876 12178 8932 12348
rect 8876 12126 8878 12178
rect 8930 12126 8932 12178
rect 8876 12114 8932 12126
rect 8540 12066 8596 12078
rect 8540 12014 8542 12066
rect 8594 12014 8596 12066
rect 8540 10052 8596 12014
rect 9604 11956 9660 11966
rect 9548 11954 9660 11956
rect 9548 11902 9606 11954
rect 9658 11902 9660 11954
rect 9548 11890 9660 11902
rect 9192 11788 9456 11798
rect 9248 11732 9296 11788
rect 9352 11732 9400 11788
rect 9192 11722 9456 11732
rect 9192 10220 9456 10230
rect 9248 10164 9296 10220
rect 9352 10164 9400 10220
rect 9192 10154 9456 10164
rect 8540 9996 8708 10052
rect 8204 9828 8260 9838
rect 7028 9212 7476 9268
rect 7980 9716 8036 9726
rect 5684 8306 5740 8316
rect 5796 8370 5908 8382
rect 5796 8318 5798 8370
rect 5850 8318 5908 8370
rect 5796 8316 5908 8318
rect 5796 8260 5852 8316
rect 5796 8194 5852 8204
rect 6532 7868 6796 7878
rect 6588 7812 6636 7868
rect 6692 7812 6740 7868
rect 6532 7802 6796 7812
rect 4732 5906 4900 5908
rect 4732 5854 4734 5906
rect 4786 5854 4900 5906
rect 4732 5852 4900 5854
rect 4956 7476 5012 7486
rect 4732 5842 4788 5852
rect 3612 5506 3668 5516
rect 3872 5516 4136 5526
rect 3276 5404 3444 5460
rect 3928 5460 3976 5516
rect 4032 5460 4080 5516
rect 3872 5450 4136 5460
rect 3276 5124 3332 5404
rect 3500 5124 3556 5134
rect 3276 5122 3556 5124
rect 3276 5070 3502 5122
rect 3554 5070 3556 5122
rect 3276 5068 3556 5070
rect 3500 5058 3556 5068
rect 3612 5124 3668 5134
rect 4620 5124 4676 5134
rect 3052 4900 3108 4910
rect 3052 4338 3108 4844
rect 3612 4788 3668 5068
rect 4376 5066 4432 5078
rect 4376 5014 4378 5066
rect 4430 5014 4432 5066
rect 4620 5030 4676 5068
rect 3612 4732 3984 4788
rect 3052 4286 3054 4338
rect 3106 4286 3108 4338
rect 3928 4394 3984 4732
rect 3928 4342 3930 4394
rect 3982 4342 3984 4394
rect 4172 4452 4228 4462
rect 4376 4452 4432 5014
rect 4956 4900 5012 7420
rect 5236 7476 5292 7486
rect 5236 7382 5292 7420
rect 6532 6300 6796 6310
rect 6588 6244 6636 6300
rect 6692 6244 6740 6300
rect 6532 6234 6796 6244
rect 6804 5908 6860 5918
rect 6804 5814 6860 5852
rect 6972 5906 7028 9212
rect 7420 9044 7476 9054
rect 7420 8950 7476 8988
rect 7756 9042 7812 9054
rect 7756 8990 7758 9042
rect 7810 8990 7812 9042
rect 7420 8372 7476 8382
rect 7196 8260 7252 8270
rect 6972 5854 6974 5906
rect 7026 5854 7028 5906
rect 6972 5842 7028 5854
rect 7084 5908 7140 5918
rect 7084 5814 7140 5852
rect 6412 5684 6468 5694
rect 6412 5682 6580 5684
rect 6412 5630 6414 5682
rect 6466 5630 6580 5682
rect 6412 5628 6580 5630
rect 6412 5618 6468 5628
rect 6524 5178 6580 5628
rect 7196 5348 7252 8204
rect 7420 5796 7476 8316
rect 7644 7700 7700 7710
rect 7644 7252 7700 7644
rect 7588 7196 7700 7252
rect 7588 6746 7644 7196
rect 7588 6694 7590 6746
rect 7642 6694 7644 6746
rect 7588 6682 7644 6694
rect 7756 6690 7812 8990
rect 7868 9044 7924 9054
rect 7868 8874 7924 8988
rect 7868 8822 7870 8874
rect 7922 8822 7924 8874
rect 7868 8810 7924 8822
rect 7980 6916 8036 9660
rect 8204 9156 8260 9772
rect 8372 9604 8428 9614
rect 8372 9602 8596 9604
rect 8372 9550 8374 9602
rect 8426 9550 8596 9602
rect 8372 9548 8596 9550
rect 8372 9538 8428 9548
rect 8428 9380 8484 9390
rect 8204 9100 8372 9156
rect 8204 8932 8260 8942
rect 8204 8370 8260 8876
rect 8204 8318 8206 8370
rect 8258 8318 8260 8370
rect 8204 8306 8260 8318
rect 7756 6638 7758 6690
rect 7810 6638 7812 6690
rect 7756 6626 7812 6638
rect 7868 6860 8036 6916
rect 7868 5908 7924 6860
rect 7980 6692 8036 6702
rect 8204 6692 8260 6702
rect 7980 6690 8148 6692
rect 7980 6638 7982 6690
rect 8034 6638 8148 6690
rect 7980 6636 8148 6638
rect 7980 6626 8036 6636
rect 7980 6356 8036 6366
rect 7980 6020 8036 6300
rect 8092 6132 8148 6636
rect 8204 6610 8206 6636
rect 8258 6610 8260 6636
rect 8204 6356 8260 6610
rect 8316 6468 8372 9100
rect 8428 9070 8484 9324
rect 8428 9018 8430 9070
rect 8482 9018 8484 9070
rect 8428 8820 8484 9018
rect 8428 8754 8484 8764
rect 8540 9156 8596 9548
rect 8652 9380 8708 9996
rect 8652 9314 8708 9324
rect 8764 9826 8820 9838
rect 8764 9774 8766 9826
rect 8818 9774 8820 9826
rect 8540 8484 8596 9100
rect 8652 9044 8708 9054
rect 8764 9044 8820 9774
rect 9436 9828 9492 9838
rect 9548 9828 9604 11890
rect 9436 9826 9604 9828
rect 9436 9774 9438 9826
rect 9490 9774 9604 9826
rect 9436 9772 9604 9774
rect 9436 9762 9492 9772
rect 9548 9658 9604 9670
rect 9548 9606 9550 9658
rect 9602 9606 9604 9658
rect 9548 9154 9604 9606
rect 9548 9102 9550 9154
rect 9602 9102 9604 9154
rect 9548 9090 9604 9102
rect 9772 9156 9828 12684
rect 9884 12180 9940 12796
rect 9996 12290 10052 13468
rect 9996 12238 9998 12290
rect 10050 12238 10052 12290
rect 9996 12226 10052 12238
rect 10332 12404 10388 12414
rect 9884 12086 9940 12124
rect 10164 12180 10220 12190
rect 10164 12086 10220 12124
rect 10332 12178 10388 12348
rect 10332 12126 10334 12178
rect 10386 12126 10388 12178
rect 10332 12114 10388 12126
rect 10780 9156 10836 9166
rect 9772 9100 10052 9156
rect 8652 9042 8820 9044
rect 8652 8990 8654 9042
rect 8706 8990 8820 9042
rect 8652 8988 8820 8990
rect 8652 8932 8708 8988
rect 9044 8986 9100 8998
rect 8652 8866 8708 8876
rect 8876 8930 8932 8942
rect 8876 8878 8878 8930
rect 8930 8878 8932 8930
rect 8540 8418 8596 8428
rect 8540 8260 8596 8270
rect 8876 8260 8932 8878
rect 9044 8934 9046 8986
rect 9098 8934 9100 8986
rect 9044 8932 9100 8934
rect 9044 8866 9100 8876
rect 9716 8986 9772 8998
rect 9716 8934 9718 8986
rect 9770 8934 9772 8986
rect 9192 8652 9456 8662
rect 9248 8596 9296 8652
rect 9352 8596 9400 8652
rect 9192 8586 9456 8596
rect 9324 8484 9380 8494
rect 9548 8484 9604 8494
rect 9380 8428 9492 8484
rect 9324 8418 9380 8428
rect 9100 8260 9156 8270
rect 8540 8258 8708 8260
rect 8540 8206 8542 8258
rect 8594 8206 8708 8258
rect 8540 8204 8708 8206
rect 8876 8258 9156 8260
rect 8876 8206 9102 8258
rect 9154 8206 9156 8258
rect 9436 8258 9492 8428
rect 8876 8204 9156 8206
rect 8540 8194 8596 8204
rect 8316 6412 8428 6468
rect 8204 6290 8260 6300
rect 8092 6076 8260 6132
rect 7980 5964 8148 6020
rect 7868 5852 8036 5908
rect 7420 5740 7588 5796
rect 7308 5684 7364 5694
rect 7364 5628 7420 5684
rect 7308 5618 7420 5628
rect 6524 5126 6526 5178
rect 6578 5126 6580 5178
rect 7084 5292 7252 5348
rect 6524 5114 6580 5126
rect 6748 5124 6804 5134
rect 6748 5042 6750 5068
rect 6802 5042 6804 5068
rect 6748 5030 6804 5042
rect 4788 4564 4844 4574
rect 4956 4564 5012 4844
rect 6532 4732 6796 4742
rect 6588 4676 6636 4732
rect 6692 4676 6740 4732
rect 6532 4666 6796 4676
rect 4788 4562 5012 4564
rect 4788 4510 4790 4562
rect 4842 4510 5012 4562
rect 4788 4508 5012 4510
rect 7084 4564 7140 5292
rect 7364 5178 7420 5618
rect 7532 5460 7588 5740
rect 7812 5684 7868 5694
rect 7812 5590 7868 5628
rect 7532 5404 7812 5460
rect 7196 5124 7252 5134
rect 7364 5126 7366 5178
rect 7418 5126 7420 5178
rect 7364 5114 7420 5126
rect 7644 5236 7700 5246
rect 7644 5122 7700 5180
rect 7196 5030 7252 5068
rect 7644 5070 7646 5122
rect 7698 5070 7700 5122
rect 7644 5058 7700 5070
rect 7756 5122 7812 5404
rect 7980 5348 8036 5852
rect 8092 5906 8148 5964
rect 8092 5854 8094 5906
rect 8146 5854 8148 5906
rect 8092 5842 8148 5854
rect 8204 6018 8260 6076
rect 8204 5966 8206 6018
rect 8258 5966 8260 6018
rect 8204 5908 8260 5966
rect 8372 5962 8428 6412
rect 8372 5910 8374 5962
rect 8426 5910 8428 5962
rect 8372 5898 8428 5910
rect 8540 5906 8596 5918
rect 7980 5134 8036 5292
rect 7756 5070 7758 5122
rect 7810 5070 7812 5122
rect 7756 5012 7812 5070
rect 7924 5122 8036 5134
rect 7924 5070 7926 5122
rect 7978 5070 8036 5122
rect 7924 5068 8036 5070
rect 7924 5058 7980 5068
rect 7756 4946 7812 4956
rect 4788 4498 4844 4508
rect 7084 4498 7140 4508
rect 7756 4564 7812 4574
rect 7756 4470 7812 4508
rect 4172 4450 4432 4452
rect 4172 4398 4174 4450
rect 4226 4398 4432 4450
rect 4172 4396 4432 4398
rect 4172 4386 4228 4396
rect 3928 4330 3984 4342
rect 8092 4340 8148 4350
rect 8204 4340 8260 5852
rect 8540 5854 8542 5906
rect 8594 5854 8596 5906
rect 8316 5348 8372 5358
rect 8540 5348 8596 5854
rect 8316 5346 8596 5348
rect 8316 5294 8318 5346
rect 8370 5294 8596 5346
rect 8316 5292 8596 5294
rect 8316 5282 8372 5292
rect 8652 5236 8708 8204
rect 9100 8194 9156 8204
rect 9268 8202 9324 8214
rect 9268 8150 9270 8202
rect 9322 8150 9324 8202
rect 9436 8206 9438 8258
rect 9490 8206 9492 8258
rect 9436 8194 9492 8206
rect 9716 8484 9772 8934
rect 9828 8484 9884 8494
rect 9716 8482 9884 8484
rect 9716 8430 9830 8482
rect 9882 8430 9884 8482
rect 9716 8428 9884 8430
rect 9548 8258 9604 8428
rect 9828 8418 9884 8428
rect 9548 8206 9550 8258
rect 9602 8206 9604 8258
rect 9548 8194 9604 8206
rect 9268 7700 9324 8150
rect 9268 7634 9324 7644
rect 9192 7084 9456 7094
rect 9248 7028 9296 7084
rect 9352 7028 9400 7084
rect 9192 7018 9456 7028
rect 9996 6692 10052 9100
rect 10220 9044 10276 9054
rect 10220 8950 10276 8988
rect 10780 9042 10836 9100
rect 10780 8990 10782 9042
rect 10834 8990 10836 9042
rect 10780 8978 10836 8990
rect 10462 8818 10518 8830
rect 10462 8766 10464 8818
rect 10516 8766 10518 8818
rect 10462 8482 10518 8766
rect 10462 8430 10464 8482
rect 10516 8430 10518 8482
rect 10462 8418 10518 8430
rect 10892 8372 10948 13916
rect 11116 13906 11172 13916
rect 11788 13972 11844 13982
rect 11788 13914 11844 13916
rect 11788 13862 11790 13914
rect 11842 13862 11844 13914
rect 11788 13850 11844 13862
rect 12012 13972 12068 13982
rect 12236 13972 12292 15262
rect 12012 13802 12068 13916
rect 11676 13746 11732 13758
rect 11676 13694 11678 13746
rect 11730 13694 11732 13746
rect 12012 13750 12014 13802
rect 12066 13750 12068 13802
rect 12012 13738 12068 13750
rect 12124 13916 12292 13972
rect 12572 15301 12574 15353
rect 12626 15301 12628 15353
rect 12572 14532 12628 15301
rect 12572 13972 12628 14476
rect 11676 13076 11732 13694
rect 11564 12404 11620 12414
rect 11564 12310 11620 12348
rect 11676 12180 11732 13020
rect 12124 13188 12180 13916
rect 12572 13906 12628 13916
rect 12796 15314 12852 15326
rect 12796 15262 12798 15314
rect 12850 15262 12852 15314
rect 12236 13746 12292 13758
rect 12236 13694 12238 13746
rect 12290 13694 12292 13746
rect 12236 13300 12292 13694
rect 12236 13234 12292 13244
rect 12796 13300 12852 15262
rect 12796 13234 12852 13244
rect 12012 12964 12068 12974
rect 12124 12964 12180 13132
rect 12348 13076 12404 13086
rect 12012 12962 12180 12964
rect 12012 12910 12014 12962
rect 12066 12910 12180 12962
rect 12012 12908 12180 12910
rect 12236 12964 12292 12987
rect 12348 12982 12404 13020
rect 12012 12898 12068 12908
rect 12236 12895 12238 12908
rect 12290 12895 12292 12908
rect 12236 12883 12292 12895
rect 11852 12572 12116 12582
rect 11908 12516 11956 12572
rect 12012 12516 12060 12572
rect 11852 12506 12116 12516
rect 11900 12180 11956 12190
rect 12012 12180 12068 12190
rect 11676 12178 12068 12180
rect 11676 12126 11902 12178
rect 11954 12126 12014 12178
rect 12066 12126 12068 12178
rect 11676 12124 12068 12126
rect 11900 12114 11956 12124
rect 12012 12114 12068 12124
rect 12236 12180 12292 12190
rect 12236 12086 12292 12124
rect 12516 11956 12572 11966
rect 12516 11954 12740 11956
rect 12516 11902 12518 11954
rect 12570 11902 12740 11954
rect 12516 11900 12740 11902
rect 12516 11890 12572 11900
rect 11852 11004 12116 11014
rect 11908 10948 11956 11004
rect 12012 10948 12060 11004
rect 11852 10938 12116 10948
rect 11852 9436 12116 9446
rect 11908 9380 11956 9436
rect 12012 9380 12060 9436
rect 11852 9370 12116 9380
rect 12684 9156 12740 11900
rect 12684 9090 12740 9100
rect 11004 9044 11060 9054
rect 11004 9042 11172 9044
rect 11004 8990 11006 9042
rect 11058 8990 11172 9042
rect 11004 8988 11172 8990
rect 11004 8978 11060 8988
rect 10892 8306 10948 8316
rect 11004 8482 11060 8494
rect 11004 8430 11006 8482
rect 11058 8430 11060 8482
rect 9996 6626 10052 6636
rect 8876 5908 8932 5918
rect 8876 5346 8932 5852
rect 9192 5516 9456 5526
rect 9248 5460 9296 5516
rect 9352 5460 9400 5516
rect 9192 5450 9456 5460
rect 8876 5294 8878 5346
rect 8930 5294 8932 5346
rect 8876 5282 8932 5294
rect 9604 5348 9660 5358
rect 8652 5170 8708 5180
rect 9212 5236 9268 5246
rect 9212 5122 9268 5180
rect 9604 5234 9660 5292
rect 9604 5182 9606 5234
rect 9658 5182 9660 5234
rect 9604 5170 9660 5182
rect 9212 5070 9214 5122
rect 9266 5070 9268 5122
rect 9212 5058 9268 5070
rect 10668 5124 10724 5134
rect 10668 5030 10724 5068
rect 11004 5122 11060 8430
rect 11116 6692 11172 8988
rect 12348 9042 12404 9054
rect 12348 8990 12350 9042
rect 12402 8990 12404 9042
rect 11284 8932 11340 8942
rect 11284 8838 11340 8876
rect 12124 8932 12180 8942
rect 12124 8260 12180 8876
rect 12236 8874 12292 8886
rect 12236 8822 12238 8874
rect 12290 8822 12292 8874
rect 12236 8484 12292 8822
rect 12236 8418 12292 8428
rect 12124 8204 12292 8260
rect 11852 7868 12116 7878
rect 11908 7812 11956 7868
rect 12012 7812 12060 7868
rect 11852 7802 12116 7812
rect 11116 5908 11172 6636
rect 11852 6300 12116 6310
rect 11908 6244 11956 6300
rect 12012 6244 12060 6300
rect 11852 6234 12116 6244
rect 12236 6132 12292 8204
rect 11340 6074 11396 6086
rect 11340 6022 11342 6074
rect 11394 6022 11396 6074
rect 11228 5908 11284 5918
rect 11116 5906 11284 5908
rect 11116 5854 11230 5906
rect 11282 5854 11284 5906
rect 11116 5852 11284 5854
rect 11004 5070 11006 5122
rect 11058 5070 11060 5122
rect 11004 5058 11060 5070
rect 11228 5124 11284 5852
rect 11228 5058 11284 5068
rect 8708 5012 8764 5022
rect 8708 4562 8764 4956
rect 11340 4900 11396 6022
rect 11788 6076 12292 6132
rect 11564 5921 11620 5933
rect 11564 5869 11566 5921
rect 11618 5869 11620 5921
rect 11564 5348 11620 5869
rect 11564 5122 11620 5292
rect 11564 5070 11566 5122
rect 11618 5070 11620 5122
rect 11564 5058 11620 5070
rect 11676 5124 11732 5134
rect 11396 4844 11620 4900
rect 11340 4834 11396 4844
rect 8708 4510 8710 4562
rect 8762 4510 8764 4562
rect 8708 4498 8764 4510
rect 8092 4338 8260 4340
rect 3052 4274 3108 4286
rect 8092 4286 8094 4338
rect 8146 4286 8260 4338
rect 8092 4284 8260 4286
rect 11564 4350 11620 4844
rect 11676 4564 11732 5068
rect 11788 5122 11844 6076
rect 11900 5906 11956 5918
rect 11900 5854 11902 5906
rect 11954 5854 11956 5906
rect 11900 5348 11956 5854
rect 12068 5684 12124 5694
rect 12348 5684 12404 8990
rect 12908 8372 12964 16156
rect 13132 9716 13188 16268
rect 13356 14308 13412 17388
rect 14252 16324 14308 17614
rect 14364 17668 14420 17678
rect 14364 17574 14420 17612
rect 14924 17444 14980 18956
rect 15036 18674 15092 19180
rect 16044 19234 16100 19246
rect 18284 19236 18340 19246
rect 16044 19182 16046 19234
rect 16098 19182 16100 19234
rect 15764 19012 15820 19022
rect 15764 18918 15820 18956
rect 15036 18622 15038 18674
rect 15090 18622 15092 18674
rect 15036 18610 15092 18622
rect 16044 18452 16100 19182
rect 17724 19234 18340 19236
rect 17724 19182 18286 19234
rect 18338 19182 18340 19234
rect 17724 19180 18340 19182
rect 17172 18844 17436 18854
rect 17228 18788 17276 18844
rect 17332 18788 17380 18844
rect 17172 18778 17436 18788
rect 16044 18386 16100 18396
rect 14512 16492 14776 16502
rect 14568 16436 14616 16492
rect 14672 16436 14720 16492
rect 14512 16426 14776 16436
rect 14924 16324 14980 17388
rect 17172 17276 17436 17286
rect 17228 17220 17276 17276
rect 17332 17220 17380 17276
rect 17172 17210 17436 17220
rect 14252 16268 14420 16324
rect 14252 16100 14308 16110
rect 14252 16006 14308 16044
rect 13916 15092 13972 15102
rect 13804 14532 13860 14542
rect 13804 14438 13860 14476
rect 13524 14420 13580 14430
rect 13524 14418 13748 14420
rect 13524 14366 13526 14418
rect 13578 14366 13748 14418
rect 13524 14364 13748 14366
rect 13524 14354 13580 14364
rect 13356 14242 13412 14252
rect 13524 13524 13580 13534
rect 13524 13430 13580 13468
rect 13524 12852 13580 12862
rect 13524 12758 13580 12796
rect 13244 12404 13300 12414
rect 13244 12178 13300 12348
rect 13244 12126 13246 12178
rect 13298 12126 13300 12178
rect 13244 12114 13300 12126
rect 13580 12205 13636 12217
rect 13580 12153 13582 12205
rect 13634 12153 13636 12205
rect 13580 9828 13636 12153
rect 13692 12180 13748 14364
rect 13804 13748 13860 13758
rect 13916 13748 13972 15036
rect 13804 13746 13972 13748
rect 13804 13694 13806 13746
rect 13858 13694 13972 13746
rect 13804 13692 13972 13694
rect 13804 13682 13860 13692
rect 13804 13188 13860 13198
rect 13804 12962 13860 13132
rect 13804 12910 13806 12962
rect 13858 12910 13860 12962
rect 13804 12898 13860 12910
rect 13916 12962 13972 13692
rect 14028 14530 14084 14542
rect 14028 14478 14030 14530
rect 14082 14478 14084 14530
rect 14028 13746 14084 14478
rect 14028 13694 14030 13746
rect 14082 13694 14084 13746
rect 14028 13076 14084 13694
rect 14252 13748 14308 13758
rect 14028 13010 14084 13020
rect 14140 13524 14196 13534
rect 13916 12910 13918 12962
rect 13970 12910 13972 12962
rect 13916 12898 13972 12910
rect 14028 12740 14084 12750
rect 14028 12346 14084 12684
rect 14028 12294 14030 12346
rect 14082 12294 14084 12346
rect 14028 12282 14084 12294
rect 13692 12114 13748 12124
rect 13916 12180 13972 12190
rect 14140 12180 14196 13468
rect 14252 13074 14308 13692
rect 14364 13188 14420 16268
rect 14812 16268 14980 16324
rect 14700 16042 14756 16054
rect 14700 15990 14702 16042
rect 14754 15990 14756 16042
rect 14700 15204 14756 15990
rect 14812 15764 14868 16268
rect 14924 16100 14980 16110
rect 15372 16100 15428 16110
rect 14924 16006 14980 16044
rect 15036 16098 15428 16100
rect 15036 16046 15374 16098
rect 15426 16046 15428 16098
rect 15036 16044 15428 16046
rect 15036 15930 15092 16044
rect 15372 16034 15428 16044
rect 15036 15878 15038 15930
rect 15090 15878 15092 15930
rect 15036 15866 15092 15878
rect 15708 15876 15764 15886
rect 15260 15874 15764 15876
rect 15260 15822 15710 15874
rect 15762 15822 15764 15874
rect 15260 15820 15764 15822
rect 14812 15708 15092 15764
rect 14924 15329 14980 15341
rect 14924 15316 14926 15329
rect 14978 15316 14980 15329
rect 14924 15237 14980 15260
rect 14812 15204 14868 15214
rect 14700 15202 14868 15204
rect 14700 15150 14814 15202
rect 14866 15150 14868 15202
rect 14700 15148 14868 15150
rect 15036 15148 15092 15708
rect 14812 15092 14868 15148
rect 14812 15026 14868 15036
rect 14924 15092 15092 15148
rect 15260 15314 15316 15820
rect 15708 15810 15764 15820
rect 17172 15708 17436 15718
rect 17228 15652 17276 15708
rect 17332 15652 17380 15708
rect 17172 15642 17436 15652
rect 15260 15262 15262 15314
rect 15314 15262 15316 15314
rect 14512 14924 14776 14934
rect 14568 14868 14616 14924
rect 14672 14868 14720 14924
rect 14512 14858 14776 14868
rect 14512 13356 14776 13366
rect 14568 13300 14616 13356
rect 14672 13300 14720 13356
rect 14512 13290 14776 13300
rect 14588 13188 14644 13198
rect 14364 13132 14532 13188
rect 14252 13022 14254 13074
rect 14306 13022 14308 13074
rect 14252 13010 14308 13022
rect 14364 12964 14420 12974
rect 14364 12895 14366 12908
rect 14418 12895 14420 12908
rect 14364 12870 14420 12895
rect 13916 12178 14196 12180
rect 13916 12126 13918 12178
rect 13970 12126 14196 12178
rect 13916 12124 14196 12126
rect 14476 12628 14532 13132
rect 14588 12964 14644 13132
rect 14588 12898 14644 12908
rect 14700 12962 14756 12974
rect 14700 12910 14702 12962
rect 14754 12910 14756 12962
rect 13916 12114 13972 12124
rect 14476 11956 14532 12572
rect 14140 11900 14532 11956
rect 14700 11956 14756 12910
rect 14028 9938 14084 9950
rect 14028 9886 14030 9938
rect 14082 9886 14084 9938
rect 13580 9826 13748 9828
rect 13580 9774 13582 9826
rect 13634 9774 13748 9826
rect 13580 9772 13748 9774
rect 13580 9762 13636 9772
rect 13132 9660 13524 9716
rect 13468 9166 13524 9660
rect 13024 9156 13080 9166
rect 13468 9154 13580 9166
rect 13468 9102 13526 9154
rect 13578 9102 13580 9154
rect 13468 9100 13580 9102
rect 13024 9080 13080 9100
rect 13524 9090 13580 9100
rect 13024 9028 13026 9080
rect 13078 9028 13080 9080
rect 13024 9016 13080 9028
rect 12908 8316 13412 8372
rect 13356 8258 13412 8316
rect 13356 8206 13358 8258
rect 13410 8206 13412 8258
rect 13356 6916 13412 8206
rect 13356 6850 13412 6860
rect 13580 8258 13636 8270
rect 13580 8206 13582 8258
rect 13634 8206 13636 8258
rect 13580 6692 13636 8206
rect 13580 6626 13636 6636
rect 12068 5682 12180 5684
rect 12068 5630 12070 5682
rect 12122 5630 12180 5682
rect 12068 5618 12180 5630
rect 11900 5282 11956 5292
rect 11788 5070 11790 5122
rect 11842 5070 11844 5122
rect 11788 5058 11844 5070
rect 12012 5234 12068 5246
rect 12012 5182 12014 5234
rect 12066 5182 12068 5234
rect 12012 5124 12068 5182
rect 12012 5058 12068 5068
rect 12124 4900 12180 5618
rect 12348 5236 12404 5628
rect 13524 5796 13580 5806
rect 12684 5348 12740 5358
rect 12348 5170 12404 5180
rect 12572 5236 12628 5246
rect 12236 5124 12292 5134
rect 12236 5030 12292 5068
rect 12572 5107 12628 5180
rect 12684 5234 12740 5292
rect 13524 5346 13580 5740
rect 13524 5294 13526 5346
rect 13578 5294 13580 5346
rect 13524 5282 13580 5294
rect 12684 5182 12686 5234
rect 12738 5182 12740 5234
rect 12684 5170 12740 5182
rect 12572 5055 12574 5107
rect 12626 5055 12628 5107
rect 12572 5043 12628 5055
rect 13692 5122 13748 9772
rect 13916 9811 13972 9823
rect 13916 9759 13918 9811
rect 13970 9759 13972 9811
rect 13916 9156 13972 9759
rect 14028 9268 14084 9886
rect 14028 9202 14084 9212
rect 13916 9090 13972 9100
rect 13804 9070 13860 9082
rect 13804 9044 13806 9070
rect 13858 9044 13860 9070
rect 14028 9070 14084 9082
rect 14028 9018 14030 9070
rect 14082 9044 14084 9070
rect 14140 9044 14196 11900
rect 14700 11890 14756 11900
rect 14512 11788 14776 11798
rect 14568 11732 14616 11788
rect 14672 11732 14720 11788
rect 14512 11722 14776 11732
rect 14512 10220 14776 10230
rect 14568 10164 14616 10220
rect 14672 10164 14720 10220
rect 14512 10154 14776 10164
rect 14364 10052 14420 10062
rect 14364 9098 14420 9996
rect 14924 9492 14980 15092
rect 15260 14532 15316 15262
rect 15260 14466 15316 14476
rect 17172 14140 17436 14150
rect 17228 14084 17276 14140
rect 17332 14084 17380 14140
rect 17172 14074 17436 14084
rect 17276 13748 17332 13758
rect 17164 13746 17332 13748
rect 17164 13694 17278 13746
rect 17330 13694 17332 13746
rect 17164 13692 17332 13694
rect 16828 13076 16884 13086
rect 16380 12962 16436 12974
rect 16380 12910 16382 12962
rect 16434 12910 16436 12962
rect 15316 12628 15372 12638
rect 15316 12402 15372 12572
rect 16380 12628 16436 12910
rect 16828 12923 16884 13020
rect 16828 12871 16830 12923
rect 16882 12871 16884 12923
rect 16828 12859 16884 12871
rect 17052 12962 17108 12974
rect 17052 12910 17054 12962
rect 17106 12910 17108 12962
rect 16380 12562 16436 12572
rect 15316 12350 15318 12402
rect 15370 12350 15372 12402
rect 15316 12338 15372 12350
rect 15148 12178 15204 12190
rect 15148 12126 15150 12178
rect 15202 12126 15204 12178
rect 15148 10052 15204 12126
rect 17052 11396 17108 12910
rect 17164 12794 17220 13692
rect 17276 13682 17332 13692
rect 17612 13522 17668 13534
rect 17612 13470 17614 13522
rect 17666 13470 17668 13522
rect 17612 12964 17668 13470
rect 17612 12870 17668 12908
rect 17164 12742 17166 12794
rect 17218 12742 17220 12794
rect 17164 12730 17220 12742
rect 17172 12572 17436 12582
rect 17228 12516 17276 12572
rect 17332 12516 17380 12572
rect 17172 12506 17436 12516
rect 17724 12180 17780 19180
rect 18284 19170 18340 19180
rect 19068 19234 19124 19246
rect 19068 19182 19070 19234
rect 19122 19182 19124 19234
rect 17836 18450 17892 18462
rect 17836 18398 17838 18450
rect 17890 18398 17892 18450
rect 17836 12740 17892 18398
rect 18172 18452 18228 18462
rect 18172 18358 18228 18396
rect 19068 18452 19124 19182
rect 19628 19236 19684 19964
rect 19740 19954 19796 19964
rect 20636 20018 20692 20030
rect 20636 19966 20638 20018
rect 20690 19966 20692 20018
rect 19832 19628 20096 19638
rect 19888 19572 19936 19628
rect 19992 19572 20040 19628
rect 19832 19562 20096 19572
rect 20636 19460 20692 19966
rect 21756 20018 21812 20030
rect 21756 19966 21758 20018
rect 21810 19966 21812 20018
rect 20636 19394 20692 19404
rect 21532 19460 21588 19470
rect 21756 19460 21812 19966
rect 21532 19458 21812 19460
rect 21532 19406 21534 19458
rect 21586 19406 21812 19458
rect 21532 19404 21812 19406
rect 21532 19394 21588 19404
rect 19628 19170 19684 19180
rect 19740 19234 19796 19246
rect 19740 19182 19742 19234
rect 19794 19182 19796 19234
rect 19516 19066 19572 19078
rect 19516 19014 19518 19066
rect 19570 19014 19572 19066
rect 19516 18788 19572 19014
rect 19740 19012 19796 19182
rect 19740 18946 19796 18956
rect 20076 19234 20132 19246
rect 20076 19182 20078 19234
rect 20130 19182 20132 19234
rect 19068 18386 19124 18396
rect 19292 18732 19572 18788
rect 19292 18450 19348 18732
rect 20076 18574 20132 19182
rect 21196 19234 21252 19246
rect 21196 19182 21198 19234
rect 21250 19182 21252 19234
rect 20412 19012 20468 19022
rect 20412 18918 20468 18956
rect 20860 19012 20916 19022
rect 20076 18562 20188 18574
rect 20076 18510 20134 18562
rect 20186 18510 20188 18562
rect 20076 18508 20188 18510
rect 20132 18498 20188 18508
rect 19292 18398 19294 18450
rect 19346 18398 19348 18450
rect 19292 18386 19348 18398
rect 19628 18452 19684 18462
rect 19628 18358 19684 18396
rect 19852 18452 19908 18462
rect 19852 18358 19908 18396
rect 20580 18452 20636 18462
rect 20580 18358 20636 18396
rect 20860 18450 20916 18956
rect 20860 18398 20862 18450
rect 20914 18398 20916 18450
rect 20860 18386 20916 18398
rect 20972 18452 21028 18462
rect 21196 18452 21252 19182
rect 22316 19124 22372 19134
rect 20972 18450 21252 18452
rect 20972 18398 20974 18450
rect 21026 18398 21252 18450
rect 20972 18396 21252 18398
rect 21588 18452 21644 18462
rect 18956 18340 19012 18350
rect 18956 18246 19012 18284
rect 19832 18060 20096 18070
rect 19888 18004 19936 18060
rect 19992 18004 20040 18060
rect 19832 17994 20096 18004
rect 18284 16884 18340 16894
rect 18228 16882 18340 16884
rect 18228 16830 18286 16882
rect 18338 16830 18340 16882
rect 18228 16818 18340 16830
rect 18228 16322 18284 16818
rect 18620 16658 18676 16670
rect 18620 16606 18622 16658
rect 18674 16606 18676 16658
rect 18620 16548 18676 16606
rect 18620 16482 18676 16492
rect 19832 16492 20096 16502
rect 19888 16436 19936 16492
rect 19992 16436 20040 16492
rect 19832 16426 20096 16436
rect 19348 16324 19404 16334
rect 18228 16270 18230 16322
rect 18282 16270 18284 16322
rect 18228 16258 18284 16270
rect 18508 16322 19404 16324
rect 18508 16270 19350 16322
rect 19402 16270 19404 16322
rect 18508 16268 19404 16270
rect 18508 16098 18564 16268
rect 19348 16258 19404 16268
rect 18508 16046 18510 16098
rect 18562 16046 18564 16098
rect 18508 15358 18564 16046
rect 18284 15314 18340 15326
rect 18284 15262 18286 15314
rect 18338 15262 18340 15314
rect 18508 15306 18510 15358
rect 18562 15306 18564 15358
rect 18732 16098 18788 16110
rect 18732 16046 18734 16098
rect 18786 16046 18788 16098
rect 18508 15294 18564 15306
rect 18620 15316 18676 15326
rect 18060 13076 18116 13086
rect 18060 12982 18116 13020
rect 17836 12674 17892 12684
rect 17948 12918 18004 12930
rect 17948 12866 17950 12918
rect 18002 12866 18004 12918
rect 17948 12404 18004 12866
rect 18284 12516 18340 15262
rect 18620 15202 18676 15260
rect 18620 15150 18622 15202
rect 18674 15150 18676 15202
rect 18620 15138 18676 15150
rect 18284 12450 18340 12460
rect 18508 12516 18564 12526
rect 17948 12338 18004 12348
rect 17052 11330 17108 11340
rect 17612 12124 17780 12180
rect 18060 12180 18116 12190
rect 18340 12180 18396 12190
rect 18060 12178 18396 12180
rect 18060 12126 18062 12178
rect 18114 12126 18342 12178
rect 18394 12126 18396 12178
rect 18060 12124 18396 12126
rect 17172 11004 17436 11014
rect 17228 10948 17276 11004
rect 17332 10948 17380 11004
rect 17172 10938 17436 10948
rect 15148 9986 15204 9996
rect 14082 9018 14196 9044
rect 14028 8988 14196 9018
rect 14252 9070 14308 9082
rect 14252 9018 14254 9070
rect 14306 9018 14308 9070
rect 14364 9046 14366 9098
rect 14418 9046 14420 9098
rect 14364 9034 14420 9046
rect 14588 9436 14980 9492
rect 17172 9436 17436 9446
rect 13804 8494 13860 8988
rect 13804 8482 13916 8494
rect 13804 8430 13862 8482
rect 13914 8430 13916 8482
rect 13804 8428 13916 8430
rect 13860 8418 13916 8428
rect 14252 8036 14308 9018
rect 14588 8932 14644 9436
rect 17228 9380 17276 9436
rect 17332 9380 17380 9436
rect 17172 9370 17436 9380
rect 14958 9268 15014 9278
rect 14958 9080 15014 9212
rect 17612 9156 17668 12124
rect 18060 12114 18116 12124
rect 18340 12114 18396 12124
rect 17724 11954 17780 11966
rect 17724 11902 17726 11954
rect 17778 11902 17780 11954
rect 17724 11396 17780 11902
rect 17724 11330 17780 11340
rect 17948 11956 18004 11966
rect 17948 10836 18004 11900
rect 18508 11844 18564 12460
rect 17612 9090 17668 9100
rect 17724 10834 18004 10836
rect 17724 10782 17950 10834
rect 18002 10782 18004 10834
rect 17724 10780 18004 10782
rect 14700 9044 14756 9054
rect 14700 8950 14756 8988
rect 14812 9042 14868 9054
rect 14812 8990 14814 9042
rect 14866 8990 14868 9042
rect 14958 9028 14960 9080
rect 15012 9028 15014 9080
rect 14958 9016 15014 9028
rect 14252 7970 14308 7980
rect 14364 8876 14644 8932
rect 14196 6020 14252 6030
rect 14364 6020 14420 8876
rect 14812 8820 14868 8990
rect 14812 8754 14868 8764
rect 15372 8818 15428 8830
rect 15372 8766 15374 8818
rect 15426 8766 15428 8818
rect 14512 8652 14776 8662
rect 14568 8596 14616 8652
rect 14672 8596 14720 8652
rect 14512 8586 14776 8596
rect 15372 8372 15428 8766
rect 15372 8306 15428 8316
rect 17500 8372 17556 8382
rect 17500 8220 17556 8316
rect 17500 8168 17502 8220
rect 17554 8168 17556 8220
rect 17500 8156 17556 8168
rect 17724 8260 17780 10780
rect 17948 10770 18004 10780
rect 18284 11788 18564 11844
rect 18620 12178 18676 12190
rect 18620 12126 18622 12178
rect 18674 12126 18676 12178
rect 18284 10610 18340 11788
rect 18620 11620 18676 12126
rect 18620 11554 18676 11564
rect 18732 12178 18788 16046
rect 18844 16100 18900 16110
rect 18844 16006 18900 16044
rect 19068 16100 19124 16110
rect 19068 16098 19236 16100
rect 19068 16046 19070 16098
rect 19122 16046 19236 16098
rect 19068 16044 19236 16046
rect 19068 16034 19124 16044
rect 19180 15482 19236 16044
rect 19180 15430 19182 15482
rect 19234 15430 19236 15482
rect 19180 15418 19236 15430
rect 20300 15596 20580 15652
rect 19404 15329 19460 15341
rect 19068 15316 19124 15326
rect 19068 15222 19124 15260
rect 19404 15277 19406 15329
rect 19458 15277 19460 15329
rect 19404 13636 19460 15277
rect 19832 14924 20096 14934
rect 19888 14868 19936 14924
rect 19992 14868 20040 14924
rect 19832 14858 20096 14868
rect 20300 14308 20356 15596
rect 20076 13773 20132 13785
rect 19740 13748 19796 13758
rect 19740 13654 19796 13692
rect 20076 13721 20078 13773
rect 20130 13721 20132 13773
rect 19404 13570 19460 13580
rect 20076 13524 20132 13721
rect 20076 13468 20244 13524
rect 19832 13356 20096 13366
rect 19888 13300 19936 13356
rect 19992 13300 20040 13356
rect 19832 13290 20096 13300
rect 20188 13076 20244 13468
rect 20188 13010 20244 13020
rect 20300 12852 20356 14252
rect 20412 15482 20468 15494
rect 20412 15430 20414 15482
rect 20466 15430 20468 15482
rect 20412 13746 20468 15430
rect 20524 15314 20580 15596
rect 20972 15382 21028 18396
rect 21588 18358 21644 18396
rect 22316 18452 22372 19068
rect 22492 18844 22756 18854
rect 22548 18788 22596 18844
rect 22652 18788 22700 18844
rect 22492 18778 22756 18788
rect 22316 18358 22372 18396
rect 21980 18228 22036 18238
rect 21980 18226 22260 18228
rect 21980 18174 21982 18226
rect 22034 18174 22260 18226
rect 21980 18172 22260 18174
rect 21980 18162 22036 18172
rect 21588 16996 21644 17006
rect 21588 16902 21644 16940
rect 20524 15262 20526 15314
rect 20578 15262 20580 15314
rect 20524 15250 20580 15262
rect 20916 15370 21028 15382
rect 20916 15318 20918 15370
rect 20970 15318 21028 15370
rect 20916 15260 21028 15318
rect 20972 15092 21028 15260
rect 21196 16884 21252 16894
rect 21196 15314 21252 16828
rect 21980 16884 22036 16894
rect 21980 16790 22036 16828
rect 21196 15262 21198 15314
rect 21250 15262 21252 15314
rect 21196 15250 21252 15262
rect 20972 15036 21364 15092
rect 21196 14532 21252 14542
rect 20524 14530 21252 14532
rect 20524 14478 21198 14530
rect 21250 14478 21252 14530
rect 20524 14476 21252 14478
rect 20524 13914 20580 14476
rect 21196 14466 21252 14476
rect 20524 13862 20526 13914
rect 20578 13862 20580 13914
rect 20524 13850 20580 13862
rect 20412 13694 20414 13746
rect 20466 13694 20468 13746
rect 20412 13682 20468 13694
rect 21308 13748 21364 15036
rect 21532 14308 21588 14318
rect 21532 14214 21588 14252
rect 21458 13783 21514 13795
rect 21458 13748 21460 13783
rect 21308 13731 21460 13748
rect 21512 13731 21514 13783
rect 21308 13692 21514 13731
rect 21644 13746 21700 13758
rect 21644 13694 21646 13746
rect 21698 13694 21700 13746
rect 21084 13636 21140 13646
rect 21084 13542 21140 13580
rect 20804 13300 20860 13310
rect 20804 13074 20860 13244
rect 20804 13022 20806 13074
rect 20858 13022 20860 13074
rect 20804 13010 20860 13022
rect 20972 13076 21028 13086
rect 20300 12786 20356 12796
rect 18732 12126 18734 12178
rect 18786 12126 18788 12178
rect 18620 11396 18676 11406
rect 18620 11302 18676 11340
rect 18284 10558 18286 10610
rect 18338 10558 18340 10610
rect 18172 10052 18228 10062
rect 18284 10052 18340 10558
rect 17948 10050 18340 10052
rect 17948 9998 18174 10050
rect 18226 9998 18340 10050
rect 17948 9996 18340 9998
rect 17836 9828 17892 9866
rect 17836 9762 17892 9772
rect 17172 7868 17436 7878
rect 17228 7812 17276 7868
rect 17332 7812 17380 7868
rect 17172 7802 17436 7812
rect 14512 7084 14776 7094
rect 14568 7028 14616 7084
rect 14672 7028 14720 7084
rect 14512 7018 14776 7028
rect 14196 6018 14420 6020
rect 14196 5966 14198 6018
rect 14250 5966 14420 6018
rect 14196 5964 14420 5966
rect 14588 6916 14644 6926
rect 14588 6132 14644 6860
rect 17172 6300 17436 6310
rect 17228 6244 17276 6300
rect 17332 6244 17380 6300
rect 17172 6234 17436 6244
rect 15036 6132 15092 6142
rect 14588 6130 15092 6132
rect 14588 6078 15038 6130
rect 15090 6078 15092 6130
rect 14588 6076 15092 6078
rect 14196 5954 14252 5964
rect 14476 5908 14532 5918
rect 14476 5814 14532 5852
rect 14588 5906 14644 6076
rect 15036 6066 15092 6076
rect 14588 5854 14590 5906
rect 14642 5854 14644 5906
rect 14588 5842 14644 5854
rect 15372 5906 15428 5918
rect 15372 5854 15374 5906
rect 15426 5854 15428 5906
rect 15372 5796 15428 5854
rect 16828 5908 16884 5918
rect 15932 5796 15988 5806
rect 15428 5740 15540 5796
rect 15372 5730 15428 5740
rect 14512 5516 14776 5526
rect 14568 5460 14616 5516
rect 14672 5460 14720 5516
rect 14512 5450 14776 5460
rect 14028 5348 14084 5358
rect 13692 5070 13694 5122
rect 13746 5070 13748 5122
rect 13580 5012 13636 5022
rect 12572 4900 12628 4910
rect 12124 4844 12292 4900
rect 11852 4732 12116 4742
rect 11908 4676 11956 4732
rect 12012 4676 12060 4732
rect 11852 4666 12116 4676
rect 11676 4508 12068 4564
rect 12012 4450 12068 4508
rect 12012 4398 12014 4450
rect 12066 4398 12068 4450
rect 12012 4386 12068 4398
rect 11564 4340 11676 4350
rect 11844 4340 11900 4350
rect 11564 4338 11900 4340
rect 11564 4286 11622 4338
rect 11674 4286 11846 4338
rect 11898 4286 11900 4338
rect 11564 4284 11900 4286
rect 8092 4274 8148 4284
rect 11620 4274 11676 4284
rect 11844 4274 11900 4284
rect 12236 4338 12292 4844
rect 12236 4286 12238 4338
rect 12290 4286 12292 4338
rect 12572 4394 12628 4844
rect 13580 4574 13636 4956
rect 13692 4900 13748 5070
rect 13804 5124 13860 5134
rect 13804 5030 13860 5068
rect 14028 5122 14084 5292
rect 14028 5070 14030 5122
rect 14082 5070 14084 5122
rect 14028 5058 14084 5070
rect 15260 5122 15316 5134
rect 15260 5070 15262 5122
rect 15314 5070 15316 5122
rect 14308 5012 14364 5022
rect 14308 5010 14532 5012
rect 14308 4958 14310 5010
rect 14362 4958 14532 5010
rect 14308 4956 14532 4958
rect 14308 4946 14364 4956
rect 13692 4844 14196 4900
rect 13580 4564 13692 4574
rect 13580 4508 13636 4564
rect 13636 4470 13692 4508
rect 14140 4562 14196 4844
rect 14140 4510 14142 4562
rect 14194 4510 14196 4562
rect 14140 4498 14196 4510
rect 12572 4342 12574 4394
rect 12626 4342 12628 4394
rect 12572 4330 12628 4342
rect 14476 4338 14532 4956
rect 15260 4564 15316 5070
rect 15484 5083 15540 5740
rect 15596 5684 15652 5694
rect 15596 5234 15652 5628
rect 15596 5182 15598 5234
rect 15650 5182 15652 5234
rect 15596 5170 15652 5182
rect 15484 5031 15486 5083
rect 15538 5031 15540 5083
rect 15932 5122 15988 5740
rect 15932 5070 15934 5122
rect 15986 5070 15988 5122
rect 15932 5058 15988 5070
rect 16828 5460 16884 5852
rect 16828 5122 16884 5404
rect 17164 5572 17220 5582
rect 17164 5236 17220 5516
rect 17164 5142 17220 5180
rect 16828 5070 16830 5122
rect 16882 5070 16884 5122
rect 16828 5058 16884 5070
rect 17724 5122 17780 8204
rect 17836 9604 17892 9614
rect 17836 8258 17892 9548
rect 17948 9042 18004 9996
rect 18172 9986 18228 9996
rect 18508 9210 18564 9222
rect 18508 9158 18510 9210
rect 18562 9158 18564 9210
rect 17948 8990 17950 9042
rect 18002 8990 18004 9042
rect 17948 8978 18004 8990
rect 18172 9081 18228 9093
rect 18172 9029 18174 9081
rect 18226 9029 18228 9081
rect 18508 9044 18564 9158
rect 18172 8820 18228 9029
rect 17836 8206 17838 8258
rect 17890 8206 17892 8258
rect 17836 8194 17892 8206
rect 18060 8764 18228 8820
rect 18284 8988 18508 9044
rect 18060 8146 18116 8764
rect 18284 8372 18340 8988
rect 18508 8978 18564 8988
rect 18620 9042 18676 9054
rect 18620 8990 18622 9042
rect 18674 8990 18676 9042
rect 18228 8316 18340 8372
rect 18228 8314 18284 8316
rect 18228 8262 18230 8314
rect 18282 8262 18284 8314
rect 18228 8250 18284 8262
rect 18452 8260 18508 8270
rect 18452 8166 18508 8204
rect 18060 8094 18062 8146
rect 18114 8094 18116 8146
rect 17892 7700 17948 7710
rect 17892 7606 17948 7644
rect 18060 7474 18116 8094
rect 18340 8148 18396 8158
rect 18340 7698 18396 8092
rect 18340 7646 18342 7698
rect 18394 7646 18396 7698
rect 18340 7634 18396 7646
rect 18620 8146 18676 8990
rect 18620 8094 18622 8146
rect 18674 8094 18676 8146
rect 18060 7422 18062 7474
rect 18114 7422 18116 7474
rect 18060 7410 18116 7422
rect 18508 7476 18564 7486
rect 18620 7476 18676 8094
rect 18508 7474 18676 7476
rect 18508 7422 18510 7474
rect 18562 7422 18676 7474
rect 18508 7420 18676 7422
rect 18508 7410 18564 7420
rect 18508 5572 18564 5582
rect 18732 5572 18788 12126
rect 19068 12516 19124 12526
rect 19068 12178 19124 12460
rect 19516 12404 19572 12414
rect 19348 12234 19404 12246
rect 19348 12224 19350 12234
rect 19068 12126 19070 12178
rect 19122 12126 19124 12178
rect 19068 12114 19124 12126
rect 19292 12182 19350 12224
rect 19402 12182 19404 12234
rect 19292 12168 19404 12182
rect 19516 12180 19572 12348
rect 20188 12236 20468 12292
rect 20188 12222 20244 12236
rect 19852 12180 19908 12190
rect 19516 12178 19908 12180
rect 18844 12068 18900 12078
rect 18844 11394 18900 12012
rect 19124 11620 19180 11630
rect 19292 11620 19348 12168
rect 19516 12126 19854 12178
rect 19906 12126 19908 12178
rect 20188 12170 20190 12222
rect 20242 12170 20244 12222
rect 20188 12158 20244 12170
rect 19516 12124 19908 12126
rect 19516 12066 19572 12124
rect 19852 12114 19908 12124
rect 19516 12014 19518 12066
rect 19570 12014 19572 12066
rect 19516 12002 19572 12014
rect 20300 12068 20356 12078
rect 20412 12068 20468 12236
rect 20748 12068 20804 12078
rect 20412 12066 20804 12068
rect 20412 12014 20750 12066
rect 20802 12014 20804 12066
rect 20412 12012 20804 12014
rect 20300 11974 20356 12012
rect 20748 12002 20804 12012
rect 19832 11788 20096 11798
rect 19888 11732 19936 11788
rect 19992 11732 20040 11788
rect 19832 11722 20096 11732
rect 19180 11564 19348 11620
rect 19124 11526 19180 11564
rect 18844 11342 18846 11394
rect 18898 11342 18900 11394
rect 18844 11330 18900 11342
rect 19832 10220 20096 10230
rect 19888 10164 19936 10220
rect 19992 10164 20040 10220
rect 19832 10154 20096 10164
rect 20412 10052 20468 10062
rect 20972 10052 21028 13020
rect 19068 9828 19124 9838
rect 19068 9734 19124 9772
rect 19292 9828 19348 9838
rect 18900 9604 18956 9614
rect 18900 9510 18956 9548
rect 19292 9380 19348 9772
rect 20188 9828 20244 9838
rect 19460 9716 19516 9726
rect 19460 9622 19516 9660
rect 19292 9324 19460 9380
rect 18956 9044 19012 9054
rect 19292 9042 19348 9054
rect 18956 8950 19012 8988
rect 19124 8986 19180 8998
rect 19124 8934 19126 8986
rect 19178 8934 19180 8986
rect 19124 8932 19180 8934
rect 19124 8484 19180 8876
rect 19124 8418 19180 8428
rect 19292 8990 19294 9042
rect 19346 8990 19348 9042
rect 18844 8258 18900 8270
rect 18844 8206 18846 8258
rect 18898 8206 18900 8258
rect 18844 8148 18900 8206
rect 18844 8082 18900 8092
rect 19068 8202 19124 8214
rect 19068 8150 19070 8202
rect 19122 8150 19124 8202
rect 19068 7700 19124 8150
rect 19292 8148 19348 8990
rect 19404 9042 19460 9324
rect 19404 8990 19406 9042
rect 19458 8990 19460 9042
rect 19404 8978 19460 8990
rect 19684 9044 19740 9054
rect 19684 8950 19740 8988
rect 19832 8652 20096 8662
rect 19888 8596 19936 8652
rect 19992 8596 20040 8652
rect 19832 8586 20096 8596
rect 19292 8082 19348 8092
rect 20188 7924 20244 9772
rect 20300 9044 20356 9054
rect 20300 8950 20356 8988
rect 20412 8428 20468 9996
rect 20748 9996 21028 10052
rect 20524 9828 20580 9838
rect 20524 9734 20580 9772
rect 20748 9604 20804 9996
rect 20636 9268 20692 9278
rect 20636 9174 20692 9212
rect 20636 8932 20692 8942
rect 20636 8484 20692 8876
rect 20412 8372 20580 8428
rect 20188 7868 20300 7924
rect 19068 7634 19124 7644
rect 20244 7530 20300 7868
rect 20244 7478 20246 7530
rect 20298 7478 20300 7530
rect 20244 7466 20300 7478
rect 19516 7364 19572 7374
rect 18564 5516 18788 5572
rect 19404 5906 19460 5918
rect 19404 5854 19406 5906
rect 19458 5854 19460 5906
rect 17724 5070 17726 5122
rect 17778 5070 17780 5122
rect 15484 5019 15540 5031
rect 17724 4900 17780 5070
rect 17724 4834 17780 4844
rect 17836 5236 17892 5246
rect 17836 4954 17892 5180
rect 18060 5124 18116 5147
rect 18060 5055 18062 5068
rect 18114 5055 18116 5068
rect 18508 5122 18564 5516
rect 18620 5348 18676 5358
rect 18620 5290 18676 5292
rect 18620 5238 18622 5290
rect 18674 5238 18676 5290
rect 19404 5348 19460 5854
rect 19516 5906 19572 7308
rect 20412 7364 20468 7374
rect 20412 7270 20468 7308
rect 19832 7084 20096 7094
rect 19888 7028 19936 7084
rect 19992 7028 20040 7084
rect 19832 7018 20096 7028
rect 20524 6468 20580 8372
rect 20300 6412 20580 6468
rect 20636 7474 20692 8428
rect 20636 7422 20638 7474
rect 20690 7422 20692 7474
rect 19516 5854 19518 5906
rect 19570 5854 19572 5906
rect 19516 5842 19572 5854
rect 20076 5908 20132 5918
rect 20076 5814 20132 5852
rect 20300 5908 20356 6412
rect 20412 6132 20468 6142
rect 20636 6132 20692 7422
rect 20412 6130 20692 6132
rect 20412 6078 20414 6130
rect 20466 6078 20692 6130
rect 20412 6076 20692 6078
rect 20412 6066 20468 6076
rect 20356 5852 20580 5908
rect 20300 5842 20356 5852
rect 19796 5684 19852 5694
rect 19404 5282 19460 5292
rect 19628 5682 19852 5684
rect 19628 5630 19798 5682
rect 19850 5630 19852 5682
rect 19628 5628 19852 5630
rect 18620 5226 18676 5238
rect 19292 5236 19348 5246
rect 19628 5236 19684 5628
rect 19796 5618 19852 5628
rect 20300 5684 20356 5694
rect 19832 5516 20096 5526
rect 19888 5460 19936 5516
rect 19992 5460 20040 5516
rect 19832 5450 20096 5460
rect 19628 5180 19908 5236
rect 18508 5070 18510 5122
rect 18562 5070 18564 5122
rect 18508 5058 18564 5070
rect 18844 5124 18900 5134
rect 18060 5043 18116 5055
rect 18844 5030 18900 5068
rect 19292 5122 19348 5180
rect 19292 5070 19294 5122
rect 19346 5070 19348 5122
rect 19292 5058 19348 5070
rect 19404 5092 19628 5124
rect 19404 5068 19574 5092
rect 17836 4902 17838 4954
rect 17890 4902 17892 4954
rect 17172 4732 17436 4742
rect 17228 4676 17276 4732
rect 17332 4676 17380 4732
rect 17172 4666 17436 4676
rect 15260 4498 15316 4508
rect 17444 4564 17500 4574
rect 17444 4470 17500 4508
rect 12236 4274 12292 4286
rect 14476 4286 14478 4338
rect 14530 4286 14532 4338
rect 14476 4274 14532 4286
rect 17612 4340 17668 4350
rect 17836 4340 17892 4902
rect 19404 4562 19460 5068
rect 19572 5040 19574 5068
rect 19626 5040 19628 5092
rect 19572 5028 19628 5040
rect 19740 5012 19796 5022
rect 19628 4954 19684 4966
rect 19628 4902 19630 4954
rect 19682 4902 19684 4954
rect 19628 4900 19684 4902
rect 19740 4900 19796 4956
rect 19628 4844 19796 4900
rect 19404 4510 19406 4562
rect 19458 4510 19460 4562
rect 19404 4498 19460 4510
rect 17612 4338 17892 4340
rect 17612 4286 17614 4338
rect 17666 4286 17892 4338
rect 17612 4284 17892 4286
rect 19740 4340 19796 4350
rect 19852 4340 19908 5180
rect 20020 5012 20076 5022
rect 20020 4450 20076 4956
rect 20020 4398 20022 4450
rect 20074 4398 20076 4450
rect 20020 4386 20076 4398
rect 19740 4338 19908 4340
rect 19740 4286 19742 4338
rect 19794 4286 19908 4338
rect 19740 4284 19908 4286
rect 20300 4338 20356 5628
rect 20524 5346 20580 5852
rect 20524 5294 20526 5346
rect 20578 5294 20580 5346
rect 20524 5282 20580 5294
rect 20300 4286 20302 4338
rect 20354 4286 20356 4338
rect 17612 4274 17668 4284
rect 19740 4274 19796 4284
rect 20300 4274 20356 4286
rect 20524 4340 20580 4350
rect 20524 4246 20580 4284
rect 20748 4170 20804 9548
rect 20860 9828 20916 9838
rect 21308 9828 21364 13692
rect 21644 13188 21700 13694
rect 21644 13122 21700 13132
rect 21756 13746 21812 13758
rect 21756 13694 21758 13746
rect 21810 13694 21812 13746
rect 21476 13076 21532 13086
rect 21476 12982 21532 13020
rect 21420 12066 21476 12078
rect 21420 12014 21422 12066
rect 21474 12014 21476 12066
rect 21420 10050 21476 12014
rect 21588 10498 21644 10510
rect 21588 10446 21590 10498
rect 21642 10446 21644 10498
rect 21588 10388 21644 10446
rect 21588 10322 21644 10332
rect 21420 9998 21422 10050
rect 21474 9998 21476 10050
rect 21420 9986 21476 9998
rect 21756 10052 21812 13694
rect 21980 13188 22036 13198
rect 21980 13094 22036 13132
rect 21756 9986 21812 9996
rect 21980 10386 22036 10398
rect 21980 10334 21982 10386
rect 22034 10334 22036 10386
rect 20860 9826 21364 9828
rect 20860 9774 20862 9826
rect 20914 9774 21364 9826
rect 20860 9772 21364 9774
rect 21812 9828 21868 9838
rect 20860 9268 20916 9772
rect 21812 9734 21868 9772
rect 21980 9826 22036 10334
rect 21980 9774 21982 9826
rect 22034 9774 22036 9826
rect 21980 9762 22036 9774
rect 22092 9826 22148 9838
rect 22092 9774 22094 9826
rect 22146 9774 22148 9826
rect 20860 9202 20916 9212
rect 22092 8932 22148 9774
rect 22092 8866 22148 8876
rect 21980 8260 22036 8270
rect 21980 8166 22036 8204
rect 21588 8148 21644 8158
rect 21588 8054 21644 8092
rect 20972 8036 21028 8046
rect 20972 7530 21028 7980
rect 22204 8036 22260 18172
rect 22492 17276 22756 17286
rect 22548 17220 22596 17276
rect 22652 17220 22700 17276
rect 22492 17210 22756 17220
rect 22316 16996 22372 17006
rect 22316 16882 22372 16940
rect 22316 16830 22318 16882
rect 22370 16830 22372 16882
rect 22316 16212 22372 16830
rect 22316 16146 22372 16156
rect 22492 15708 22756 15718
rect 22548 15652 22596 15708
rect 22652 15652 22700 15708
rect 22492 15642 22756 15652
rect 22492 14140 22756 14150
rect 22548 14084 22596 14140
rect 22652 14084 22700 14140
rect 22492 14074 22756 14084
rect 22316 13300 22372 13310
rect 22316 12962 22372 13244
rect 22316 12910 22318 12962
rect 22370 12910 22372 12962
rect 22316 12898 22372 12910
rect 22492 12572 22756 12582
rect 22548 12516 22596 12572
rect 22652 12516 22700 12572
rect 22492 12506 22756 12516
rect 22492 11004 22756 11014
rect 22548 10948 22596 11004
rect 22652 10948 22700 11004
rect 22492 10938 22756 10948
rect 22316 10610 22372 10622
rect 22316 10558 22318 10610
rect 22370 10558 22372 10610
rect 22316 10388 22372 10558
rect 22316 10322 22372 10332
rect 22492 9436 22756 9446
rect 22548 9380 22596 9436
rect 22652 9380 22700 9436
rect 22492 9370 22756 9380
rect 22204 7970 22260 7980
rect 22316 8258 22372 8270
rect 22316 8206 22318 8258
rect 22370 8206 22372 8258
rect 22316 8148 22372 8206
rect 20972 7478 20974 7530
rect 21026 7478 21028 7530
rect 20972 7466 21028 7478
rect 22316 7476 22372 8092
rect 22492 7868 22756 7878
rect 22548 7812 22596 7868
rect 22652 7812 22700 7868
rect 22492 7802 22756 7812
rect 22316 7410 22372 7420
rect 22492 6300 22756 6310
rect 22548 6244 22596 6300
rect 22652 6244 22700 6300
rect 22492 6234 22756 6244
rect 20860 5796 20916 5806
rect 20860 5236 20916 5740
rect 20860 5122 20916 5180
rect 21980 5236 22036 5246
rect 21980 5142 22036 5180
rect 20860 5070 20862 5122
rect 20914 5070 20916 5122
rect 20860 4338 20916 5070
rect 21588 5124 21644 5134
rect 21588 5030 21644 5068
rect 22316 5124 22372 5134
rect 22316 4564 22372 5068
rect 22492 4732 22756 4742
rect 22548 4676 22596 4732
rect 22652 4676 22700 4732
rect 22492 4666 22756 4676
rect 22316 4498 22372 4508
rect 20860 4286 20862 4338
rect 20914 4286 20916 4338
rect 20860 4274 20916 4286
rect 21196 4340 21252 4350
rect 21196 4246 21252 4284
rect 21700 4340 21756 4350
rect 20748 4118 20750 4170
rect 20802 4118 20804 4170
rect 21700 4228 21756 4284
rect 21700 4226 21812 4228
rect 21700 4174 21702 4226
rect 21754 4174 21812 4226
rect 21700 4162 21812 4174
rect 20748 4106 20804 4118
rect 3872 3948 4136 3958
rect 3928 3892 3976 3948
rect 4032 3892 4080 3948
rect 3872 3882 4136 3892
rect 9192 3948 9456 3958
rect 9248 3892 9296 3948
rect 9352 3892 9400 3948
rect 9192 3882 9456 3892
rect 14512 3948 14776 3958
rect 14568 3892 14616 3948
rect 14672 3892 14720 3948
rect 14512 3882 14776 3892
rect 19832 3948 20096 3958
rect 19888 3892 19936 3948
rect 19992 3892 20040 3948
rect 19832 3882 20096 3892
rect 21756 3668 21812 4162
rect 22148 4226 22204 4238
rect 22148 4174 22150 4226
rect 22202 4174 22204 4226
rect 22148 3668 22204 4174
rect 21756 3612 22204 3668
rect 6532 3164 6796 3174
rect 6588 3108 6636 3164
rect 6692 3108 6740 3164
rect 6532 3098 6796 3108
rect 11852 3164 12116 3174
rect 11908 3108 11956 3164
rect 12012 3108 12060 3164
rect 11852 3098 12116 3108
rect 17172 3164 17436 3174
rect 17228 3108 17276 3164
rect 17332 3108 17380 3164
rect 17172 3098 17436 3108
rect 21756 1652 21812 3612
rect 22492 3164 22756 3174
rect 22548 3108 22596 3164
rect 22652 3108 22700 3164
rect 22492 3098 22756 3108
rect 21756 1586 21812 1596
<< via2 >>
rect 6532 20410 6588 20412
rect 6532 20358 6534 20410
rect 6534 20358 6586 20410
rect 6586 20358 6588 20410
rect 6532 20356 6588 20358
rect 6636 20410 6692 20412
rect 6636 20358 6638 20410
rect 6638 20358 6690 20410
rect 6690 20358 6692 20410
rect 6636 20356 6692 20358
rect 6740 20410 6796 20412
rect 6740 20358 6742 20410
rect 6742 20358 6794 20410
rect 6794 20358 6796 20410
rect 6740 20356 6796 20358
rect 11852 20410 11908 20412
rect 11852 20358 11854 20410
rect 11854 20358 11906 20410
rect 11906 20358 11908 20410
rect 11852 20356 11908 20358
rect 11956 20410 12012 20412
rect 11956 20358 11958 20410
rect 11958 20358 12010 20410
rect 12010 20358 12012 20410
rect 11956 20356 12012 20358
rect 12060 20410 12116 20412
rect 12060 20358 12062 20410
rect 12062 20358 12114 20410
rect 12114 20358 12116 20410
rect 12060 20356 12116 20358
rect 17172 20410 17228 20412
rect 17172 20358 17174 20410
rect 17174 20358 17226 20410
rect 17226 20358 17228 20410
rect 17172 20356 17228 20358
rect 17276 20410 17332 20412
rect 17276 20358 17278 20410
rect 17278 20358 17330 20410
rect 17330 20358 17332 20410
rect 17276 20356 17332 20358
rect 17380 20410 17436 20412
rect 17380 20358 17382 20410
rect 17382 20358 17434 20410
rect 17434 20358 17436 20410
rect 17380 20356 17436 20358
rect 20076 21980 20132 22036
rect 19852 20076 19908 20132
rect 20972 20130 21028 20132
rect 20972 20078 20974 20130
rect 20974 20078 21026 20130
rect 21026 20078 21028 20130
rect 20972 20076 21028 20078
rect 22492 20410 22548 20412
rect 22492 20358 22494 20410
rect 22494 20358 22546 20410
rect 22546 20358 22548 20410
rect 22492 20356 22548 20358
rect 22596 20410 22652 20412
rect 22596 20358 22598 20410
rect 22598 20358 22650 20410
rect 22650 20358 22652 20410
rect 22596 20356 22652 20358
rect 22700 20410 22756 20412
rect 22700 20358 22702 20410
rect 22702 20358 22754 20410
rect 22754 20358 22756 20410
rect 22700 20356 22756 20358
rect 5852 19964 5908 20020
rect 3872 19626 3928 19628
rect 3872 19574 3874 19626
rect 3874 19574 3926 19626
rect 3926 19574 3928 19626
rect 3872 19572 3928 19574
rect 3976 19626 4032 19628
rect 3976 19574 3978 19626
rect 3978 19574 4030 19626
rect 4030 19574 4032 19626
rect 3976 19572 4032 19574
rect 4080 19626 4136 19628
rect 4080 19574 4082 19626
rect 4082 19574 4134 19626
rect 4134 19574 4136 19626
rect 4080 19572 4136 19574
rect 4508 19458 4564 19460
rect 4508 19406 4510 19458
rect 4510 19406 4562 19458
rect 4562 19406 4564 19458
rect 4508 19404 4564 19406
rect 9212 20018 9268 20020
rect 9212 19966 9214 20018
rect 9214 19966 9266 20018
rect 9266 19966 9268 20018
rect 9212 19964 9268 19966
rect 9192 19626 9248 19628
rect 9192 19574 9194 19626
rect 9194 19574 9246 19626
rect 9246 19574 9248 19626
rect 9192 19572 9248 19574
rect 9296 19626 9352 19628
rect 9296 19574 9298 19626
rect 9298 19574 9350 19626
rect 9350 19574 9352 19626
rect 9296 19572 9352 19574
rect 9400 19626 9456 19628
rect 9400 19574 9402 19626
rect 9402 19574 9454 19626
rect 9454 19574 9456 19626
rect 9400 19572 9456 19574
rect 6412 19404 6468 19460
rect 3388 18508 3444 18564
rect 4060 19234 4116 19236
rect 4060 19182 4062 19234
rect 4062 19182 4114 19234
rect 4114 19182 4116 19234
rect 4060 19180 4116 19182
rect 5012 19180 5068 19236
rect 5180 19234 5236 19236
rect 5180 19182 5182 19234
rect 5182 19182 5234 19234
rect 5234 19182 5236 19234
rect 5180 19180 5236 19182
rect 3556 17948 3612 18004
rect 4508 18508 4564 18564
rect 3500 17724 3556 17780
rect 3872 18058 3928 18060
rect 3872 18006 3874 18058
rect 3874 18006 3926 18058
rect 3926 18006 3928 18058
rect 3872 18004 3928 18006
rect 3976 18058 4032 18060
rect 3976 18006 3978 18058
rect 3978 18006 4030 18058
rect 4030 18006 4032 18058
rect 3976 18004 4032 18006
rect 4080 18058 4136 18060
rect 4080 18006 4082 18058
rect 4082 18006 4134 18058
rect 4134 18006 4136 18058
rect 4080 18004 4136 18006
rect 6532 18842 6588 18844
rect 6532 18790 6534 18842
rect 6534 18790 6586 18842
rect 6586 18790 6588 18842
rect 6532 18788 6588 18790
rect 6636 18842 6692 18844
rect 6636 18790 6638 18842
rect 6638 18790 6690 18842
rect 6690 18790 6692 18842
rect 6636 18788 6692 18790
rect 6740 18842 6796 18844
rect 6740 18790 6742 18842
rect 6742 18790 6794 18842
rect 6794 18790 6796 18842
rect 6740 18788 6796 18790
rect 5516 18508 5572 18564
rect 7644 18508 7700 18564
rect 3948 17724 4004 17780
rect 3724 16882 3780 16884
rect 3724 16830 3726 16882
rect 3726 16830 3778 16882
rect 3778 16830 3780 16882
rect 3724 16828 3780 16830
rect 7756 18338 7812 18340
rect 7756 18286 7758 18338
rect 7758 18286 7810 18338
rect 7810 18286 7812 18338
rect 7756 18284 7812 18286
rect 3872 16490 3928 16492
rect 3872 16438 3874 16490
rect 3874 16438 3926 16490
rect 3926 16438 3928 16490
rect 3872 16436 3928 16438
rect 3976 16490 4032 16492
rect 3976 16438 3978 16490
rect 3978 16438 4030 16490
rect 4030 16438 4032 16490
rect 3976 16436 4032 16438
rect 4080 16490 4136 16492
rect 4080 16438 4082 16490
rect 4082 16438 4134 16490
rect 4134 16438 4136 16490
rect 4080 16436 4136 16438
rect 2828 15372 2884 15428
rect 3612 16044 3668 16100
rect 4508 17500 4564 17556
rect 4508 17052 4564 17108
rect 4844 17612 4900 17668
rect 3836 15372 3892 15428
rect 4396 16098 4452 16100
rect 4396 16046 4398 16098
rect 4398 16046 4450 16098
rect 4450 16046 4452 16098
rect 4396 16044 4452 16046
rect 3948 15260 4004 15316
rect 6532 17274 6588 17276
rect 6532 17222 6534 17274
rect 6534 17222 6586 17274
rect 6586 17222 6588 17274
rect 6532 17220 6588 17222
rect 6636 17274 6692 17276
rect 6636 17222 6638 17274
rect 6638 17222 6690 17274
rect 6690 17222 6692 17274
rect 6636 17220 6692 17222
rect 6740 17274 6796 17276
rect 6740 17222 6742 17274
rect 6742 17222 6794 17274
rect 6794 17222 6796 17274
rect 6740 17220 6796 17222
rect 4844 16882 4900 16884
rect 4844 16830 4846 16882
rect 4846 16830 4898 16882
rect 4898 16830 4900 16882
rect 4844 16828 4900 16830
rect 4732 16044 4788 16100
rect 4676 15260 4732 15316
rect 3872 14922 3928 14924
rect 3872 14870 3874 14922
rect 3874 14870 3926 14922
rect 3926 14870 3928 14922
rect 3872 14868 3928 14870
rect 3976 14922 4032 14924
rect 3976 14870 3978 14922
rect 3978 14870 4030 14922
rect 4030 14870 4032 14922
rect 3976 14868 4032 14870
rect 4080 14922 4136 14924
rect 4080 14870 4082 14922
rect 4082 14870 4134 14922
rect 4134 14870 4136 14922
rect 4080 14868 4136 14870
rect 4172 13858 4228 13860
rect 4172 13806 4174 13858
rect 4174 13806 4226 13858
rect 4226 13806 4228 13858
rect 4172 13804 4228 13806
rect 3872 13354 3928 13356
rect 3872 13302 3874 13354
rect 3874 13302 3926 13354
rect 3926 13302 3928 13354
rect 3872 13300 3928 13302
rect 3976 13354 4032 13356
rect 3976 13302 3978 13354
rect 3978 13302 4030 13354
rect 4030 13302 4032 13354
rect 3976 13300 4032 13302
rect 4080 13354 4136 13356
rect 4080 13302 4082 13354
rect 4082 13302 4134 13354
rect 4134 13302 4136 13354
rect 4080 13300 4136 13302
rect 4284 13020 4340 13076
rect 3872 11786 3928 11788
rect 3872 11734 3874 11786
rect 3874 11734 3926 11786
rect 3926 11734 3928 11786
rect 3872 11732 3928 11734
rect 3976 11786 4032 11788
rect 3976 11734 3978 11786
rect 3978 11734 4030 11786
rect 4030 11734 4032 11786
rect 3976 11732 4032 11734
rect 4080 11786 4136 11788
rect 4080 11734 4082 11786
rect 4082 11734 4134 11786
rect 4134 11734 4136 11786
rect 4080 11732 4136 11734
rect 3164 11394 3220 11396
rect 3164 11342 3166 11394
rect 3166 11342 3218 11394
rect 3218 11342 3220 11394
rect 3164 11340 3220 11342
rect 3948 11340 4004 11396
rect 7980 16940 8036 16996
rect 7532 16044 7588 16100
rect 6532 15706 6588 15708
rect 6532 15654 6534 15706
rect 6534 15654 6586 15706
rect 6586 15654 6588 15706
rect 6532 15652 6588 15654
rect 6636 15706 6692 15708
rect 6636 15654 6638 15706
rect 6638 15654 6690 15706
rect 6690 15654 6692 15706
rect 6636 15652 6692 15654
rect 6740 15706 6796 15708
rect 6740 15654 6742 15706
rect 6742 15654 6794 15706
rect 6794 15654 6796 15706
rect 6740 15652 6796 15654
rect 4620 14252 4676 14308
rect 5180 14588 5236 14644
rect 4508 13020 4564 13076
rect 3872 10218 3928 10220
rect 3872 10166 3874 10218
rect 3874 10166 3926 10218
rect 3926 10166 3928 10218
rect 3872 10164 3928 10166
rect 3976 10218 4032 10220
rect 3976 10166 3978 10218
rect 3978 10166 4030 10218
rect 4030 10166 4032 10218
rect 3976 10164 4032 10166
rect 4080 10218 4136 10220
rect 4080 10166 4082 10218
rect 4082 10166 4134 10218
rect 4134 10166 4136 10218
rect 4080 10164 4136 10166
rect 4508 11367 4564 11396
rect 4508 11340 4510 11367
rect 4510 11340 4562 11367
rect 4562 11340 4564 11367
rect 3724 9884 3780 9940
rect 3872 8650 3928 8652
rect 3872 8598 3874 8650
rect 3874 8598 3926 8650
rect 3926 8598 3928 8650
rect 3872 8596 3928 8598
rect 3976 8650 4032 8652
rect 3976 8598 3978 8650
rect 3978 8598 4030 8650
rect 4030 8598 4032 8650
rect 3976 8596 4032 8598
rect 4080 8650 4136 8652
rect 4080 8598 4082 8650
rect 4082 8598 4134 8650
rect 4134 8598 4136 8650
rect 4080 8596 4136 8598
rect 4396 9714 4452 9716
rect 4396 9662 4398 9714
rect 4398 9662 4450 9714
rect 4450 9662 4452 9714
rect 4396 9660 4452 9662
rect 4844 13746 4900 13748
rect 4844 13694 4846 13746
rect 4846 13694 4898 13746
rect 4898 13694 4900 13746
rect 4844 13692 4900 13694
rect 4844 9884 4900 9940
rect 4732 9772 4788 9828
rect 5796 14642 5852 14644
rect 5796 14590 5798 14642
rect 5798 14590 5850 14642
rect 5850 14590 5852 14642
rect 5796 14588 5852 14590
rect 5684 14252 5740 14308
rect 6532 14138 6588 14140
rect 6532 14086 6534 14138
rect 6534 14086 6586 14138
rect 6586 14086 6588 14138
rect 6532 14084 6588 14086
rect 6636 14138 6692 14140
rect 6636 14086 6638 14138
rect 6638 14086 6690 14138
rect 6690 14086 6692 14138
rect 6636 14084 6692 14086
rect 6740 14138 6796 14140
rect 6740 14086 6742 14138
rect 6742 14086 6794 14138
rect 6794 14086 6796 14138
rect 6740 14084 6796 14086
rect 4732 8876 4788 8932
rect 4508 8316 4564 8372
rect 3892 7644 3948 7700
rect 4620 8258 4676 8260
rect 4620 8206 4622 8258
rect 4622 8206 4674 8258
rect 4674 8206 4676 8258
rect 4620 8204 4676 8206
rect 4676 7698 4732 7700
rect 4676 7646 4678 7698
rect 4678 7646 4730 7698
rect 4730 7646 4732 7698
rect 4676 7644 4732 7646
rect 4508 7474 4564 7476
rect 4508 7422 4510 7474
rect 4510 7422 4562 7474
rect 4562 7422 4564 7474
rect 4508 7420 4564 7422
rect 3872 7082 3928 7084
rect 3872 7030 3874 7082
rect 3874 7030 3926 7082
rect 3926 7030 3928 7082
rect 3872 7028 3928 7030
rect 3976 7082 4032 7084
rect 3976 7030 3978 7082
rect 3978 7030 4030 7082
rect 4030 7030 4032 7082
rect 3976 7028 4032 7030
rect 4080 7082 4136 7084
rect 4080 7030 4082 7082
rect 4082 7030 4134 7082
rect 4134 7030 4136 7082
rect 4080 7028 4136 7030
rect 3855 5852 3911 5908
rect 4956 9212 5012 9268
rect 5124 8370 5180 8372
rect 5124 8318 5126 8370
rect 5126 8318 5178 8370
rect 5178 8318 5180 8370
rect 5124 8316 5180 8318
rect 8652 18508 8708 18564
rect 11852 18842 11908 18844
rect 11852 18790 11854 18842
rect 11854 18790 11906 18842
rect 11906 18790 11908 18842
rect 11852 18788 11908 18790
rect 11956 18842 12012 18844
rect 11956 18790 11958 18842
rect 11958 18790 12010 18842
rect 12010 18790 12012 18842
rect 11956 18788 12012 18790
rect 12060 18842 12116 18844
rect 12060 18790 12062 18842
rect 12062 18790 12114 18842
rect 12114 18790 12116 18842
rect 12060 18788 12116 18790
rect 9436 18508 9492 18564
rect 9996 18450 10052 18452
rect 9996 18398 9998 18450
rect 9998 18398 10050 18450
rect 10050 18398 10052 18450
rect 9996 18396 10052 18398
rect 9660 18284 9716 18340
rect 9192 18058 9248 18060
rect 9192 18006 9194 18058
rect 9194 18006 9246 18058
rect 9246 18006 9248 18058
rect 9192 18004 9248 18006
rect 9296 18058 9352 18060
rect 9296 18006 9298 18058
rect 9298 18006 9350 18058
rect 9350 18006 9352 18058
rect 9296 18004 9352 18006
rect 9400 18058 9456 18060
rect 9400 18006 9402 18058
rect 9402 18006 9454 18058
rect 9454 18006 9456 18058
rect 9400 18004 9456 18006
rect 8876 17666 8932 17668
rect 8876 17614 8878 17666
rect 8878 17614 8930 17666
rect 8930 17614 8932 17666
rect 8876 17612 8932 17614
rect 8484 17388 8540 17444
rect 8484 16940 8540 16996
rect 8876 16940 8932 16996
rect 14512 19626 14568 19628
rect 14512 19574 14514 19626
rect 14514 19574 14566 19626
rect 14566 19574 14568 19626
rect 14512 19572 14568 19574
rect 14616 19626 14672 19628
rect 14616 19574 14618 19626
rect 14618 19574 14670 19626
rect 14670 19574 14672 19626
rect 14616 19572 14672 19574
rect 14720 19626 14776 19628
rect 14720 19574 14722 19626
rect 14722 19574 14774 19626
rect 14774 19574 14776 19626
rect 14720 19572 14776 19574
rect 16380 19458 16436 19460
rect 16380 19406 16382 19458
rect 16382 19406 16434 19458
rect 16434 19406 16436 19458
rect 16380 19404 16436 19406
rect 17612 19404 17668 19460
rect 18620 19458 18676 19460
rect 18620 19406 18622 19458
rect 18622 19406 18674 19458
rect 18674 19406 18676 19458
rect 18620 19404 18676 19406
rect 14252 19180 14308 19236
rect 14140 18956 14196 19012
rect 14924 18956 14980 19012
rect 14028 18450 14084 18452
rect 14028 18398 14030 18450
rect 14030 18398 14082 18450
rect 14082 18398 14084 18450
rect 14028 18396 14084 18398
rect 13692 18284 13748 18340
rect 13860 18172 13916 18228
rect 14700 18172 14756 18228
rect 14512 18058 14568 18060
rect 14512 18006 14514 18058
rect 14514 18006 14566 18058
rect 14566 18006 14568 18058
rect 14512 18004 14568 18006
rect 14616 18058 14672 18060
rect 14616 18006 14618 18058
rect 14618 18006 14670 18058
rect 14670 18006 14672 18058
rect 14616 18004 14672 18006
rect 14720 18058 14776 18060
rect 14720 18006 14722 18058
rect 14722 18006 14774 18058
rect 14774 18006 14776 18058
rect 14720 18004 14776 18006
rect 12684 17612 12740 17668
rect 11852 17274 11908 17276
rect 11852 17222 11854 17274
rect 11854 17222 11906 17274
rect 11906 17222 11908 17274
rect 11852 17220 11908 17222
rect 11956 17274 12012 17276
rect 11956 17222 11958 17274
rect 11958 17222 12010 17274
rect 12010 17222 12012 17274
rect 11956 17220 12012 17222
rect 12060 17274 12116 17276
rect 12060 17222 12062 17274
rect 12062 17222 12114 17274
rect 12114 17222 12116 17274
rect 12060 17220 12116 17222
rect 11676 17052 11732 17108
rect 9192 16490 9248 16492
rect 9192 16438 9194 16490
rect 9194 16438 9246 16490
rect 9246 16438 9248 16490
rect 9192 16436 9248 16438
rect 9296 16490 9352 16492
rect 9296 16438 9298 16490
rect 9298 16438 9350 16490
rect 9350 16438 9352 16490
rect 9296 16436 9352 16438
rect 9400 16490 9456 16492
rect 9400 16438 9402 16490
rect 9402 16438 9454 16490
rect 9454 16438 9456 16490
rect 9400 16436 9456 16438
rect 8092 16044 8148 16100
rect 9192 14922 9248 14924
rect 9192 14870 9194 14922
rect 9194 14870 9246 14922
rect 9246 14870 9248 14922
rect 9192 14868 9248 14870
rect 9296 14922 9352 14924
rect 9296 14870 9298 14922
rect 9298 14870 9350 14922
rect 9350 14870 9352 14922
rect 9296 14868 9352 14870
rect 9400 14922 9456 14924
rect 9400 14870 9402 14922
rect 9402 14870 9454 14922
rect 9454 14870 9456 14922
rect 9400 14868 9456 14870
rect 7980 14588 8036 14644
rect 7196 13804 7252 13860
rect 8092 13804 8148 13860
rect 7308 13692 7364 13748
rect 7420 13468 7476 13524
rect 7868 13132 7924 13188
rect 6532 12570 6588 12572
rect 6532 12518 6534 12570
rect 6534 12518 6586 12570
rect 6586 12518 6588 12570
rect 6532 12516 6588 12518
rect 6636 12570 6692 12572
rect 6636 12518 6638 12570
rect 6638 12518 6690 12570
rect 6690 12518 6692 12570
rect 6636 12516 6692 12518
rect 6740 12570 6796 12572
rect 6740 12518 6742 12570
rect 6742 12518 6794 12570
rect 6794 12518 6796 12570
rect 6740 12516 6796 12518
rect 6532 11002 6588 11004
rect 6532 10950 6534 11002
rect 6534 10950 6586 11002
rect 6586 10950 6588 11002
rect 6532 10948 6588 10950
rect 6636 11002 6692 11004
rect 6636 10950 6638 11002
rect 6638 10950 6690 11002
rect 6690 10950 6692 11002
rect 6636 10948 6692 10950
rect 6740 11002 6796 11004
rect 6740 10950 6742 11002
rect 6742 10950 6794 11002
rect 6794 10950 6796 11002
rect 6740 10948 6796 10950
rect 6300 9938 6356 9940
rect 6300 9886 6302 9938
rect 6302 9886 6354 9938
rect 6354 9886 6356 9938
rect 6300 9884 6356 9886
rect 6076 9660 6132 9716
rect 6468 9660 6524 9716
rect 6916 9714 6972 9716
rect 6916 9662 6918 9714
rect 6918 9662 6970 9714
rect 6970 9662 6972 9714
rect 6916 9660 6972 9662
rect 6532 9434 6588 9436
rect 6532 9382 6534 9434
rect 6534 9382 6586 9434
rect 6586 9382 6588 9434
rect 6532 9380 6588 9382
rect 6636 9434 6692 9436
rect 6636 9382 6638 9434
rect 6638 9382 6690 9434
rect 6690 9382 6692 9434
rect 6636 9380 6692 9382
rect 6740 9434 6796 9436
rect 6740 9382 6742 9434
rect 6742 9382 6794 9434
rect 6794 9382 6796 9434
rect 6740 9380 6796 9382
rect 6076 8988 6132 9044
rect 8316 13132 8372 13188
rect 11340 16882 11396 16884
rect 11340 16830 11342 16882
rect 11342 16830 11394 16882
rect 11394 16830 11396 16882
rect 11340 16828 11396 16830
rect 12236 17052 12292 17108
rect 12012 16863 12014 16884
rect 12014 16863 12066 16884
rect 12066 16863 12068 16884
rect 13580 17666 13636 17668
rect 13580 17614 13582 17666
rect 13582 17614 13634 17666
rect 13634 17614 13636 17666
rect 13580 17612 13636 17614
rect 13132 16994 13188 16996
rect 13132 16942 13134 16994
rect 13134 16942 13186 16994
rect 13186 16942 13188 16994
rect 13132 16940 13188 16942
rect 12012 16828 12068 16863
rect 11852 15706 11908 15708
rect 11852 15654 11854 15706
rect 11854 15654 11906 15706
rect 11906 15654 11908 15706
rect 11852 15652 11908 15654
rect 11956 15706 12012 15708
rect 11956 15654 11958 15706
rect 11958 15654 12010 15706
rect 12010 15654 12012 15706
rect 11956 15652 12012 15654
rect 12060 15706 12116 15708
rect 12060 15654 12062 15706
rect 12062 15654 12114 15706
rect 12114 15654 12116 15706
rect 12060 15652 12116 15654
rect 12796 16828 12852 16884
rect 11852 14138 11908 14140
rect 11852 14086 11854 14138
rect 11854 14086 11906 14138
rect 11906 14086 11908 14138
rect 11852 14084 11908 14086
rect 11956 14138 12012 14140
rect 11956 14086 11958 14138
rect 11958 14086 12010 14138
rect 12010 14086 12012 14138
rect 11956 14084 12012 14086
rect 12060 14138 12116 14140
rect 12060 14086 12062 14138
rect 12062 14086 12114 14138
rect 12114 14086 12116 14138
rect 12060 14084 12116 14086
rect 11116 13916 11172 13972
rect 8764 13746 8820 13748
rect 8764 13694 8766 13746
rect 8766 13694 8818 13746
rect 8818 13694 8820 13746
rect 8764 13692 8820 13694
rect 9996 13468 10052 13524
rect 9192 13354 9248 13356
rect 9192 13302 9194 13354
rect 9194 13302 9246 13354
rect 9246 13302 9248 13354
rect 9192 13300 9248 13302
rect 9296 13354 9352 13356
rect 9296 13302 9298 13354
rect 9298 13302 9350 13354
rect 9350 13302 9352 13354
rect 9296 13300 9352 13302
rect 9400 13354 9456 13356
rect 9400 13302 9402 13354
rect 9402 13302 9454 13354
rect 9454 13302 9456 13354
rect 9400 13300 9456 13302
rect 8428 12348 8484 12404
rect 9884 12796 9940 12852
rect 8876 12684 8932 12740
rect 9772 12684 9828 12740
rect 8764 12236 8820 12292
rect 8876 12348 8932 12404
rect 7532 12124 7588 12180
rect 8652 12141 8654 12180
rect 8654 12141 8706 12180
rect 8706 12141 8708 12180
rect 8652 12124 8708 12141
rect 9192 11786 9248 11788
rect 9192 11734 9194 11786
rect 9194 11734 9246 11786
rect 9246 11734 9248 11786
rect 9192 11732 9248 11734
rect 9296 11786 9352 11788
rect 9296 11734 9298 11786
rect 9298 11734 9350 11786
rect 9350 11734 9352 11786
rect 9296 11732 9352 11734
rect 9400 11786 9456 11788
rect 9400 11734 9402 11786
rect 9402 11734 9454 11786
rect 9454 11734 9456 11786
rect 9400 11732 9456 11734
rect 9192 10218 9248 10220
rect 9192 10166 9194 10218
rect 9194 10166 9246 10218
rect 9246 10166 9248 10218
rect 9192 10164 9248 10166
rect 9296 10218 9352 10220
rect 9296 10166 9298 10218
rect 9298 10166 9350 10218
rect 9350 10166 9352 10218
rect 9296 10164 9352 10166
rect 9400 10218 9456 10220
rect 9400 10166 9402 10218
rect 9402 10166 9454 10218
rect 9454 10166 9456 10218
rect 9400 10164 9456 10166
rect 8204 9826 8260 9828
rect 8204 9774 8206 9826
rect 8206 9774 8258 9826
rect 8258 9774 8260 9826
rect 8204 9772 8260 9774
rect 6972 9212 7028 9268
rect 7980 9660 8036 9716
rect 5684 8316 5740 8372
rect 5796 8204 5852 8260
rect 6532 7866 6588 7868
rect 6532 7814 6534 7866
rect 6534 7814 6586 7866
rect 6586 7814 6588 7866
rect 6532 7812 6588 7814
rect 6636 7866 6692 7868
rect 6636 7814 6638 7866
rect 6638 7814 6690 7866
rect 6690 7814 6692 7866
rect 6636 7812 6692 7814
rect 6740 7866 6796 7868
rect 6740 7814 6742 7866
rect 6742 7814 6794 7866
rect 6794 7814 6796 7866
rect 6740 7812 6796 7814
rect 4956 7420 5012 7476
rect 3612 5516 3668 5572
rect 3872 5514 3928 5516
rect 3872 5462 3874 5514
rect 3874 5462 3926 5514
rect 3926 5462 3928 5514
rect 3872 5460 3928 5462
rect 3976 5514 4032 5516
rect 3976 5462 3978 5514
rect 3978 5462 4030 5514
rect 4030 5462 4032 5514
rect 3976 5460 4032 5462
rect 4080 5514 4136 5516
rect 4080 5462 4082 5514
rect 4082 5462 4134 5514
rect 4134 5462 4136 5514
rect 4080 5460 4136 5462
rect 3612 5068 3668 5124
rect 4620 5122 4676 5124
rect 3052 4844 3108 4900
rect 4620 5070 4622 5122
rect 4622 5070 4674 5122
rect 4674 5070 4676 5122
rect 4620 5068 4676 5070
rect 5236 7474 5292 7476
rect 5236 7422 5238 7474
rect 5238 7422 5290 7474
rect 5290 7422 5292 7474
rect 5236 7420 5292 7422
rect 6532 6298 6588 6300
rect 6532 6246 6534 6298
rect 6534 6246 6586 6298
rect 6586 6246 6588 6298
rect 6532 6244 6588 6246
rect 6636 6298 6692 6300
rect 6636 6246 6638 6298
rect 6638 6246 6690 6298
rect 6690 6246 6692 6298
rect 6636 6244 6692 6246
rect 6740 6298 6796 6300
rect 6740 6246 6742 6298
rect 6742 6246 6794 6298
rect 6794 6246 6796 6298
rect 6740 6244 6796 6246
rect 6804 5906 6860 5908
rect 6804 5854 6806 5906
rect 6806 5854 6858 5906
rect 6858 5854 6860 5906
rect 6804 5852 6860 5854
rect 7420 9042 7476 9044
rect 7420 8990 7422 9042
rect 7422 8990 7474 9042
rect 7474 8990 7476 9042
rect 7420 8988 7476 8990
rect 7420 8316 7476 8372
rect 7196 8204 7252 8260
rect 7084 5906 7140 5908
rect 7084 5854 7086 5906
rect 7086 5854 7138 5906
rect 7138 5854 7140 5906
rect 7084 5852 7140 5854
rect 7644 7644 7700 7700
rect 7868 8988 7924 9044
rect 8428 9324 8484 9380
rect 8204 8876 8260 8932
rect 7980 6300 8036 6356
rect 8204 6662 8260 6692
rect 8204 6636 8206 6662
rect 8206 6636 8258 6662
rect 8258 6636 8260 6662
rect 8428 8764 8484 8820
rect 8652 9324 8708 9380
rect 8540 9100 8596 9156
rect 10332 12348 10388 12404
rect 9884 12178 9940 12180
rect 9884 12126 9886 12178
rect 9886 12126 9938 12178
rect 9938 12126 9940 12178
rect 9884 12124 9940 12126
rect 10164 12178 10220 12180
rect 10164 12126 10166 12178
rect 10166 12126 10218 12178
rect 10218 12126 10220 12178
rect 10164 12124 10220 12126
rect 8652 8876 8708 8932
rect 8540 8428 8596 8484
rect 9044 8876 9100 8932
rect 9192 8650 9248 8652
rect 9192 8598 9194 8650
rect 9194 8598 9246 8650
rect 9246 8598 9248 8650
rect 9192 8596 9248 8598
rect 9296 8650 9352 8652
rect 9296 8598 9298 8650
rect 9298 8598 9350 8650
rect 9350 8598 9352 8650
rect 9296 8596 9352 8598
rect 9400 8650 9456 8652
rect 9400 8598 9402 8650
rect 9402 8598 9454 8650
rect 9454 8598 9456 8650
rect 9400 8596 9456 8598
rect 9324 8428 9380 8484
rect 8204 6300 8260 6356
rect 7308 5628 7364 5684
rect 6748 5094 6804 5124
rect 6748 5068 6750 5094
rect 6750 5068 6802 5094
rect 6802 5068 6804 5094
rect 4956 4844 5012 4900
rect 6532 4730 6588 4732
rect 6532 4678 6534 4730
rect 6534 4678 6586 4730
rect 6586 4678 6588 4730
rect 6532 4676 6588 4678
rect 6636 4730 6692 4732
rect 6636 4678 6638 4730
rect 6638 4678 6690 4730
rect 6690 4678 6692 4730
rect 6636 4676 6692 4678
rect 6740 4730 6796 4732
rect 6740 4678 6742 4730
rect 6742 4678 6794 4730
rect 6794 4678 6796 4730
rect 6740 4676 6796 4678
rect 7812 5682 7868 5684
rect 7812 5630 7814 5682
rect 7814 5630 7866 5682
rect 7866 5630 7868 5682
rect 7812 5628 7868 5630
rect 7196 5122 7252 5124
rect 7196 5070 7198 5122
rect 7198 5070 7250 5122
rect 7250 5070 7252 5122
rect 7644 5180 7700 5236
rect 7196 5068 7252 5070
rect 8204 5852 8260 5908
rect 7980 5292 8036 5348
rect 7756 4956 7812 5012
rect 7084 4508 7140 4564
rect 7756 4562 7812 4564
rect 7756 4510 7758 4562
rect 7758 4510 7810 4562
rect 7810 4510 7812 4562
rect 7756 4508 7812 4510
rect 9548 8428 9604 8484
rect 9268 7644 9324 7700
rect 9192 7082 9248 7084
rect 9192 7030 9194 7082
rect 9194 7030 9246 7082
rect 9246 7030 9248 7082
rect 9192 7028 9248 7030
rect 9296 7082 9352 7084
rect 9296 7030 9298 7082
rect 9298 7030 9350 7082
rect 9350 7030 9352 7082
rect 9296 7028 9352 7030
rect 9400 7082 9456 7084
rect 9400 7030 9402 7082
rect 9402 7030 9454 7082
rect 9454 7030 9456 7082
rect 9400 7028 9456 7030
rect 10780 9100 10836 9156
rect 10220 9042 10276 9044
rect 10220 8990 10222 9042
rect 10222 8990 10274 9042
rect 10274 8990 10276 9042
rect 10220 8988 10276 8990
rect 11788 13916 11844 13972
rect 12012 13916 12068 13972
rect 12572 14476 12628 14532
rect 12572 13916 12628 13972
rect 11676 13020 11732 13076
rect 11564 12402 11620 12404
rect 11564 12350 11566 12402
rect 11566 12350 11618 12402
rect 11618 12350 11620 12402
rect 11564 12348 11620 12350
rect 12236 13244 12292 13300
rect 12796 13244 12852 13300
rect 12124 13132 12180 13188
rect 12348 13074 12404 13076
rect 12348 13022 12350 13074
rect 12350 13022 12402 13074
rect 12402 13022 12404 13074
rect 12348 13020 12404 13022
rect 12236 12947 12292 12964
rect 12236 12908 12238 12947
rect 12238 12908 12290 12947
rect 12290 12908 12292 12947
rect 11852 12570 11908 12572
rect 11852 12518 11854 12570
rect 11854 12518 11906 12570
rect 11906 12518 11908 12570
rect 11852 12516 11908 12518
rect 11956 12570 12012 12572
rect 11956 12518 11958 12570
rect 11958 12518 12010 12570
rect 12010 12518 12012 12570
rect 11956 12516 12012 12518
rect 12060 12570 12116 12572
rect 12060 12518 12062 12570
rect 12062 12518 12114 12570
rect 12114 12518 12116 12570
rect 12060 12516 12116 12518
rect 12236 12178 12292 12180
rect 12236 12126 12238 12178
rect 12238 12126 12290 12178
rect 12290 12126 12292 12178
rect 12236 12124 12292 12126
rect 11852 11002 11908 11004
rect 11852 10950 11854 11002
rect 11854 10950 11906 11002
rect 11906 10950 11908 11002
rect 11852 10948 11908 10950
rect 11956 11002 12012 11004
rect 11956 10950 11958 11002
rect 11958 10950 12010 11002
rect 12010 10950 12012 11002
rect 11956 10948 12012 10950
rect 12060 11002 12116 11004
rect 12060 10950 12062 11002
rect 12062 10950 12114 11002
rect 12114 10950 12116 11002
rect 12060 10948 12116 10950
rect 11852 9434 11908 9436
rect 11852 9382 11854 9434
rect 11854 9382 11906 9434
rect 11906 9382 11908 9434
rect 11852 9380 11908 9382
rect 11956 9434 12012 9436
rect 11956 9382 11958 9434
rect 11958 9382 12010 9434
rect 12010 9382 12012 9434
rect 11956 9380 12012 9382
rect 12060 9434 12116 9436
rect 12060 9382 12062 9434
rect 12062 9382 12114 9434
rect 12114 9382 12116 9434
rect 12060 9380 12116 9382
rect 12684 9100 12740 9156
rect 10892 8316 10948 8372
rect 9996 6636 10052 6692
rect 8876 5852 8932 5908
rect 9192 5514 9248 5516
rect 9192 5462 9194 5514
rect 9194 5462 9246 5514
rect 9246 5462 9248 5514
rect 9192 5460 9248 5462
rect 9296 5514 9352 5516
rect 9296 5462 9298 5514
rect 9298 5462 9350 5514
rect 9350 5462 9352 5514
rect 9296 5460 9352 5462
rect 9400 5514 9456 5516
rect 9400 5462 9402 5514
rect 9402 5462 9454 5514
rect 9454 5462 9456 5514
rect 9400 5460 9456 5462
rect 9604 5292 9660 5348
rect 8652 5180 8708 5236
rect 9212 5180 9268 5236
rect 10668 5122 10724 5124
rect 10668 5070 10670 5122
rect 10670 5070 10722 5122
rect 10722 5070 10724 5122
rect 10668 5068 10724 5070
rect 11284 8930 11340 8932
rect 11284 8878 11286 8930
rect 11286 8878 11338 8930
rect 11338 8878 11340 8930
rect 11284 8876 11340 8878
rect 12124 8876 12180 8932
rect 12236 8428 12292 8484
rect 11852 7866 11908 7868
rect 11852 7814 11854 7866
rect 11854 7814 11906 7866
rect 11906 7814 11908 7866
rect 11852 7812 11908 7814
rect 11956 7866 12012 7868
rect 11956 7814 11958 7866
rect 11958 7814 12010 7866
rect 12010 7814 12012 7866
rect 11956 7812 12012 7814
rect 12060 7866 12116 7868
rect 12060 7814 12062 7866
rect 12062 7814 12114 7866
rect 12114 7814 12116 7866
rect 12060 7812 12116 7814
rect 11116 6636 11172 6692
rect 11852 6298 11908 6300
rect 11852 6246 11854 6298
rect 11854 6246 11906 6298
rect 11906 6246 11908 6298
rect 11852 6244 11908 6246
rect 11956 6298 12012 6300
rect 11956 6246 11958 6298
rect 11958 6246 12010 6298
rect 12010 6246 12012 6298
rect 11956 6244 12012 6246
rect 12060 6298 12116 6300
rect 12060 6246 12062 6298
rect 12062 6246 12114 6298
rect 12114 6246 12116 6298
rect 12060 6244 12116 6246
rect 11228 5068 11284 5124
rect 8708 4956 8764 5012
rect 11564 5292 11620 5348
rect 11676 5068 11732 5124
rect 11340 4844 11396 4900
rect 14364 17666 14420 17668
rect 14364 17614 14366 17666
rect 14366 17614 14418 17666
rect 14418 17614 14420 17666
rect 14364 17612 14420 17614
rect 15764 19010 15820 19012
rect 15764 18958 15766 19010
rect 15766 18958 15818 19010
rect 15818 18958 15820 19010
rect 15764 18956 15820 18958
rect 17172 18842 17228 18844
rect 17172 18790 17174 18842
rect 17174 18790 17226 18842
rect 17226 18790 17228 18842
rect 17172 18788 17228 18790
rect 17276 18842 17332 18844
rect 17276 18790 17278 18842
rect 17278 18790 17330 18842
rect 17330 18790 17332 18842
rect 17276 18788 17332 18790
rect 17380 18842 17436 18844
rect 17380 18790 17382 18842
rect 17382 18790 17434 18842
rect 17434 18790 17436 18842
rect 17380 18788 17436 18790
rect 16044 18396 16100 18452
rect 14924 17388 14980 17444
rect 14512 16490 14568 16492
rect 14512 16438 14514 16490
rect 14514 16438 14566 16490
rect 14566 16438 14568 16490
rect 14512 16436 14568 16438
rect 14616 16490 14672 16492
rect 14616 16438 14618 16490
rect 14618 16438 14670 16490
rect 14670 16438 14672 16490
rect 14616 16436 14672 16438
rect 14720 16490 14776 16492
rect 14720 16438 14722 16490
rect 14722 16438 14774 16490
rect 14774 16438 14776 16490
rect 14720 16436 14776 16438
rect 17172 17274 17228 17276
rect 17172 17222 17174 17274
rect 17174 17222 17226 17274
rect 17226 17222 17228 17274
rect 17172 17220 17228 17222
rect 17276 17274 17332 17276
rect 17276 17222 17278 17274
rect 17278 17222 17330 17274
rect 17330 17222 17332 17274
rect 17276 17220 17332 17222
rect 17380 17274 17436 17276
rect 17380 17222 17382 17274
rect 17382 17222 17434 17274
rect 17434 17222 17436 17274
rect 17380 17220 17436 17222
rect 14252 16098 14308 16100
rect 14252 16046 14254 16098
rect 14254 16046 14306 16098
rect 14306 16046 14308 16098
rect 14252 16044 14308 16046
rect 13916 15036 13972 15092
rect 13804 14530 13860 14532
rect 13804 14478 13806 14530
rect 13806 14478 13858 14530
rect 13858 14478 13860 14530
rect 13804 14476 13860 14478
rect 13356 14252 13412 14308
rect 13524 13522 13580 13524
rect 13524 13470 13526 13522
rect 13526 13470 13578 13522
rect 13578 13470 13580 13522
rect 13524 13468 13580 13470
rect 13524 12850 13580 12852
rect 13524 12798 13526 12850
rect 13526 12798 13578 12850
rect 13578 12798 13580 12850
rect 13524 12796 13580 12798
rect 13244 12348 13300 12404
rect 13804 13132 13860 13188
rect 14252 13692 14308 13748
rect 14028 13020 14084 13076
rect 14140 13468 14196 13524
rect 14028 12684 14084 12740
rect 13692 12124 13748 12180
rect 14924 16098 14980 16100
rect 14924 16046 14926 16098
rect 14926 16046 14978 16098
rect 14978 16046 14980 16098
rect 14924 16044 14980 16046
rect 14924 15277 14926 15316
rect 14926 15277 14978 15316
rect 14978 15277 14980 15316
rect 14924 15260 14980 15277
rect 14812 15036 14868 15092
rect 17172 15706 17228 15708
rect 17172 15654 17174 15706
rect 17174 15654 17226 15706
rect 17226 15654 17228 15706
rect 17172 15652 17228 15654
rect 17276 15706 17332 15708
rect 17276 15654 17278 15706
rect 17278 15654 17330 15706
rect 17330 15654 17332 15706
rect 17276 15652 17332 15654
rect 17380 15706 17436 15708
rect 17380 15654 17382 15706
rect 17382 15654 17434 15706
rect 17434 15654 17436 15706
rect 17380 15652 17436 15654
rect 14512 14922 14568 14924
rect 14512 14870 14514 14922
rect 14514 14870 14566 14922
rect 14566 14870 14568 14922
rect 14512 14868 14568 14870
rect 14616 14922 14672 14924
rect 14616 14870 14618 14922
rect 14618 14870 14670 14922
rect 14670 14870 14672 14922
rect 14616 14868 14672 14870
rect 14720 14922 14776 14924
rect 14720 14870 14722 14922
rect 14722 14870 14774 14922
rect 14774 14870 14776 14922
rect 14720 14868 14776 14870
rect 14512 13354 14568 13356
rect 14512 13302 14514 13354
rect 14514 13302 14566 13354
rect 14566 13302 14568 13354
rect 14512 13300 14568 13302
rect 14616 13354 14672 13356
rect 14616 13302 14618 13354
rect 14618 13302 14670 13354
rect 14670 13302 14672 13354
rect 14616 13300 14672 13302
rect 14720 13354 14776 13356
rect 14720 13302 14722 13354
rect 14722 13302 14774 13354
rect 14774 13302 14776 13354
rect 14720 13300 14776 13302
rect 14364 12947 14420 12964
rect 14364 12908 14366 12947
rect 14366 12908 14418 12947
rect 14418 12908 14420 12947
rect 14588 13132 14644 13188
rect 14588 12908 14644 12964
rect 14476 12572 14532 12628
rect 14700 11900 14756 11956
rect 13024 9100 13080 9156
rect 13356 6860 13412 6916
rect 13580 6636 13636 6692
rect 11900 5292 11956 5348
rect 12012 5068 12068 5124
rect 12348 5628 12404 5684
rect 13524 5740 13580 5796
rect 12684 5292 12740 5348
rect 12348 5180 12404 5236
rect 12572 5180 12628 5236
rect 12236 5122 12292 5124
rect 12236 5070 12238 5122
rect 12238 5070 12290 5122
rect 12290 5070 12292 5122
rect 12236 5068 12292 5070
rect 14028 9212 14084 9268
rect 13916 9100 13972 9156
rect 13804 9018 13806 9044
rect 13806 9018 13858 9044
rect 13858 9018 13860 9044
rect 13804 8988 13860 9018
rect 14512 11786 14568 11788
rect 14512 11734 14514 11786
rect 14514 11734 14566 11786
rect 14566 11734 14568 11786
rect 14512 11732 14568 11734
rect 14616 11786 14672 11788
rect 14616 11734 14618 11786
rect 14618 11734 14670 11786
rect 14670 11734 14672 11786
rect 14616 11732 14672 11734
rect 14720 11786 14776 11788
rect 14720 11734 14722 11786
rect 14722 11734 14774 11786
rect 14774 11734 14776 11786
rect 14720 11732 14776 11734
rect 14512 10218 14568 10220
rect 14512 10166 14514 10218
rect 14514 10166 14566 10218
rect 14566 10166 14568 10218
rect 14512 10164 14568 10166
rect 14616 10218 14672 10220
rect 14616 10166 14618 10218
rect 14618 10166 14670 10218
rect 14670 10166 14672 10218
rect 14616 10164 14672 10166
rect 14720 10218 14776 10220
rect 14720 10166 14722 10218
rect 14722 10166 14774 10218
rect 14774 10166 14776 10218
rect 14720 10164 14776 10166
rect 14364 9996 14420 10052
rect 15260 14476 15316 14532
rect 17172 14138 17228 14140
rect 17172 14086 17174 14138
rect 17174 14086 17226 14138
rect 17226 14086 17228 14138
rect 17172 14084 17228 14086
rect 17276 14138 17332 14140
rect 17276 14086 17278 14138
rect 17278 14086 17330 14138
rect 17330 14086 17332 14138
rect 17276 14084 17332 14086
rect 17380 14138 17436 14140
rect 17380 14086 17382 14138
rect 17382 14086 17434 14138
rect 17434 14086 17436 14138
rect 17380 14084 17436 14086
rect 16828 13020 16884 13076
rect 15316 12572 15372 12628
rect 16380 12572 16436 12628
rect 17612 12962 17668 12964
rect 17612 12910 17614 12962
rect 17614 12910 17666 12962
rect 17666 12910 17668 12962
rect 17612 12908 17668 12910
rect 17172 12570 17228 12572
rect 17172 12518 17174 12570
rect 17174 12518 17226 12570
rect 17226 12518 17228 12570
rect 17172 12516 17228 12518
rect 17276 12570 17332 12572
rect 17276 12518 17278 12570
rect 17278 12518 17330 12570
rect 17330 12518 17332 12570
rect 17276 12516 17332 12518
rect 17380 12570 17436 12572
rect 17380 12518 17382 12570
rect 17382 12518 17434 12570
rect 17434 12518 17436 12570
rect 17380 12516 17436 12518
rect 18172 18450 18228 18452
rect 18172 18398 18174 18450
rect 18174 18398 18226 18450
rect 18226 18398 18228 18450
rect 18172 18396 18228 18398
rect 19832 19626 19888 19628
rect 19832 19574 19834 19626
rect 19834 19574 19886 19626
rect 19886 19574 19888 19626
rect 19832 19572 19888 19574
rect 19936 19626 19992 19628
rect 19936 19574 19938 19626
rect 19938 19574 19990 19626
rect 19990 19574 19992 19626
rect 19936 19572 19992 19574
rect 20040 19626 20096 19628
rect 20040 19574 20042 19626
rect 20042 19574 20094 19626
rect 20094 19574 20096 19626
rect 20040 19572 20096 19574
rect 20636 19404 20692 19460
rect 19628 19180 19684 19236
rect 19740 18956 19796 19012
rect 19068 18396 19124 18452
rect 20412 19010 20468 19012
rect 20412 18958 20414 19010
rect 20414 18958 20466 19010
rect 20466 18958 20468 19010
rect 20412 18956 20468 18958
rect 20860 18956 20916 19012
rect 19628 18450 19684 18452
rect 19628 18398 19630 18450
rect 19630 18398 19682 18450
rect 19682 18398 19684 18450
rect 19628 18396 19684 18398
rect 19852 18450 19908 18452
rect 19852 18398 19854 18450
rect 19854 18398 19906 18450
rect 19906 18398 19908 18450
rect 19852 18396 19908 18398
rect 20580 18450 20636 18452
rect 20580 18398 20582 18450
rect 20582 18398 20634 18450
rect 20634 18398 20636 18450
rect 20580 18396 20636 18398
rect 22316 19068 22372 19124
rect 21588 18450 21644 18452
rect 21588 18398 21590 18450
rect 21590 18398 21642 18450
rect 21642 18398 21644 18450
rect 21588 18396 21644 18398
rect 18956 18338 19012 18340
rect 18956 18286 18958 18338
rect 18958 18286 19010 18338
rect 19010 18286 19012 18338
rect 18956 18284 19012 18286
rect 19832 18058 19888 18060
rect 19832 18006 19834 18058
rect 19834 18006 19886 18058
rect 19886 18006 19888 18058
rect 19832 18004 19888 18006
rect 19936 18058 19992 18060
rect 19936 18006 19938 18058
rect 19938 18006 19990 18058
rect 19990 18006 19992 18058
rect 19936 18004 19992 18006
rect 20040 18058 20096 18060
rect 20040 18006 20042 18058
rect 20042 18006 20094 18058
rect 20094 18006 20096 18058
rect 20040 18004 20096 18006
rect 18620 16492 18676 16548
rect 19832 16490 19888 16492
rect 19832 16438 19834 16490
rect 19834 16438 19886 16490
rect 19886 16438 19888 16490
rect 19832 16436 19888 16438
rect 19936 16490 19992 16492
rect 19936 16438 19938 16490
rect 19938 16438 19990 16490
rect 19990 16438 19992 16490
rect 19936 16436 19992 16438
rect 20040 16490 20096 16492
rect 20040 16438 20042 16490
rect 20042 16438 20094 16490
rect 20094 16438 20096 16490
rect 20040 16436 20096 16438
rect 18060 13074 18116 13076
rect 18060 13022 18062 13074
rect 18062 13022 18114 13074
rect 18114 13022 18116 13074
rect 18060 13020 18116 13022
rect 17836 12684 17892 12740
rect 18620 15260 18676 15316
rect 18284 12460 18340 12516
rect 18508 12460 18564 12516
rect 17948 12348 18004 12404
rect 17052 11340 17108 11396
rect 17172 11002 17228 11004
rect 17172 10950 17174 11002
rect 17174 10950 17226 11002
rect 17226 10950 17228 11002
rect 17172 10948 17228 10950
rect 17276 11002 17332 11004
rect 17276 10950 17278 11002
rect 17278 10950 17330 11002
rect 17330 10950 17332 11002
rect 17276 10948 17332 10950
rect 17380 11002 17436 11004
rect 17380 10950 17382 11002
rect 17382 10950 17434 11002
rect 17434 10950 17436 11002
rect 17380 10948 17436 10950
rect 15148 9996 15204 10052
rect 17172 9434 17228 9436
rect 17172 9382 17174 9434
rect 17174 9382 17226 9434
rect 17226 9382 17228 9434
rect 17172 9380 17228 9382
rect 17276 9434 17332 9436
rect 17276 9382 17278 9434
rect 17278 9382 17330 9434
rect 17330 9382 17332 9434
rect 17276 9380 17332 9382
rect 17380 9434 17436 9436
rect 17380 9382 17382 9434
rect 17382 9382 17434 9434
rect 17434 9382 17436 9434
rect 17380 9380 17436 9382
rect 14958 9212 15014 9268
rect 17724 11340 17780 11396
rect 17948 11900 18004 11956
rect 17612 9100 17668 9156
rect 14700 9042 14756 9044
rect 14700 8990 14702 9042
rect 14702 8990 14754 9042
rect 14754 8990 14756 9042
rect 14700 8988 14756 8990
rect 14252 7980 14308 8036
rect 14812 8764 14868 8820
rect 14512 8650 14568 8652
rect 14512 8598 14514 8650
rect 14514 8598 14566 8650
rect 14566 8598 14568 8650
rect 14512 8596 14568 8598
rect 14616 8650 14672 8652
rect 14616 8598 14618 8650
rect 14618 8598 14670 8650
rect 14670 8598 14672 8650
rect 14616 8596 14672 8598
rect 14720 8650 14776 8652
rect 14720 8598 14722 8650
rect 14722 8598 14774 8650
rect 14774 8598 14776 8650
rect 14720 8596 14776 8598
rect 15372 8316 15428 8372
rect 17500 8316 17556 8372
rect 18620 11564 18676 11620
rect 18844 16098 18900 16100
rect 18844 16046 18846 16098
rect 18846 16046 18898 16098
rect 18898 16046 18900 16098
rect 18844 16044 18900 16046
rect 19068 15314 19124 15316
rect 19068 15262 19070 15314
rect 19070 15262 19122 15314
rect 19122 15262 19124 15314
rect 19068 15260 19124 15262
rect 19832 14922 19888 14924
rect 19832 14870 19834 14922
rect 19834 14870 19886 14922
rect 19886 14870 19888 14922
rect 19832 14868 19888 14870
rect 19936 14922 19992 14924
rect 19936 14870 19938 14922
rect 19938 14870 19990 14922
rect 19990 14870 19992 14922
rect 19936 14868 19992 14870
rect 20040 14922 20096 14924
rect 20040 14870 20042 14922
rect 20042 14870 20094 14922
rect 20094 14870 20096 14922
rect 20040 14868 20096 14870
rect 20300 14252 20356 14308
rect 19740 13746 19796 13748
rect 19740 13694 19742 13746
rect 19742 13694 19794 13746
rect 19794 13694 19796 13746
rect 19740 13692 19796 13694
rect 19404 13580 19460 13636
rect 19832 13354 19888 13356
rect 19832 13302 19834 13354
rect 19834 13302 19886 13354
rect 19886 13302 19888 13354
rect 19832 13300 19888 13302
rect 19936 13354 19992 13356
rect 19936 13302 19938 13354
rect 19938 13302 19990 13354
rect 19990 13302 19992 13354
rect 19936 13300 19992 13302
rect 20040 13354 20096 13356
rect 20040 13302 20042 13354
rect 20042 13302 20094 13354
rect 20094 13302 20096 13354
rect 20040 13300 20096 13302
rect 20188 13020 20244 13076
rect 22492 18842 22548 18844
rect 22492 18790 22494 18842
rect 22494 18790 22546 18842
rect 22546 18790 22548 18842
rect 22492 18788 22548 18790
rect 22596 18842 22652 18844
rect 22596 18790 22598 18842
rect 22598 18790 22650 18842
rect 22650 18790 22652 18842
rect 22596 18788 22652 18790
rect 22700 18842 22756 18844
rect 22700 18790 22702 18842
rect 22702 18790 22754 18842
rect 22754 18790 22756 18842
rect 22700 18788 22756 18790
rect 22316 18450 22372 18452
rect 22316 18398 22318 18450
rect 22318 18398 22370 18450
rect 22370 18398 22372 18450
rect 22316 18396 22372 18398
rect 21588 16994 21644 16996
rect 21588 16942 21590 16994
rect 21590 16942 21642 16994
rect 21642 16942 21644 16994
rect 21588 16940 21644 16942
rect 21196 16828 21252 16884
rect 21980 16882 22036 16884
rect 21980 16830 21982 16882
rect 21982 16830 22034 16882
rect 22034 16830 22036 16882
rect 21980 16828 22036 16830
rect 21532 14306 21588 14308
rect 21532 14254 21534 14306
rect 21534 14254 21586 14306
rect 21586 14254 21588 14306
rect 21532 14252 21588 14254
rect 21084 13634 21140 13636
rect 21084 13582 21086 13634
rect 21086 13582 21138 13634
rect 21138 13582 21140 13634
rect 21084 13580 21140 13582
rect 20804 13244 20860 13300
rect 20972 13020 21028 13076
rect 20300 12796 20356 12852
rect 18620 11394 18676 11396
rect 18620 11342 18622 11394
rect 18622 11342 18674 11394
rect 18674 11342 18676 11394
rect 18620 11340 18676 11342
rect 17836 9826 17892 9828
rect 17836 9774 17838 9826
rect 17838 9774 17890 9826
rect 17890 9774 17892 9826
rect 17836 9772 17892 9774
rect 17724 8204 17780 8260
rect 17172 7866 17228 7868
rect 17172 7814 17174 7866
rect 17174 7814 17226 7866
rect 17226 7814 17228 7866
rect 17172 7812 17228 7814
rect 17276 7866 17332 7868
rect 17276 7814 17278 7866
rect 17278 7814 17330 7866
rect 17330 7814 17332 7866
rect 17276 7812 17332 7814
rect 17380 7866 17436 7868
rect 17380 7814 17382 7866
rect 17382 7814 17434 7866
rect 17434 7814 17436 7866
rect 17380 7812 17436 7814
rect 14512 7082 14568 7084
rect 14512 7030 14514 7082
rect 14514 7030 14566 7082
rect 14566 7030 14568 7082
rect 14512 7028 14568 7030
rect 14616 7082 14672 7084
rect 14616 7030 14618 7082
rect 14618 7030 14670 7082
rect 14670 7030 14672 7082
rect 14616 7028 14672 7030
rect 14720 7082 14776 7084
rect 14720 7030 14722 7082
rect 14722 7030 14774 7082
rect 14774 7030 14776 7082
rect 14720 7028 14776 7030
rect 14588 6860 14644 6916
rect 17172 6298 17228 6300
rect 17172 6246 17174 6298
rect 17174 6246 17226 6298
rect 17226 6246 17228 6298
rect 17172 6244 17228 6246
rect 17276 6298 17332 6300
rect 17276 6246 17278 6298
rect 17278 6246 17330 6298
rect 17330 6246 17332 6298
rect 17276 6244 17332 6246
rect 17380 6298 17436 6300
rect 17380 6246 17382 6298
rect 17382 6246 17434 6298
rect 17434 6246 17436 6298
rect 17380 6244 17436 6246
rect 14476 5906 14532 5908
rect 14476 5854 14478 5906
rect 14478 5854 14530 5906
rect 14530 5854 14532 5906
rect 14476 5852 14532 5854
rect 16828 5852 16884 5908
rect 15372 5740 15428 5796
rect 14512 5514 14568 5516
rect 14512 5462 14514 5514
rect 14514 5462 14566 5514
rect 14566 5462 14568 5514
rect 14512 5460 14568 5462
rect 14616 5514 14672 5516
rect 14616 5462 14618 5514
rect 14618 5462 14670 5514
rect 14670 5462 14672 5514
rect 14616 5460 14672 5462
rect 14720 5514 14776 5516
rect 14720 5462 14722 5514
rect 14722 5462 14774 5514
rect 14774 5462 14776 5514
rect 14720 5460 14776 5462
rect 14028 5292 14084 5348
rect 13580 4956 13636 5012
rect 11852 4730 11908 4732
rect 11852 4678 11854 4730
rect 11854 4678 11906 4730
rect 11906 4678 11908 4730
rect 11852 4676 11908 4678
rect 11956 4730 12012 4732
rect 11956 4678 11958 4730
rect 11958 4678 12010 4730
rect 12010 4678 12012 4730
rect 11956 4676 12012 4678
rect 12060 4730 12116 4732
rect 12060 4678 12062 4730
rect 12062 4678 12114 4730
rect 12114 4678 12116 4730
rect 12060 4676 12116 4678
rect 12572 4844 12628 4900
rect 13804 5122 13860 5124
rect 13804 5070 13806 5122
rect 13806 5070 13858 5122
rect 13858 5070 13860 5122
rect 13804 5068 13860 5070
rect 13636 4562 13692 4564
rect 13636 4510 13638 4562
rect 13638 4510 13690 4562
rect 13690 4510 13692 4562
rect 13636 4508 13692 4510
rect 15932 5740 15988 5796
rect 15596 5628 15652 5684
rect 16828 5404 16884 5460
rect 17164 5516 17220 5572
rect 17164 5234 17220 5236
rect 17164 5182 17166 5234
rect 17166 5182 17218 5234
rect 17218 5182 17220 5234
rect 17164 5180 17220 5182
rect 17836 9548 17892 9604
rect 18508 8988 18564 9044
rect 18452 8258 18508 8260
rect 18452 8206 18454 8258
rect 18454 8206 18506 8258
rect 18506 8206 18508 8258
rect 18452 8204 18508 8206
rect 17892 7698 17948 7700
rect 17892 7646 17894 7698
rect 17894 7646 17946 7698
rect 17946 7646 17948 7698
rect 17892 7644 17948 7646
rect 18340 8092 18396 8148
rect 19068 12460 19124 12516
rect 19516 12348 19572 12404
rect 18844 12012 18900 12068
rect 20300 12066 20356 12068
rect 20300 12014 20302 12066
rect 20302 12014 20354 12066
rect 20354 12014 20356 12066
rect 20300 12012 20356 12014
rect 19832 11786 19888 11788
rect 19832 11734 19834 11786
rect 19834 11734 19886 11786
rect 19886 11734 19888 11786
rect 19832 11732 19888 11734
rect 19936 11786 19992 11788
rect 19936 11734 19938 11786
rect 19938 11734 19990 11786
rect 19990 11734 19992 11786
rect 19936 11732 19992 11734
rect 20040 11786 20096 11788
rect 20040 11734 20042 11786
rect 20042 11734 20094 11786
rect 20094 11734 20096 11786
rect 20040 11732 20096 11734
rect 19124 11618 19180 11620
rect 19124 11566 19126 11618
rect 19126 11566 19178 11618
rect 19178 11566 19180 11618
rect 19124 11564 19180 11566
rect 19832 10218 19888 10220
rect 19832 10166 19834 10218
rect 19834 10166 19886 10218
rect 19886 10166 19888 10218
rect 19832 10164 19888 10166
rect 19936 10218 19992 10220
rect 19936 10166 19938 10218
rect 19938 10166 19990 10218
rect 19990 10166 19992 10218
rect 19936 10164 19992 10166
rect 20040 10218 20096 10220
rect 20040 10166 20042 10218
rect 20042 10166 20094 10218
rect 20094 10166 20096 10218
rect 20040 10164 20096 10166
rect 20412 9996 20468 10052
rect 19068 9826 19124 9828
rect 19068 9774 19070 9826
rect 19070 9774 19122 9826
rect 19122 9774 19124 9826
rect 19068 9772 19124 9774
rect 19292 9772 19348 9828
rect 18900 9602 18956 9604
rect 18900 9550 18902 9602
rect 18902 9550 18954 9602
rect 18954 9550 18956 9602
rect 18900 9548 18956 9550
rect 20188 9772 20244 9828
rect 19460 9714 19516 9716
rect 19460 9662 19462 9714
rect 19462 9662 19514 9714
rect 19514 9662 19516 9714
rect 19460 9660 19516 9662
rect 18956 9042 19012 9044
rect 18956 8990 18958 9042
rect 18958 8990 19010 9042
rect 19010 8990 19012 9042
rect 18956 8988 19012 8990
rect 19124 8876 19180 8932
rect 19124 8428 19180 8484
rect 18844 8092 18900 8148
rect 19684 9042 19740 9044
rect 19684 8990 19686 9042
rect 19686 8990 19738 9042
rect 19738 8990 19740 9042
rect 19684 8988 19740 8990
rect 19832 8650 19888 8652
rect 19832 8598 19834 8650
rect 19834 8598 19886 8650
rect 19886 8598 19888 8650
rect 19832 8596 19888 8598
rect 19936 8650 19992 8652
rect 19936 8598 19938 8650
rect 19938 8598 19990 8650
rect 19990 8598 19992 8650
rect 19936 8596 19992 8598
rect 20040 8650 20096 8652
rect 20040 8598 20042 8650
rect 20042 8598 20094 8650
rect 20094 8598 20096 8650
rect 20040 8596 20096 8598
rect 19292 8092 19348 8148
rect 20300 9042 20356 9044
rect 20300 8990 20302 9042
rect 20302 8990 20354 9042
rect 20354 8990 20356 9042
rect 20300 8988 20356 8990
rect 20524 9826 20580 9828
rect 20524 9774 20526 9826
rect 20526 9774 20578 9826
rect 20578 9774 20580 9826
rect 20524 9772 20580 9774
rect 20748 9548 20804 9604
rect 20636 9266 20692 9268
rect 20636 9214 20638 9266
rect 20638 9214 20690 9266
rect 20690 9214 20692 9266
rect 20636 9212 20692 9214
rect 20636 8876 20692 8932
rect 20636 8428 20692 8484
rect 19068 7644 19124 7700
rect 19516 7308 19572 7364
rect 18508 5516 18564 5572
rect 17724 4844 17780 4900
rect 17836 5180 17892 5236
rect 18060 5107 18116 5124
rect 18060 5068 18062 5107
rect 18062 5068 18114 5107
rect 18114 5068 18116 5107
rect 18620 5292 18676 5348
rect 20412 7362 20468 7364
rect 20412 7310 20414 7362
rect 20414 7310 20466 7362
rect 20466 7310 20468 7362
rect 20412 7308 20468 7310
rect 19832 7082 19888 7084
rect 19832 7030 19834 7082
rect 19834 7030 19886 7082
rect 19886 7030 19888 7082
rect 19832 7028 19888 7030
rect 19936 7082 19992 7084
rect 19936 7030 19938 7082
rect 19938 7030 19990 7082
rect 19990 7030 19992 7082
rect 19936 7028 19992 7030
rect 20040 7082 20096 7084
rect 20040 7030 20042 7082
rect 20042 7030 20094 7082
rect 20094 7030 20096 7082
rect 20040 7028 20096 7030
rect 20076 5906 20132 5908
rect 20076 5854 20078 5906
rect 20078 5854 20130 5906
rect 20130 5854 20132 5906
rect 20076 5852 20132 5854
rect 20300 5852 20356 5908
rect 19404 5292 19460 5348
rect 19292 5180 19348 5236
rect 20300 5628 20356 5684
rect 19832 5514 19888 5516
rect 19832 5462 19834 5514
rect 19834 5462 19886 5514
rect 19886 5462 19888 5514
rect 19832 5460 19888 5462
rect 19936 5514 19992 5516
rect 19936 5462 19938 5514
rect 19938 5462 19990 5514
rect 19990 5462 19992 5514
rect 19936 5460 19992 5462
rect 20040 5514 20096 5516
rect 20040 5462 20042 5514
rect 20042 5462 20094 5514
rect 20094 5462 20096 5514
rect 20040 5460 20096 5462
rect 18844 5122 18900 5124
rect 18844 5070 18846 5122
rect 18846 5070 18898 5122
rect 18898 5070 18900 5122
rect 18844 5068 18900 5070
rect 17172 4730 17228 4732
rect 17172 4678 17174 4730
rect 17174 4678 17226 4730
rect 17226 4678 17228 4730
rect 17172 4676 17228 4678
rect 17276 4730 17332 4732
rect 17276 4678 17278 4730
rect 17278 4678 17330 4730
rect 17330 4678 17332 4730
rect 17276 4676 17332 4678
rect 17380 4730 17436 4732
rect 17380 4678 17382 4730
rect 17382 4678 17434 4730
rect 17434 4678 17436 4730
rect 17380 4676 17436 4678
rect 15260 4508 15316 4564
rect 17444 4562 17500 4564
rect 17444 4510 17446 4562
rect 17446 4510 17498 4562
rect 17498 4510 17500 4562
rect 17444 4508 17500 4510
rect 19740 4956 19796 5012
rect 20020 4956 20076 5012
rect 20524 4338 20580 4340
rect 20524 4286 20526 4338
rect 20526 4286 20578 4338
rect 20578 4286 20580 4338
rect 20524 4284 20580 4286
rect 21644 13132 21700 13188
rect 21476 13074 21532 13076
rect 21476 13022 21478 13074
rect 21478 13022 21530 13074
rect 21530 13022 21532 13074
rect 21476 13020 21532 13022
rect 21588 10332 21644 10388
rect 21980 13186 22036 13188
rect 21980 13134 21982 13186
rect 21982 13134 22034 13186
rect 22034 13134 22036 13186
rect 21980 13132 22036 13134
rect 21756 9996 21812 10052
rect 21812 9826 21868 9828
rect 21812 9774 21814 9826
rect 21814 9774 21866 9826
rect 21866 9774 21868 9826
rect 21812 9772 21868 9774
rect 20860 9212 20916 9268
rect 22092 8876 22148 8932
rect 21980 8258 22036 8260
rect 21980 8206 21982 8258
rect 21982 8206 22034 8258
rect 22034 8206 22036 8258
rect 21980 8204 22036 8206
rect 21588 8146 21644 8148
rect 21588 8094 21590 8146
rect 21590 8094 21642 8146
rect 21642 8094 21644 8146
rect 21588 8092 21644 8094
rect 20972 7980 21028 8036
rect 22492 17274 22548 17276
rect 22492 17222 22494 17274
rect 22494 17222 22546 17274
rect 22546 17222 22548 17274
rect 22492 17220 22548 17222
rect 22596 17274 22652 17276
rect 22596 17222 22598 17274
rect 22598 17222 22650 17274
rect 22650 17222 22652 17274
rect 22596 17220 22652 17222
rect 22700 17274 22756 17276
rect 22700 17222 22702 17274
rect 22702 17222 22754 17274
rect 22754 17222 22756 17274
rect 22700 17220 22756 17222
rect 22316 16940 22372 16996
rect 22316 16156 22372 16212
rect 22492 15706 22548 15708
rect 22492 15654 22494 15706
rect 22494 15654 22546 15706
rect 22546 15654 22548 15706
rect 22492 15652 22548 15654
rect 22596 15706 22652 15708
rect 22596 15654 22598 15706
rect 22598 15654 22650 15706
rect 22650 15654 22652 15706
rect 22596 15652 22652 15654
rect 22700 15706 22756 15708
rect 22700 15654 22702 15706
rect 22702 15654 22754 15706
rect 22754 15654 22756 15706
rect 22700 15652 22756 15654
rect 22492 14138 22548 14140
rect 22492 14086 22494 14138
rect 22494 14086 22546 14138
rect 22546 14086 22548 14138
rect 22492 14084 22548 14086
rect 22596 14138 22652 14140
rect 22596 14086 22598 14138
rect 22598 14086 22650 14138
rect 22650 14086 22652 14138
rect 22596 14084 22652 14086
rect 22700 14138 22756 14140
rect 22700 14086 22702 14138
rect 22702 14086 22754 14138
rect 22754 14086 22756 14138
rect 22700 14084 22756 14086
rect 22316 13244 22372 13300
rect 22492 12570 22548 12572
rect 22492 12518 22494 12570
rect 22494 12518 22546 12570
rect 22546 12518 22548 12570
rect 22492 12516 22548 12518
rect 22596 12570 22652 12572
rect 22596 12518 22598 12570
rect 22598 12518 22650 12570
rect 22650 12518 22652 12570
rect 22596 12516 22652 12518
rect 22700 12570 22756 12572
rect 22700 12518 22702 12570
rect 22702 12518 22754 12570
rect 22754 12518 22756 12570
rect 22700 12516 22756 12518
rect 22492 11002 22548 11004
rect 22492 10950 22494 11002
rect 22494 10950 22546 11002
rect 22546 10950 22548 11002
rect 22492 10948 22548 10950
rect 22596 11002 22652 11004
rect 22596 10950 22598 11002
rect 22598 10950 22650 11002
rect 22650 10950 22652 11002
rect 22596 10948 22652 10950
rect 22700 11002 22756 11004
rect 22700 10950 22702 11002
rect 22702 10950 22754 11002
rect 22754 10950 22756 11002
rect 22700 10948 22756 10950
rect 22316 10332 22372 10388
rect 22492 9434 22548 9436
rect 22492 9382 22494 9434
rect 22494 9382 22546 9434
rect 22546 9382 22548 9434
rect 22492 9380 22548 9382
rect 22596 9434 22652 9436
rect 22596 9382 22598 9434
rect 22598 9382 22650 9434
rect 22650 9382 22652 9434
rect 22596 9380 22652 9382
rect 22700 9434 22756 9436
rect 22700 9382 22702 9434
rect 22702 9382 22754 9434
rect 22754 9382 22756 9434
rect 22700 9380 22756 9382
rect 22204 7980 22260 8036
rect 22316 8092 22372 8148
rect 22492 7866 22548 7868
rect 22492 7814 22494 7866
rect 22494 7814 22546 7866
rect 22546 7814 22548 7866
rect 22492 7812 22548 7814
rect 22596 7866 22652 7868
rect 22596 7814 22598 7866
rect 22598 7814 22650 7866
rect 22650 7814 22652 7866
rect 22596 7812 22652 7814
rect 22700 7866 22756 7868
rect 22700 7814 22702 7866
rect 22702 7814 22754 7866
rect 22754 7814 22756 7866
rect 22700 7812 22756 7814
rect 22316 7420 22372 7476
rect 22492 6298 22548 6300
rect 22492 6246 22494 6298
rect 22494 6246 22546 6298
rect 22546 6246 22548 6298
rect 22492 6244 22548 6246
rect 22596 6298 22652 6300
rect 22596 6246 22598 6298
rect 22598 6246 22650 6298
rect 22650 6246 22652 6298
rect 22596 6244 22652 6246
rect 22700 6298 22756 6300
rect 22700 6246 22702 6298
rect 22702 6246 22754 6298
rect 22754 6246 22756 6298
rect 22700 6244 22756 6246
rect 20860 5740 20916 5796
rect 20860 5180 20916 5236
rect 21980 5234 22036 5236
rect 21980 5182 21982 5234
rect 21982 5182 22034 5234
rect 22034 5182 22036 5234
rect 21980 5180 22036 5182
rect 21588 5122 21644 5124
rect 21588 5070 21590 5122
rect 21590 5070 21642 5122
rect 21642 5070 21644 5122
rect 21588 5068 21644 5070
rect 22316 5122 22372 5124
rect 22316 5070 22318 5122
rect 22318 5070 22370 5122
rect 22370 5070 22372 5122
rect 22316 5068 22372 5070
rect 22492 4730 22548 4732
rect 22492 4678 22494 4730
rect 22494 4678 22546 4730
rect 22546 4678 22548 4730
rect 22492 4676 22548 4678
rect 22596 4730 22652 4732
rect 22596 4678 22598 4730
rect 22598 4678 22650 4730
rect 22650 4678 22652 4730
rect 22596 4676 22652 4678
rect 22700 4730 22756 4732
rect 22700 4678 22702 4730
rect 22702 4678 22754 4730
rect 22754 4678 22756 4730
rect 22700 4676 22756 4678
rect 22316 4508 22372 4564
rect 21196 4338 21252 4340
rect 21196 4286 21198 4338
rect 21198 4286 21250 4338
rect 21250 4286 21252 4338
rect 21196 4284 21252 4286
rect 21700 4284 21756 4340
rect 3872 3946 3928 3948
rect 3872 3894 3874 3946
rect 3874 3894 3926 3946
rect 3926 3894 3928 3946
rect 3872 3892 3928 3894
rect 3976 3946 4032 3948
rect 3976 3894 3978 3946
rect 3978 3894 4030 3946
rect 4030 3894 4032 3946
rect 3976 3892 4032 3894
rect 4080 3946 4136 3948
rect 4080 3894 4082 3946
rect 4082 3894 4134 3946
rect 4134 3894 4136 3946
rect 4080 3892 4136 3894
rect 9192 3946 9248 3948
rect 9192 3894 9194 3946
rect 9194 3894 9246 3946
rect 9246 3894 9248 3946
rect 9192 3892 9248 3894
rect 9296 3946 9352 3948
rect 9296 3894 9298 3946
rect 9298 3894 9350 3946
rect 9350 3894 9352 3946
rect 9296 3892 9352 3894
rect 9400 3946 9456 3948
rect 9400 3894 9402 3946
rect 9402 3894 9454 3946
rect 9454 3894 9456 3946
rect 9400 3892 9456 3894
rect 14512 3946 14568 3948
rect 14512 3894 14514 3946
rect 14514 3894 14566 3946
rect 14566 3894 14568 3946
rect 14512 3892 14568 3894
rect 14616 3946 14672 3948
rect 14616 3894 14618 3946
rect 14618 3894 14670 3946
rect 14670 3894 14672 3946
rect 14616 3892 14672 3894
rect 14720 3946 14776 3948
rect 14720 3894 14722 3946
rect 14722 3894 14774 3946
rect 14774 3894 14776 3946
rect 14720 3892 14776 3894
rect 19832 3946 19888 3948
rect 19832 3894 19834 3946
rect 19834 3894 19886 3946
rect 19886 3894 19888 3946
rect 19832 3892 19888 3894
rect 19936 3946 19992 3948
rect 19936 3894 19938 3946
rect 19938 3894 19990 3946
rect 19990 3894 19992 3946
rect 19936 3892 19992 3894
rect 20040 3946 20096 3948
rect 20040 3894 20042 3946
rect 20042 3894 20094 3946
rect 20094 3894 20096 3946
rect 20040 3892 20096 3894
rect 6532 3162 6588 3164
rect 6532 3110 6534 3162
rect 6534 3110 6586 3162
rect 6586 3110 6588 3162
rect 6532 3108 6588 3110
rect 6636 3162 6692 3164
rect 6636 3110 6638 3162
rect 6638 3110 6690 3162
rect 6690 3110 6692 3162
rect 6636 3108 6692 3110
rect 6740 3162 6796 3164
rect 6740 3110 6742 3162
rect 6742 3110 6794 3162
rect 6794 3110 6796 3162
rect 6740 3108 6796 3110
rect 11852 3162 11908 3164
rect 11852 3110 11854 3162
rect 11854 3110 11906 3162
rect 11906 3110 11908 3162
rect 11852 3108 11908 3110
rect 11956 3162 12012 3164
rect 11956 3110 11958 3162
rect 11958 3110 12010 3162
rect 12010 3110 12012 3162
rect 11956 3108 12012 3110
rect 12060 3162 12116 3164
rect 12060 3110 12062 3162
rect 12062 3110 12114 3162
rect 12114 3110 12116 3162
rect 12060 3108 12116 3110
rect 17172 3162 17228 3164
rect 17172 3110 17174 3162
rect 17174 3110 17226 3162
rect 17226 3110 17228 3162
rect 17172 3108 17228 3110
rect 17276 3162 17332 3164
rect 17276 3110 17278 3162
rect 17278 3110 17330 3162
rect 17330 3110 17332 3162
rect 17276 3108 17332 3110
rect 17380 3162 17436 3164
rect 17380 3110 17382 3162
rect 17382 3110 17434 3162
rect 17434 3110 17436 3162
rect 17380 3108 17436 3110
rect 22492 3162 22548 3164
rect 22492 3110 22494 3162
rect 22494 3110 22546 3162
rect 22546 3110 22548 3162
rect 22492 3108 22548 3110
rect 22596 3162 22652 3164
rect 22596 3110 22598 3162
rect 22598 3110 22650 3162
rect 22650 3110 22652 3162
rect 22596 3108 22652 3110
rect 22700 3162 22756 3164
rect 22700 3110 22702 3162
rect 22702 3110 22754 3162
rect 22754 3110 22756 3162
rect 22700 3108 22756 3110
rect 21756 1596 21812 1652
<< metal3 >>
rect 23200 22036 24000 22064
rect 20066 21980 20076 22036
rect 20132 21980 24000 22036
rect 23200 21952 24000 21980
rect 6522 20356 6532 20412
rect 6588 20356 6636 20412
rect 6692 20356 6740 20412
rect 6796 20356 6806 20412
rect 11842 20356 11852 20412
rect 11908 20356 11956 20412
rect 12012 20356 12060 20412
rect 12116 20356 12126 20412
rect 17162 20356 17172 20412
rect 17228 20356 17276 20412
rect 17332 20356 17380 20412
rect 17436 20356 17446 20412
rect 22482 20356 22492 20412
rect 22548 20356 22596 20412
rect 22652 20356 22700 20412
rect 22756 20356 22766 20412
rect 19842 20076 19852 20132
rect 19908 20076 20972 20132
rect 21028 20076 21038 20132
rect 5842 19964 5852 20020
rect 5908 19964 9212 20020
rect 9268 19964 9278 20020
rect 3862 19572 3872 19628
rect 3928 19572 3976 19628
rect 4032 19572 4080 19628
rect 4136 19572 4146 19628
rect 9182 19572 9192 19628
rect 9248 19572 9296 19628
rect 9352 19572 9400 19628
rect 9456 19572 9466 19628
rect 14502 19572 14512 19628
rect 14568 19572 14616 19628
rect 14672 19572 14720 19628
rect 14776 19572 14786 19628
rect 19822 19572 19832 19628
rect 19888 19572 19936 19628
rect 19992 19572 20040 19628
rect 20096 19572 20106 19628
rect 4498 19404 4508 19460
rect 4564 19404 6412 19460
rect 6468 19404 6478 19460
rect 16370 19404 16380 19460
rect 16436 19404 17612 19460
rect 17668 19404 17678 19460
rect 18610 19404 18620 19460
rect 18676 19404 20636 19460
rect 20692 19404 20702 19460
rect 4050 19180 4060 19236
rect 4116 19180 5012 19236
rect 5068 19180 5078 19236
rect 5170 19180 5180 19236
rect 5236 19180 14252 19236
rect 14308 19180 19628 19236
rect 19684 19180 19694 19236
rect 23200 19124 24000 19152
rect 22306 19068 22316 19124
rect 22372 19068 24000 19124
rect 23200 19040 24000 19068
rect 14130 18956 14140 19012
rect 14196 18956 14924 19012
rect 14980 18956 15764 19012
rect 15820 18956 15830 19012
rect 19730 18956 19740 19012
rect 19796 18956 20412 19012
rect 20468 18956 20860 19012
rect 20916 18956 20926 19012
rect 6522 18788 6532 18844
rect 6588 18788 6636 18844
rect 6692 18788 6740 18844
rect 6796 18788 6806 18844
rect 11842 18788 11852 18844
rect 11908 18788 11956 18844
rect 12012 18788 12060 18844
rect 12116 18788 12126 18844
rect 17162 18788 17172 18844
rect 17228 18788 17276 18844
rect 17332 18788 17380 18844
rect 17436 18788 17446 18844
rect 22482 18788 22492 18844
rect 22548 18788 22596 18844
rect 22652 18788 22700 18844
rect 22756 18788 22766 18844
rect 3378 18508 3388 18564
rect 3444 18508 4508 18564
rect 4564 18508 5516 18564
rect 5572 18508 5582 18564
rect 7634 18508 7644 18564
rect 7700 18508 8652 18564
rect 8708 18508 8718 18564
rect 9426 18508 9436 18564
rect 9492 18508 9502 18564
rect 9436 18452 9492 18508
rect 9436 18396 9996 18452
rect 10052 18396 14028 18452
rect 14084 18396 16044 18452
rect 16100 18396 16110 18452
rect 18162 18396 18172 18452
rect 18228 18396 19068 18452
rect 19124 18396 19628 18452
rect 19684 18396 19694 18452
rect 19842 18396 19852 18452
rect 19908 18396 20580 18452
rect 20636 18396 20646 18452
rect 21578 18396 21588 18452
rect 21644 18396 22316 18452
rect 22372 18396 22382 18452
rect 7746 18284 7756 18340
rect 7812 18284 9660 18340
rect 9716 18284 9726 18340
rect 13682 18284 13692 18340
rect 13748 18284 18956 18340
rect 19012 18284 19022 18340
rect 13850 18172 13860 18228
rect 13916 18172 14700 18228
rect 14756 18172 14766 18228
rect 3862 18004 3872 18060
rect 3928 18004 3976 18060
rect 4032 18004 4080 18060
rect 4136 18004 4146 18060
rect 9182 18004 9192 18060
rect 9248 18004 9296 18060
rect 9352 18004 9400 18060
rect 9456 18004 9466 18060
rect 14502 18004 14512 18060
rect 14568 18004 14616 18060
rect 14672 18004 14720 18060
rect 14776 18004 14786 18060
rect 19822 18004 19832 18060
rect 19888 18004 19936 18060
rect 19992 18004 20040 18060
rect 20096 18004 20106 18060
rect 3546 17948 3556 18004
rect 3612 17892 3668 18004
rect 3612 17836 4564 17892
rect 3490 17724 3500 17780
rect 3556 17724 3948 17780
rect 4004 17724 4014 17780
rect 4508 17556 4564 17836
rect 4834 17612 4844 17668
rect 4900 17612 8876 17668
rect 8932 17612 8942 17668
rect 12674 17612 12684 17668
rect 12740 17612 13580 17668
rect 13636 17612 14364 17668
rect 14420 17612 14430 17668
rect 4498 17500 4508 17556
rect 4564 17500 4574 17556
rect 8474 17388 8484 17444
rect 8540 17388 14924 17444
rect 14980 17388 14990 17444
rect 6522 17220 6532 17276
rect 6588 17220 6636 17276
rect 6692 17220 6740 17276
rect 6796 17220 6806 17276
rect 11842 17220 11852 17276
rect 11908 17220 11956 17276
rect 12012 17220 12060 17276
rect 12116 17220 12126 17276
rect 17162 17220 17172 17276
rect 17228 17220 17276 17276
rect 17332 17220 17380 17276
rect 17436 17220 17446 17276
rect 22482 17220 22492 17276
rect 22548 17220 22596 17276
rect 22652 17220 22700 17276
rect 22756 17220 22766 17276
rect 4498 17052 4508 17108
rect 4564 17052 11676 17108
rect 11732 17052 12236 17108
rect 12292 17052 12302 17108
rect 7970 16940 7980 16996
rect 8036 16940 8484 16996
rect 8540 16940 8550 16996
rect 8866 16940 8876 16996
rect 8932 16940 13132 16996
rect 13188 16940 13198 16996
rect 21578 16940 21588 16996
rect 21644 16940 22316 16996
rect 22372 16940 22382 16996
rect 3714 16828 3724 16884
rect 3780 16828 4844 16884
rect 4900 16828 4910 16884
rect 11330 16828 11340 16884
rect 11396 16828 12012 16884
rect 12068 16828 12796 16884
rect 12852 16828 12862 16884
rect 21186 16828 21196 16884
rect 21252 16828 21980 16884
rect 22036 16828 22046 16884
rect 18610 16492 18620 16548
rect 18676 16492 18686 16548
rect 3862 16436 3872 16492
rect 3928 16436 3976 16492
rect 4032 16436 4080 16492
rect 4136 16436 4146 16492
rect 9182 16436 9192 16492
rect 9248 16436 9296 16492
rect 9352 16436 9400 16492
rect 9456 16436 9466 16492
rect 14502 16436 14512 16492
rect 14568 16436 14616 16492
rect 14672 16436 14720 16492
rect 14776 16436 14786 16492
rect 18620 16100 18676 16492
rect 19822 16436 19832 16492
rect 19888 16436 19936 16492
rect 19992 16436 20040 16492
rect 20096 16436 20106 16492
rect 23200 16212 24000 16240
rect 22306 16156 22316 16212
rect 22372 16156 24000 16212
rect 23200 16128 24000 16156
rect 3602 16044 3612 16100
rect 3668 16044 4396 16100
rect 4452 16044 4462 16100
rect 4722 16044 4732 16100
rect 4788 16044 7532 16100
rect 7588 16044 8092 16100
rect 8148 16044 14252 16100
rect 14308 16044 14318 16100
rect 14914 16044 14924 16100
rect 14980 16044 18844 16100
rect 18900 16044 18910 16100
rect 6522 15652 6532 15708
rect 6588 15652 6636 15708
rect 6692 15652 6740 15708
rect 6796 15652 6806 15708
rect 11842 15652 11852 15708
rect 11908 15652 11956 15708
rect 12012 15652 12060 15708
rect 12116 15652 12126 15708
rect 17162 15652 17172 15708
rect 17228 15652 17276 15708
rect 17332 15652 17380 15708
rect 17436 15652 17446 15708
rect 22482 15652 22492 15708
rect 22548 15652 22596 15708
rect 22652 15652 22700 15708
rect 22756 15652 22766 15708
rect 2818 15372 2828 15428
rect 2884 15372 3836 15428
rect 3892 15372 3902 15428
rect 3938 15260 3948 15316
rect 4004 15260 4676 15316
rect 4732 15260 4742 15316
rect 14914 15260 14924 15316
rect 14980 15260 18620 15316
rect 18676 15260 19068 15316
rect 19124 15260 19134 15316
rect 13906 15036 13916 15092
rect 13972 15036 14812 15092
rect 14868 15036 14878 15092
rect 3862 14868 3872 14924
rect 3928 14868 3976 14924
rect 4032 14868 4080 14924
rect 4136 14868 4146 14924
rect 9182 14868 9192 14924
rect 9248 14868 9296 14924
rect 9352 14868 9400 14924
rect 9456 14868 9466 14924
rect 14502 14868 14512 14924
rect 14568 14868 14616 14924
rect 14672 14868 14720 14924
rect 14776 14868 14786 14924
rect 19822 14868 19832 14924
rect 19888 14868 19936 14924
rect 19992 14868 20040 14924
rect 20096 14868 20106 14924
rect 5170 14588 5180 14644
rect 5236 14588 5796 14644
rect 5852 14588 7980 14644
rect 8036 14588 8046 14644
rect 12562 14476 12572 14532
rect 12628 14476 13804 14532
rect 13860 14476 15260 14532
rect 15316 14476 15326 14532
rect 4610 14252 4620 14308
rect 4676 14252 5684 14308
rect 5740 14252 13356 14308
rect 13412 14252 13422 14308
rect 20290 14252 20300 14308
rect 20356 14252 21532 14308
rect 21588 14252 21598 14308
rect 6522 14084 6532 14140
rect 6588 14084 6636 14140
rect 6692 14084 6740 14140
rect 6796 14084 6806 14140
rect 11842 14084 11852 14140
rect 11908 14084 11956 14140
rect 12012 14084 12060 14140
rect 12116 14084 12126 14140
rect 17162 14084 17172 14140
rect 17228 14084 17276 14140
rect 17332 14084 17380 14140
rect 17436 14084 17446 14140
rect 22482 14084 22492 14140
rect 22548 14084 22596 14140
rect 22652 14084 22700 14140
rect 22756 14084 22766 14140
rect 11106 13916 11116 13972
rect 11172 13916 11788 13972
rect 11844 13916 11854 13972
rect 12002 13916 12012 13972
rect 12068 13916 12572 13972
rect 12628 13916 12638 13972
rect 4162 13804 4172 13860
rect 4228 13804 7196 13860
rect 7252 13804 8092 13860
rect 8148 13804 8158 13860
rect 4834 13692 4844 13748
rect 4900 13692 7308 13748
rect 7364 13692 7374 13748
rect 8754 13692 8764 13748
rect 8820 13692 14252 13748
rect 14308 13692 19740 13748
rect 19796 13692 19806 13748
rect 19394 13580 19404 13636
rect 19460 13580 21084 13636
rect 21140 13580 21150 13636
rect 7410 13468 7420 13524
rect 7476 13468 9996 13524
rect 10052 13468 13524 13524
rect 13580 13468 14140 13524
rect 14196 13468 14206 13524
rect 3862 13300 3872 13356
rect 3928 13300 3976 13356
rect 4032 13300 4080 13356
rect 4136 13300 4146 13356
rect 9182 13300 9192 13356
rect 9248 13300 9296 13356
rect 9352 13300 9400 13356
rect 9456 13300 9466 13356
rect 14502 13300 14512 13356
rect 14568 13300 14616 13356
rect 14672 13300 14720 13356
rect 14776 13300 14786 13356
rect 19822 13300 19832 13356
rect 19888 13300 19936 13356
rect 19992 13300 20040 13356
rect 20096 13300 20106 13356
rect 23200 13300 24000 13328
rect 12226 13244 12236 13300
rect 12292 13244 12796 13300
rect 12852 13244 13860 13300
rect 20794 13244 20804 13300
rect 20860 13244 22316 13300
rect 22372 13244 24000 13300
rect 13804 13188 13860 13244
rect 23200 13216 24000 13244
rect 7858 13132 7868 13188
rect 7924 13132 8316 13188
rect 8372 13132 12124 13188
rect 12180 13132 12190 13188
rect 13794 13132 13804 13188
rect 13860 13132 14588 13188
rect 14644 13132 14654 13188
rect 21634 13132 21644 13188
rect 21700 13132 21980 13188
rect 22036 13132 22046 13188
rect 4274 13020 4284 13076
rect 4340 13020 4508 13076
rect 4564 13020 10332 13076
rect 10388 13020 10398 13076
rect 11666 13020 11676 13076
rect 11732 13020 12348 13076
rect 12404 13020 12414 13076
rect 14018 13020 14028 13076
rect 14084 13020 16828 13076
rect 16884 13020 18060 13076
rect 18116 13020 18126 13076
rect 20178 13020 20188 13076
rect 20244 13020 20972 13076
rect 21028 13020 21476 13076
rect 21532 13020 21542 13076
rect 12226 12908 12236 12964
rect 12292 12908 14364 12964
rect 14420 12908 14430 12964
rect 14578 12908 14588 12964
rect 14644 12908 17612 12964
rect 17668 12908 17678 12964
rect 14364 12852 14420 12908
rect 9874 12796 9884 12852
rect 9940 12796 13524 12852
rect 13580 12796 13590 12852
rect 14364 12796 20300 12852
rect 20356 12796 20366 12852
rect 8866 12684 8876 12740
rect 8932 12684 9772 12740
rect 9828 12684 12292 12740
rect 14018 12684 14028 12740
rect 14084 12684 17836 12740
rect 17892 12684 17902 12740
rect 12236 12628 12292 12684
rect 12236 12572 14476 12628
rect 14532 12572 14542 12628
rect 15092 12572 15316 12628
rect 15372 12572 16380 12628
rect 16436 12572 16446 12628
rect 6522 12516 6532 12572
rect 6588 12516 6636 12572
rect 6692 12516 6740 12572
rect 6796 12516 6806 12572
rect 11842 12516 11852 12572
rect 11908 12516 11956 12572
rect 12012 12516 12060 12572
rect 12116 12516 12126 12572
rect 8418 12348 8428 12404
rect 8484 12348 8876 12404
rect 8932 12348 10332 12404
rect 10388 12348 11564 12404
rect 11620 12348 13244 12404
rect 13300 12348 13310 12404
rect 15092 12292 15148 12572
rect 17162 12516 17172 12572
rect 17228 12516 17276 12572
rect 17332 12516 17380 12572
rect 17436 12516 17446 12572
rect 22482 12516 22492 12572
rect 22548 12516 22596 12572
rect 22652 12516 22700 12572
rect 22756 12516 22766 12572
rect 18274 12460 18284 12516
rect 18340 12460 18508 12516
rect 18564 12460 19068 12516
rect 19124 12460 19134 12516
rect 17938 12348 17948 12404
rect 18004 12348 19516 12404
rect 19572 12348 19582 12404
rect 8754 12236 8764 12292
rect 8820 12236 10164 12292
rect 10322 12236 10332 12292
rect 10388 12236 15148 12292
rect 7522 12124 7532 12180
rect 7588 12124 8652 12180
rect 8708 12124 9884 12180
rect 9940 12124 9950 12180
rect 10108 12124 10164 12236
rect 10220 12124 12236 12180
rect 12292 12124 13692 12180
rect 13748 12124 13758 12180
rect 18834 12012 18844 12068
rect 18900 12012 20300 12068
rect 20356 12012 20366 12068
rect 14690 11900 14700 11956
rect 14756 11900 17948 11956
rect 18004 11900 18014 11956
rect 3862 11732 3872 11788
rect 3928 11732 3976 11788
rect 4032 11732 4080 11788
rect 4136 11732 4146 11788
rect 9182 11732 9192 11788
rect 9248 11732 9296 11788
rect 9352 11732 9400 11788
rect 9456 11732 9466 11788
rect 14502 11732 14512 11788
rect 14568 11732 14616 11788
rect 14672 11732 14720 11788
rect 14776 11732 14786 11788
rect 19822 11732 19832 11788
rect 19888 11732 19936 11788
rect 19992 11732 20040 11788
rect 20096 11732 20106 11788
rect 18610 11564 18620 11620
rect 18676 11564 19124 11620
rect 19180 11564 19190 11620
rect 3154 11340 3164 11396
rect 3220 11340 3948 11396
rect 4004 11340 4508 11396
rect 4564 11340 4574 11396
rect 17042 11340 17052 11396
rect 17108 11340 17724 11396
rect 17780 11340 18620 11396
rect 18676 11340 18686 11396
rect 6522 10948 6532 11004
rect 6588 10948 6636 11004
rect 6692 10948 6740 11004
rect 6796 10948 6806 11004
rect 11842 10948 11852 11004
rect 11908 10948 11956 11004
rect 12012 10948 12060 11004
rect 12116 10948 12126 11004
rect 17162 10948 17172 11004
rect 17228 10948 17276 11004
rect 17332 10948 17380 11004
rect 17436 10948 17446 11004
rect 22482 10948 22492 11004
rect 22548 10948 22596 11004
rect 22652 10948 22700 11004
rect 22756 10948 22766 11004
rect 23200 10388 24000 10416
rect 21578 10332 21588 10388
rect 21644 10332 22316 10388
rect 22372 10332 24000 10388
rect 23200 10304 24000 10332
rect 3862 10164 3872 10220
rect 3928 10164 3976 10220
rect 4032 10164 4080 10220
rect 4136 10164 4146 10220
rect 9182 10164 9192 10220
rect 9248 10164 9296 10220
rect 9352 10164 9400 10220
rect 9456 10164 9466 10220
rect 14502 10164 14512 10220
rect 14568 10164 14616 10220
rect 14672 10164 14720 10220
rect 14776 10164 14786 10220
rect 19822 10164 19832 10220
rect 19888 10164 19936 10220
rect 19992 10164 20040 10220
rect 20096 10164 20106 10220
rect 14354 9996 14364 10052
rect 14420 9996 15148 10052
rect 15204 9996 20412 10052
rect 20468 9996 21756 10052
rect 21812 9996 21822 10052
rect 3714 9884 3724 9940
rect 3780 9884 4844 9940
rect 4900 9884 6300 9940
rect 6356 9884 6366 9940
rect 4722 9772 4732 9828
rect 4788 9772 8204 9828
rect 8260 9772 8270 9828
rect 17826 9772 17836 9828
rect 17892 9772 17902 9828
rect 19058 9772 19068 9828
rect 19124 9772 19292 9828
rect 19348 9772 20188 9828
rect 20244 9772 20524 9828
rect 20580 9772 21812 9828
rect 21868 9772 21878 9828
rect 17836 9716 17892 9772
rect 4386 9660 4396 9716
rect 4452 9660 6076 9716
rect 6132 9660 6142 9716
rect 6458 9660 6468 9716
rect 6524 9660 6916 9716
rect 6972 9660 7980 9716
rect 8036 9660 19460 9716
rect 19516 9660 20188 9716
rect 20132 9604 20188 9660
rect 17826 9548 17836 9604
rect 17892 9548 18900 9604
rect 18956 9548 18966 9604
rect 20132 9548 20748 9604
rect 20804 9548 20814 9604
rect 6522 9380 6532 9436
rect 6588 9380 6636 9436
rect 6692 9380 6740 9436
rect 6796 9380 6806 9436
rect 11842 9380 11852 9436
rect 11908 9380 11956 9436
rect 12012 9380 12060 9436
rect 12116 9380 12126 9436
rect 17162 9380 17172 9436
rect 17228 9380 17276 9436
rect 17332 9380 17380 9436
rect 17436 9380 17446 9436
rect 22482 9380 22492 9436
rect 22548 9380 22596 9436
rect 22652 9380 22700 9436
rect 22756 9380 22766 9436
rect 8418 9324 8428 9380
rect 8484 9324 8652 9380
rect 8708 9324 8718 9380
rect 4946 9212 4956 9268
rect 5012 9212 6972 9268
rect 7028 9212 7038 9268
rect 14018 9212 14028 9268
rect 14084 9212 14958 9268
rect 15014 9212 15148 9268
rect 20626 9212 20636 9268
rect 20692 9212 20860 9268
rect 20916 9212 20926 9268
rect 15092 9156 15148 9212
rect 8530 9100 8540 9156
rect 8596 9100 10780 9156
rect 10836 9100 10846 9156
rect 12674 9100 12684 9156
rect 12740 9100 13024 9156
rect 13080 9100 13916 9156
rect 13972 9100 13982 9156
rect 15092 9100 17612 9156
rect 17668 9100 17678 9156
rect 6066 8988 6076 9044
rect 6132 8988 7420 9044
rect 7476 8988 7486 9044
rect 7858 8988 7868 9044
rect 7924 8988 10220 9044
rect 10276 8988 10286 9044
rect 13794 8988 13804 9044
rect 13860 8988 14700 9044
rect 14756 8988 14766 9044
rect 18498 8988 18508 9044
rect 18564 8988 18956 9044
rect 19012 8988 19022 9044
rect 19674 8988 19684 9044
rect 19740 8988 20300 9044
rect 20356 8988 20366 9044
rect 4722 8876 4732 8932
rect 4788 8876 8204 8932
rect 8260 8876 8652 8932
rect 8708 8876 8718 8932
rect 9034 8876 9044 8932
rect 9100 8876 11284 8932
rect 11340 8876 11350 8932
rect 12114 8876 12124 8932
rect 12180 8876 19124 8932
rect 19180 8876 19190 8932
rect 20626 8876 20636 8932
rect 20692 8876 22092 8932
rect 22148 8876 22158 8932
rect 8418 8764 8428 8820
rect 8484 8764 14812 8820
rect 14868 8764 14878 8820
rect 3862 8596 3872 8652
rect 3928 8596 3976 8652
rect 4032 8596 4080 8652
rect 4136 8596 4146 8652
rect 9182 8596 9192 8652
rect 9248 8596 9296 8652
rect 9352 8596 9400 8652
rect 9456 8596 9466 8652
rect 14502 8596 14512 8652
rect 14568 8596 14616 8652
rect 14672 8596 14720 8652
rect 14776 8596 14786 8652
rect 19822 8596 19832 8652
rect 19888 8596 19936 8652
rect 19992 8596 20040 8652
rect 20096 8596 20106 8652
rect 8530 8428 8540 8484
rect 8596 8428 9324 8484
rect 9380 8428 9390 8484
rect 9538 8428 9548 8484
rect 9604 8428 12236 8484
rect 12292 8428 12302 8484
rect 19114 8428 19124 8484
rect 19180 8428 20636 8484
rect 20692 8428 20702 8484
rect 4498 8316 4508 8372
rect 4564 8316 5124 8372
rect 5180 8316 5684 8372
rect 5740 8316 7420 8372
rect 7476 8316 10892 8372
rect 10948 8316 10958 8372
rect 15362 8316 15372 8372
rect 15428 8316 17500 8372
rect 17556 8316 17566 8372
rect 4610 8204 4620 8260
rect 4676 8204 5796 8260
rect 5852 8204 7196 8260
rect 7252 8204 7262 8260
rect 17714 8204 17724 8260
rect 17780 8204 18452 8260
rect 18508 8204 18518 8260
rect 20132 8204 21980 8260
rect 22036 8204 22046 8260
rect 18330 8092 18340 8148
rect 18396 8092 18844 8148
rect 18900 8092 19292 8148
rect 19348 8092 19358 8148
rect 20132 8036 20188 8204
rect 21578 8092 21588 8148
rect 21644 8092 22316 8148
rect 22372 8092 22382 8148
rect 14242 7980 14252 8036
rect 14308 7980 20188 8036
rect 20962 7980 20972 8036
rect 21028 7980 22204 8036
rect 22260 7980 22270 8036
rect 6522 7812 6532 7868
rect 6588 7812 6636 7868
rect 6692 7812 6740 7868
rect 6796 7812 6806 7868
rect 11842 7812 11852 7868
rect 11908 7812 11956 7868
rect 12012 7812 12060 7868
rect 12116 7812 12126 7868
rect 17162 7812 17172 7868
rect 17228 7812 17276 7868
rect 17332 7812 17380 7868
rect 17436 7812 17446 7868
rect 22482 7812 22492 7868
rect 22548 7812 22596 7868
rect 22652 7812 22700 7868
rect 22756 7812 22766 7868
rect 3882 7644 3892 7700
rect 3948 7644 4676 7700
rect 4732 7644 7644 7700
rect 7700 7644 9268 7700
rect 9324 7644 9334 7700
rect 17882 7644 17892 7700
rect 17948 7644 19068 7700
rect 19124 7644 19134 7700
rect 23200 7476 24000 7504
rect 4498 7420 4508 7476
rect 4564 7420 4956 7476
rect 5012 7420 5236 7476
rect 5292 7420 5302 7476
rect 22306 7420 22316 7476
rect 22372 7420 24000 7476
rect 23200 7392 24000 7420
rect 19506 7308 19516 7364
rect 19572 7308 20412 7364
rect 20468 7308 20478 7364
rect 3862 7028 3872 7084
rect 3928 7028 3976 7084
rect 4032 7028 4080 7084
rect 4136 7028 4146 7084
rect 9182 7028 9192 7084
rect 9248 7028 9296 7084
rect 9352 7028 9400 7084
rect 9456 7028 9466 7084
rect 14502 7028 14512 7084
rect 14568 7028 14616 7084
rect 14672 7028 14720 7084
rect 14776 7028 14786 7084
rect 19822 7028 19832 7084
rect 19888 7028 19936 7084
rect 19992 7028 20040 7084
rect 20096 7028 20106 7084
rect 13346 6860 13356 6916
rect 13412 6860 14588 6916
rect 14644 6860 14654 6916
rect 8194 6636 8204 6692
rect 8260 6636 9996 6692
rect 10052 6636 10062 6692
rect 11106 6636 11116 6692
rect 11172 6636 13580 6692
rect 13636 6636 13646 6692
rect 7970 6300 7980 6356
rect 8036 6300 8204 6356
rect 8260 6300 8270 6356
rect 6522 6244 6532 6300
rect 6588 6244 6636 6300
rect 6692 6244 6740 6300
rect 6796 6244 6806 6300
rect 11842 6244 11852 6300
rect 11908 6244 11956 6300
rect 12012 6244 12060 6300
rect 12116 6244 12126 6300
rect 17162 6244 17172 6300
rect 17228 6244 17276 6300
rect 17332 6244 17380 6300
rect 17436 6244 17446 6300
rect 22482 6244 22492 6300
rect 22548 6244 22596 6300
rect 22652 6244 22700 6300
rect 22756 6244 22766 6300
rect 3845 5852 3855 5908
rect 3911 5852 6804 5908
rect 6860 5852 6870 5908
rect 7074 5852 7084 5908
rect 7140 5852 8204 5908
rect 8260 5852 8876 5908
rect 8932 5852 8942 5908
rect 14466 5852 14476 5908
rect 14532 5852 16828 5908
rect 16884 5852 16894 5908
rect 20066 5852 20076 5908
rect 20132 5852 20300 5908
rect 20356 5852 20366 5908
rect 13514 5740 13524 5796
rect 13580 5740 15372 5796
rect 15428 5740 15438 5796
rect 15922 5740 15932 5796
rect 15988 5740 20860 5796
rect 20916 5740 20926 5796
rect 20300 5684 20356 5740
rect 7298 5628 7308 5684
rect 7364 5628 7812 5684
rect 7868 5628 7878 5684
rect 12338 5628 12348 5684
rect 12404 5628 15596 5684
rect 15652 5628 15662 5684
rect 20290 5628 20300 5684
rect 20356 5628 20366 5684
rect 3602 5516 3612 5572
rect 3668 5516 3678 5572
rect 17154 5516 17164 5572
rect 17220 5516 18508 5572
rect 18564 5516 18574 5572
rect 3612 5124 3668 5516
rect 3862 5460 3872 5516
rect 3928 5460 3976 5516
rect 4032 5460 4080 5516
rect 4136 5460 4146 5516
rect 9182 5460 9192 5516
rect 9248 5460 9296 5516
rect 9352 5460 9400 5516
rect 9456 5460 9466 5516
rect 14502 5460 14512 5516
rect 14568 5460 14616 5516
rect 14672 5460 14720 5516
rect 14776 5460 14786 5516
rect 19822 5460 19832 5516
rect 19888 5460 19936 5516
rect 19992 5460 20040 5516
rect 20096 5460 20106 5516
rect 16818 5404 16828 5460
rect 16884 5404 19684 5460
rect 19628 5348 19684 5404
rect 7970 5292 7980 5348
rect 8036 5292 9604 5348
rect 9660 5292 9670 5348
rect 11554 5292 11564 5348
rect 11620 5292 11900 5348
rect 11956 5292 12684 5348
rect 12740 5292 12750 5348
rect 14018 5292 14028 5348
rect 14084 5292 18620 5348
rect 18676 5292 19404 5348
rect 19460 5292 19470 5348
rect 19628 5292 20020 5348
rect 7634 5180 7644 5236
rect 7700 5180 8652 5236
rect 8708 5180 9212 5236
rect 9268 5180 12348 5236
rect 12404 5180 12414 5236
rect 12562 5180 12572 5236
rect 12628 5180 17164 5236
rect 17220 5180 17230 5236
rect 17826 5180 17836 5236
rect 17892 5180 19292 5236
rect 19348 5180 19358 5236
rect 3602 5068 3612 5124
rect 3668 5068 3678 5124
rect 4610 5068 4620 5124
rect 4676 5068 6748 5124
rect 6804 5068 6814 5124
rect 7186 5068 7196 5124
rect 7252 5068 10668 5124
rect 10724 5068 10734 5124
rect 11218 5068 11228 5124
rect 11284 5068 11676 5124
rect 11732 5068 11742 5124
rect 12002 5068 12012 5124
rect 12068 5068 12236 5124
rect 12292 5068 12302 5124
rect 13794 5068 13804 5124
rect 13860 5068 13870 5124
rect 18050 5068 18060 5124
rect 18116 5068 18844 5124
rect 18900 5068 19796 5124
rect 13804 5012 13860 5068
rect 19740 5012 19796 5068
rect 7746 4956 7756 5012
rect 7812 4956 8708 5012
rect 8764 4956 8774 5012
rect 13570 4956 13580 5012
rect 13636 4956 13860 5012
rect 19730 4956 19740 5012
rect 19796 4956 19806 5012
rect 19964 4956 20020 5292
rect 20850 5180 20860 5236
rect 20916 5180 21980 5236
rect 22036 5180 22046 5236
rect 21578 5068 21588 5124
rect 21644 5068 22316 5124
rect 22372 5068 22382 5124
rect 20076 4956 20086 5012
rect 3042 4844 3052 4900
rect 3108 4844 4956 4900
rect 5012 4844 11340 4900
rect 11396 4844 11406 4900
rect 12562 4844 12572 4900
rect 12628 4844 17724 4900
rect 17780 4844 17790 4900
rect 6522 4676 6532 4732
rect 6588 4676 6636 4732
rect 6692 4676 6740 4732
rect 6796 4676 6806 4732
rect 11842 4676 11852 4732
rect 11908 4676 11956 4732
rect 12012 4676 12060 4732
rect 12116 4676 12126 4732
rect 17162 4676 17172 4732
rect 17228 4676 17276 4732
rect 17332 4676 17380 4732
rect 17436 4676 17446 4732
rect 22482 4676 22492 4732
rect 22548 4676 22596 4732
rect 22652 4676 22700 4732
rect 22756 4676 22766 4732
rect 23200 4564 24000 4592
rect 7074 4508 7084 4564
rect 7140 4508 7756 4564
rect 7812 4508 13636 4564
rect 13692 4508 13702 4564
rect 15250 4508 15260 4564
rect 15316 4508 17444 4564
rect 17500 4508 17510 4564
rect 22306 4508 22316 4564
rect 22372 4508 24000 4564
rect 23200 4480 24000 4508
rect 20514 4284 20524 4340
rect 20580 4284 21196 4340
rect 21252 4284 21700 4340
rect 21756 4284 21766 4340
rect 3862 3892 3872 3948
rect 3928 3892 3976 3948
rect 4032 3892 4080 3948
rect 4136 3892 4146 3948
rect 9182 3892 9192 3948
rect 9248 3892 9296 3948
rect 9352 3892 9400 3948
rect 9456 3892 9466 3948
rect 14502 3892 14512 3948
rect 14568 3892 14616 3948
rect 14672 3892 14720 3948
rect 14776 3892 14786 3948
rect 19822 3892 19832 3948
rect 19888 3892 19936 3948
rect 19992 3892 20040 3948
rect 20096 3892 20106 3948
rect 6522 3108 6532 3164
rect 6588 3108 6636 3164
rect 6692 3108 6740 3164
rect 6796 3108 6806 3164
rect 11842 3108 11852 3164
rect 11908 3108 11956 3164
rect 12012 3108 12060 3164
rect 12116 3108 12126 3164
rect 17162 3108 17172 3164
rect 17228 3108 17276 3164
rect 17332 3108 17380 3164
rect 17436 3108 17446 3164
rect 22482 3108 22492 3164
rect 22548 3108 22596 3164
rect 22652 3108 22700 3164
rect 22756 3108 22766 3164
rect 23200 1652 24000 1680
rect 21746 1596 21756 1652
rect 21812 1596 24000 1652
rect 23200 1568 24000 1596
<< via3 >>
rect 6532 20356 6588 20412
rect 6636 20356 6692 20412
rect 6740 20356 6796 20412
rect 11852 20356 11908 20412
rect 11956 20356 12012 20412
rect 12060 20356 12116 20412
rect 17172 20356 17228 20412
rect 17276 20356 17332 20412
rect 17380 20356 17436 20412
rect 22492 20356 22548 20412
rect 22596 20356 22652 20412
rect 22700 20356 22756 20412
rect 3872 19572 3928 19628
rect 3976 19572 4032 19628
rect 4080 19572 4136 19628
rect 9192 19572 9248 19628
rect 9296 19572 9352 19628
rect 9400 19572 9456 19628
rect 14512 19572 14568 19628
rect 14616 19572 14672 19628
rect 14720 19572 14776 19628
rect 19832 19572 19888 19628
rect 19936 19572 19992 19628
rect 20040 19572 20096 19628
rect 6532 18788 6588 18844
rect 6636 18788 6692 18844
rect 6740 18788 6796 18844
rect 11852 18788 11908 18844
rect 11956 18788 12012 18844
rect 12060 18788 12116 18844
rect 17172 18788 17228 18844
rect 17276 18788 17332 18844
rect 17380 18788 17436 18844
rect 22492 18788 22548 18844
rect 22596 18788 22652 18844
rect 22700 18788 22756 18844
rect 3872 18004 3928 18060
rect 3976 18004 4032 18060
rect 4080 18004 4136 18060
rect 9192 18004 9248 18060
rect 9296 18004 9352 18060
rect 9400 18004 9456 18060
rect 14512 18004 14568 18060
rect 14616 18004 14672 18060
rect 14720 18004 14776 18060
rect 19832 18004 19888 18060
rect 19936 18004 19992 18060
rect 20040 18004 20096 18060
rect 6532 17220 6588 17276
rect 6636 17220 6692 17276
rect 6740 17220 6796 17276
rect 11852 17220 11908 17276
rect 11956 17220 12012 17276
rect 12060 17220 12116 17276
rect 17172 17220 17228 17276
rect 17276 17220 17332 17276
rect 17380 17220 17436 17276
rect 22492 17220 22548 17276
rect 22596 17220 22652 17276
rect 22700 17220 22756 17276
rect 3872 16436 3928 16492
rect 3976 16436 4032 16492
rect 4080 16436 4136 16492
rect 9192 16436 9248 16492
rect 9296 16436 9352 16492
rect 9400 16436 9456 16492
rect 14512 16436 14568 16492
rect 14616 16436 14672 16492
rect 14720 16436 14776 16492
rect 19832 16436 19888 16492
rect 19936 16436 19992 16492
rect 20040 16436 20096 16492
rect 6532 15652 6588 15708
rect 6636 15652 6692 15708
rect 6740 15652 6796 15708
rect 11852 15652 11908 15708
rect 11956 15652 12012 15708
rect 12060 15652 12116 15708
rect 17172 15652 17228 15708
rect 17276 15652 17332 15708
rect 17380 15652 17436 15708
rect 22492 15652 22548 15708
rect 22596 15652 22652 15708
rect 22700 15652 22756 15708
rect 3872 14868 3928 14924
rect 3976 14868 4032 14924
rect 4080 14868 4136 14924
rect 9192 14868 9248 14924
rect 9296 14868 9352 14924
rect 9400 14868 9456 14924
rect 14512 14868 14568 14924
rect 14616 14868 14672 14924
rect 14720 14868 14776 14924
rect 19832 14868 19888 14924
rect 19936 14868 19992 14924
rect 20040 14868 20096 14924
rect 6532 14084 6588 14140
rect 6636 14084 6692 14140
rect 6740 14084 6796 14140
rect 11852 14084 11908 14140
rect 11956 14084 12012 14140
rect 12060 14084 12116 14140
rect 17172 14084 17228 14140
rect 17276 14084 17332 14140
rect 17380 14084 17436 14140
rect 22492 14084 22548 14140
rect 22596 14084 22652 14140
rect 22700 14084 22756 14140
rect 3872 13300 3928 13356
rect 3976 13300 4032 13356
rect 4080 13300 4136 13356
rect 9192 13300 9248 13356
rect 9296 13300 9352 13356
rect 9400 13300 9456 13356
rect 14512 13300 14568 13356
rect 14616 13300 14672 13356
rect 14720 13300 14776 13356
rect 19832 13300 19888 13356
rect 19936 13300 19992 13356
rect 20040 13300 20096 13356
rect 10332 13020 10388 13076
rect 6532 12516 6588 12572
rect 6636 12516 6692 12572
rect 6740 12516 6796 12572
rect 11852 12516 11908 12572
rect 11956 12516 12012 12572
rect 12060 12516 12116 12572
rect 17172 12516 17228 12572
rect 17276 12516 17332 12572
rect 17380 12516 17436 12572
rect 22492 12516 22548 12572
rect 22596 12516 22652 12572
rect 22700 12516 22756 12572
rect 10332 12236 10388 12292
rect 3872 11732 3928 11788
rect 3976 11732 4032 11788
rect 4080 11732 4136 11788
rect 9192 11732 9248 11788
rect 9296 11732 9352 11788
rect 9400 11732 9456 11788
rect 14512 11732 14568 11788
rect 14616 11732 14672 11788
rect 14720 11732 14776 11788
rect 19832 11732 19888 11788
rect 19936 11732 19992 11788
rect 20040 11732 20096 11788
rect 6532 10948 6588 11004
rect 6636 10948 6692 11004
rect 6740 10948 6796 11004
rect 11852 10948 11908 11004
rect 11956 10948 12012 11004
rect 12060 10948 12116 11004
rect 17172 10948 17228 11004
rect 17276 10948 17332 11004
rect 17380 10948 17436 11004
rect 22492 10948 22548 11004
rect 22596 10948 22652 11004
rect 22700 10948 22756 11004
rect 3872 10164 3928 10220
rect 3976 10164 4032 10220
rect 4080 10164 4136 10220
rect 9192 10164 9248 10220
rect 9296 10164 9352 10220
rect 9400 10164 9456 10220
rect 14512 10164 14568 10220
rect 14616 10164 14672 10220
rect 14720 10164 14776 10220
rect 19832 10164 19888 10220
rect 19936 10164 19992 10220
rect 20040 10164 20096 10220
rect 6532 9380 6588 9436
rect 6636 9380 6692 9436
rect 6740 9380 6796 9436
rect 11852 9380 11908 9436
rect 11956 9380 12012 9436
rect 12060 9380 12116 9436
rect 17172 9380 17228 9436
rect 17276 9380 17332 9436
rect 17380 9380 17436 9436
rect 22492 9380 22548 9436
rect 22596 9380 22652 9436
rect 22700 9380 22756 9436
rect 3872 8596 3928 8652
rect 3976 8596 4032 8652
rect 4080 8596 4136 8652
rect 9192 8596 9248 8652
rect 9296 8596 9352 8652
rect 9400 8596 9456 8652
rect 14512 8596 14568 8652
rect 14616 8596 14672 8652
rect 14720 8596 14776 8652
rect 19832 8596 19888 8652
rect 19936 8596 19992 8652
rect 20040 8596 20096 8652
rect 6532 7812 6588 7868
rect 6636 7812 6692 7868
rect 6740 7812 6796 7868
rect 11852 7812 11908 7868
rect 11956 7812 12012 7868
rect 12060 7812 12116 7868
rect 17172 7812 17228 7868
rect 17276 7812 17332 7868
rect 17380 7812 17436 7868
rect 22492 7812 22548 7868
rect 22596 7812 22652 7868
rect 22700 7812 22756 7868
rect 3872 7028 3928 7084
rect 3976 7028 4032 7084
rect 4080 7028 4136 7084
rect 9192 7028 9248 7084
rect 9296 7028 9352 7084
rect 9400 7028 9456 7084
rect 14512 7028 14568 7084
rect 14616 7028 14672 7084
rect 14720 7028 14776 7084
rect 19832 7028 19888 7084
rect 19936 7028 19992 7084
rect 20040 7028 20096 7084
rect 6532 6244 6588 6300
rect 6636 6244 6692 6300
rect 6740 6244 6796 6300
rect 11852 6244 11908 6300
rect 11956 6244 12012 6300
rect 12060 6244 12116 6300
rect 17172 6244 17228 6300
rect 17276 6244 17332 6300
rect 17380 6244 17436 6300
rect 22492 6244 22548 6300
rect 22596 6244 22652 6300
rect 22700 6244 22756 6300
rect 3872 5460 3928 5516
rect 3976 5460 4032 5516
rect 4080 5460 4136 5516
rect 9192 5460 9248 5516
rect 9296 5460 9352 5516
rect 9400 5460 9456 5516
rect 14512 5460 14568 5516
rect 14616 5460 14672 5516
rect 14720 5460 14776 5516
rect 19832 5460 19888 5516
rect 19936 5460 19992 5516
rect 20040 5460 20096 5516
rect 6532 4676 6588 4732
rect 6636 4676 6692 4732
rect 6740 4676 6796 4732
rect 11852 4676 11908 4732
rect 11956 4676 12012 4732
rect 12060 4676 12116 4732
rect 17172 4676 17228 4732
rect 17276 4676 17332 4732
rect 17380 4676 17436 4732
rect 22492 4676 22548 4732
rect 22596 4676 22652 4732
rect 22700 4676 22756 4732
rect 3872 3892 3928 3948
rect 3976 3892 4032 3948
rect 4080 3892 4136 3948
rect 9192 3892 9248 3948
rect 9296 3892 9352 3948
rect 9400 3892 9456 3948
rect 14512 3892 14568 3948
rect 14616 3892 14672 3948
rect 14720 3892 14776 3948
rect 19832 3892 19888 3948
rect 19936 3892 19992 3948
rect 20040 3892 20096 3948
rect 6532 3108 6588 3164
rect 6636 3108 6692 3164
rect 6740 3108 6796 3164
rect 11852 3108 11908 3164
rect 11956 3108 12012 3164
rect 12060 3108 12116 3164
rect 17172 3108 17228 3164
rect 17276 3108 17332 3164
rect 17380 3108 17436 3164
rect 22492 3108 22548 3164
rect 22596 3108 22652 3164
rect 22700 3108 22756 3164
<< metal4 >>
rect 3844 19628 4164 20444
rect 3844 19572 3872 19628
rect 3928 19572 3976 19628
rect 4032 19572 4080 19628
rect 4136 19572 4164 19628
rect 3844 18060 4164 19572
rect 3844 18004 3872 18060
rect 3928 18004 3976 18060
rect 4032 18004 4080 18060
rect 4136 18004 4164 18060
rect 3844 16492 4164 18004
rect 3844 16436 3872 16492
rect 3928 16436 3976 16492
rect 4032 16436 4080 16492
rect 4136 16436 4164 16492
rect 3844 14924 4164 16436
rect 3844 14868 3872 14924
rect 3928 14868 3976 14924
rect 4032 14868 4080 14924
rect 4136 14868 4164 14924
rect 3844 13356 4164 14868
rect 3844 13300 3872 13356
rect 3928 13300 3976 13356
rect 4032 13300 4080 13356
rect 4136 13300 4164 13356
rect 3844 11788 4164 13300
rect 3844 11732 3872 11788
rect 3928 11732 3976 11788
rect 4032 11732 4080 11788
rect 4136 11732 4164 11788
rect 3844 10220 4164 11732
rect 3844 10164 3872 10220
rect 3928 10164 3976 10220
rect 4032 10164 4080 10220
rect 4136 10164 4164 10220
rect 3844 8652 4164 10164
rect 3844 8596 3872 8652
rect 3928 8596 3976 8652
rect 4032 8596 4080 8652
rect 4136 8596 4164 8652
rect 3844 7084 4164 8596
rect 3844 7028 3872 7084
rect 3928 7028 3976 7084
rect 4032 7028 4080 7084
rect 4136 7028 4164 7084
rect 3844 5516 4164 7028
rect 3844 5460 3872 5516
rect 3928 5460 3976 5516
rect 4032 5460 4080 5516
rect 4136 5460 4164 5516
rect 3844 3948 4164 5460
rect 3844 3892 3872 3948
rect 3928 3892 3976 3948
rect 4032 3892 4080 3948
rect 4136 3892 4164 3948
rect 3844 3076 4164 3892
rect 6504 20412 6824 20444
rect 6504 20356 6532 20412
rect 6588 20356 6636 20412
rect 6692 20356 6740 20412
rect 6796 20356 6824 20412
rect 6504 18844 6824 20356
rect 6504 18788 6532 18844
rect 6588 18788 6636 18844
rect 6692 18788 6740 18844
rect 6796 18788 6824 18844
rect 6504 17276 6824 18788
rect 6504 17220 6532 17276
rect 6588 17220 6636 17276
rect 6692 17220 6740 17276
rect 6796 17220 6824 17276
rect 6504 15708 6824 17220
rect 6504 15652 6532 15708
rect 6588 15652 6636 15708
rect 6692 15652 6740 15708
rect 6796 15652 6824 15708
rect 6504 14140 6824 15652
rect 6504 14084 6532 14140
rect 6588 14084 6636 14140
rect 6692 14084 6740 14140
rect 6796 14084 6824 14140
rect 6504 12572 6824 14084
rect 6504 12516 6532 12572
rect 6588 12516 6636 12572
rect 6692 12516 6740 12572
rect 6796 12516 6824 12572
rect 6504 11004 6824 12516
rect 6504 10948 6532 11004
rect 6588 10948 6636 11004
rect 6692 10948 6740 11004
rect 6796 10948 6824 11004
rect 6504 9436 6824 10948
rect 6504 9380 6532 9436
rect 6588 9380 6636 9436
rect 6692 9380 6740 9436
rect 6796 9380 6824 9436
rect 6504 7868 6824 9380
rect 6504 7812 6532 7868
rect 6588 7812 6636 7868
rect 6692 7812 6740 7868
rect 6796 7812 6824 7868
rect 6504 6300 6824 7812
rect 6504 6244 6532 6300
rect 6588 6244 6636 6300
rect 6692 6244 6740 6300
rect 6796 6244 6824 6300
rect 6504 4732 6824 6244
rect 6504 4676 6532 4732
rect 6588 4676 6636 4732
rect 6692 4676 6740 4732
rect 6796 4676 6824 4732
rect 6504 3164 6824 4676
rect 6504 3108 6532 3164
rect 6588 3108 6636 3164
rect 6692 3108 6740 3164
rect 6796 3108 6824 3164
rect 6504 3076 6824 3108
rect 9164 19628 9484 20444
rect 9164 19572 9192 19628
rect 9248 19572 9296 19628
rect 9352 19572 9400 19628
rect 9456 19572 9484 19628
rect 9164 18060 9484 19572
rect 9164 18004 9192 18060
rect 9248 18004 9296 18060
rect 9352 18004 9400 18060
rect 9456 18004 9484 18060
rect 9164 16492 9484 18004
rect 9164 16436 9192 16492
rect 9248 16436 9296 16492
rect 9352 16436 9400 16492
rect 9456 16436 9484 16492
rect 9164 14924 9484 16436
rect 9164 14868 9192 14924
rect 9248 14868 9296 14924
rect 9352 14868 9400 14924
rect 9456 14868 9484 14924
rect 9164 13356 9484 14868
rect 9164 13300 9192 13356
rect 9248 13300 9296 13356
rect 9352 13300 9400 13356
rect 9456 13300 9484 13356
rect 9164 11788 9484 13300
rect 11824 20412 12144 20444
rect 11824 20356 11852 20412
rect 11908 20356 11956 20412
rect 12012 20356 12060 20412
rect 12116 20356 12144 20412
rect 11824 18844 12144 20356
rect 11824 18788 11852 18844
rect 11908 18788 11956 18844
rect 12012 18788 12060 18844
rect 12116 18788 12144 18844
rect 11824 17276 12144 18788
rect 11824 17220 11852 17276
rect 11908 17220 11956 17276
rect 12012 17220 12060 17276
rect 12116 17220 12144 17276
rect 11824 15708 12144 17220
rect 11824 15652 11852 15708
rect 11908 15652 11956 15708
rect 12012 15652 12060 15708
rect 12116 15652 12144 15708
rect 11824 14140 12144 15652
rect 11824 14084 11852 14140
rect 11908 14084 11956 14140
rect 12012 14084 12060 14140
rect 12116 14084 12144 14140
rect 10332 13076 10388 13086
rect 10332 12292 10388 13020
rect 10332 12226 10388 12236
rect 11824 12572 12144 14084
rect 11824 12516 11852 12572
rect 11908 12516 11956 12572
rect 12012 12516 12060 12572
rect 12116 12516 12144 12572
rect 9164 11732 9192 11788
rect 9248 11732 9296 11788
rect 9352 11732 9400 11788
rect 9456 11732 9484 11788
rect 9164 10220 9484 11732
rect 9164 10164 9192 10220
rect 9248 10164 9296 10220
rect 9352 10164 9400 10220
rect 9456 10164 9484 10220
rect 9164 8652 9484 10164
rect 9164 8596 9192 8652
rect 9248 8596 9296 8652
rect 9352 8596 9400 8652
rect 9456 8596 9484 8652
rect 9164 7084 9484 8596
rect 9164 7028 9192 7084
rect 9248 7028 9296 7084
rect 9352 7028 9400 7084
rect 9456 7028 9484 7084
rect 9164 5516 9484 7028
rect 9164 5460 9192 5516
rect 9248 5460 9296 5516
rect 9352 5460 9400 5516
rect 9456 5460 9484 5516
rect 9164 3948 9484 5460
rect 9164 3892 9192 3948
rect 9248 3892 9296 3948
rect 9352 3892 9400 3948
rect 9456 3892 9484 3948
rect 9164 3076 9484 3892
rect 11824 11004 12144 12516
rect 11824 10948 11852 11004
rect 11908 10948 11956 11004
rect 12012 10948 12060 11004
rect 12116 10948 12144 11004
rect 11824 9436 12144 10948
rect 11824 9380 11852 9436
rect 11908 9380 11956 9436
rect 12012 9380 12060 9436
rect 12116 9380 12144 9436
rect 11824 7868 12144 9380
rect 11824 7812 11852 7868
rect 11908 7812 11956 7868
rect 12012 7812 12060 7868
rect 12116 7812 12144 7868
rect 11824 6300 12144 7812
rect 11824 6244 11852 6300
rect 11908 6244 11956 6300
rect 12012 6244 12060 6300
rect 12116 6244 12144 6300
rect 11824 4732 12144 6244
rect 11824 4676 11852 4732
rect 11908 4676 11956 4732
rect 12012 4676 12060 4732
rect 12116 4676 12144 4732
rect 11824 3164 12144 4676
rect 11824 3108 11852 3164
rect 11908 3108 11956 3164
rect 12012 3108 12060 3164
rect 12116 3108 12144 3164
rect 11824 3076 12144 3108
rect 14484 19628 14804 20444
rect 14484 19572 14512 19628
rect 14568 19572 14616 19628
rect 14672 19572 14720 19628
rect 14776 19572 14804 19628
rect 14484 18060 14804 19572
rect 14484 18004 14512 18060
rect 14568 18004 14616 18060
rect 14672 18004 14720 18060
rect 14776 18004 14804 18060
rect 14484 16492 14804 18004
rect 14484 16436 14512 16492
rect 14568 16436 14616 16492
rect 14672 16436 14720 16492
rect 14776 16436 14804 16492
rect 14484 14924 14804 16436
rect 14484 14868 14512 14924
rect 14568 14868 14616 14924
rect 14672 14868 14720 14924
rect 14776 14868 14804 14924
rect 14484 13356 14804 14868
rect 14484 13300 14512 13356
rect 14568 13300 14616 13356
rect 14672 13300 14720 13356
rect 14776 13300 14804 13356
rect 14484 11788 14804 13300
rect 14484 11732 14512 11788
rect 14568 11732 14616 11788
rect 14672 11732 14720 11788
rect 14776 11732 14804 11788
rect 14484 10220 14804 11732
rect 14484 10164 14512 10220
rect 14568 10164 14616 10220
rect 14672 10164 14720 10220
rect 14776 10164 14804 10220
rect 14484 8652 14804 10164
rect 14484 8596 14512 8652
rect 14568 8596 14616 8652
rect 14672 8596 14720 8652
rect 14776 8596 14804 8652
rect 14484 7084 14804 8596
rect 14484 7028 14512 7084
rect 14568 7028 14616 7084
rect 14672 7028 14720 7084
rect 14776 7028 14804 7084
rect 14484 5516 14804 7028
rect 14484 5460 14512 5516
rect 14568 5460 14616 5516
rect 14672 5460 14720 5516
rect 14776 5460 14804 5516
rect 14484 3948 14804 5460
rect 14484 3892 14512 3948
rect 14568 3892 14616 3948
rect 14672 3892 14720 3948
rect 14776 3892 14804 3948
rect 14484 3076 14804 3892
rect 17144 20412 17464 20444
rect 17144 20356 17172 20412
rect 17228 20356 17276 20412
rect 17332 20356 17380 20412
rect 17436 20356 17464 20412
rect 17144 18844 17464 20356
rect 17144 18788 17172 18844
rect 17228 18788 17276 18844
rect 17332 18788 17380 18844
rect 17436 18788 17464 18844
rect 17144 17276 17464 18788
rect 17144 17220 17172 17276
rect 17228 17220 17276 17276
rect 17332 17220 17380 17276
rect 17436 17220 17464 17276
rect 17144 15708 17464 17220
rect 17144 15652 17172 15708
rect 17228 15652 17276 15708
rect 17332 15652 17380 15708
rect 17436 15652 17464 15708
rect 17144 14140 17464 15652
rect 17144 14084 17172 14140
rect 17228 14084 17276 14140
rect 17332 14084 17380 14140
rect 17436 14084 17464 14140
rect 17144 12572 17464 14084
rect 17144 12516 17172 12572
rect 17228 12516 17276 12572
rect 17332 12516 17380 12572
rect 17436 12516 17464 12572
rect 17144 11004 17464 12516
rect 17144 10948 17172 11004
rect 17228 10948 17276 11004
rect 17332 10948 17380 11004
rect 17436 10948 17464 11004
rect 17144 9436 17464 10948
rect 17144 9380 17172 9436
rect 17228 9380 17276 9436
rect 17332 9380 17380 9436
rect 17436 9380 17464 9436
rect 17144 7868 17464 9380
rect 17144 7812 17172 7868
rect 17228 7812 17276 7868
rect 17332 7812 17380 7868
rect 17436 7812 17464 7868
rect 17144 6300 17464 7812
rect 17144 6244 17172 6300
rect 17228 6244 17276 6300
rect 17332 6244 17380 6300
rect 17436 6244 17464 6300
rect 17144 4732 17464 6244
rect 17144 4676 17172 4732
rect 17228 4676 17276 4732
rect 17332 4676 17380 4732
rect 17436 4676 17464 4732
rect 17144 3164 17464 4676
rect 17144 3108 17172 3164
rect 17228 3108 17276 3164
rect 17332 3108 17380 3164
rect 17436 3108 17464 3164
rect 17144 3076 17464 3108
rect 19804 19628 20124 20444
rect 19804 19572 19832 19628
rect 19888 19572 19936 19628
rect 19992 19572 20040 19628
rect 20096 19572 20124 19628
rect 19804 18060 20124 19572
rect 19804 18004 19832 18060
rect 19888 18004 19936 18060
rect 19992 18004 20040 18060
rect 20096 18004 20124 18060
rect 19804 16492 20124 18004
rect 19804 16436 19832 16492
rect 19888 16436 19936 16492
rect 19992 16436 20040 16492
rect 20096 16436 20124 16492
rect 19804 14924 20124 16436
rect 19804 14868 19832 14924
rect 19888 14868 19936 14924
rect 19992 14868 20040 14924
rect 20096 14868 20124 14924
rect 19804 13356 20124 14868
rect 19804 13300 19832 13356
rect 19888 13300 19936 13356
rect 19992 13300 20040 13356
rect 20096 13300 20124 13356
rect 19804 11788 20124 13300
rect 19804 11732 19832 11788
rect 19888 11732 19936 11788
rect 19992 11732 20040 11788
rect 20096 11732 20124 11788
rect 19804 10220 20124 11732
rect 19804 10164 19832 10220
rect 19888 10164 19936 10220
rect 19992 10164 20040 10220
rect 20096 10164 20124 10220
rect 19804 8652 20124 10164
rect 19804 8596 19832 8652
rect 19888 8596 19936 8652
rect 19992 8596 20040 8652
rect 20096 8596 20124 8652
rect 19804 7084 20124 8596
rect 19804 7028 19832 7084
rect 19888 7028 19936 7084
rect 19992 7028 20040 7084
rect 20096 7028 20124 7084
rect 19804 5516 20124 7028
rect 19804 5460 19832 5516
rect 19888 5460 19936 5516
rect 19992 5460 20040 5516
rect 20096 5460 20124 5516
rect 19804 3948 20124 5460
rect 19804 3892 19832 3948
rect 19888 3892 19936 3948
rect 19992 3892 20040 3948
rect 20096 3892 20124 3948
rect 19804 3076 20124 3892
rect 22464 20412 22784 20444
rect 22464 20356 22492 20412
rect 22548 20356 22596 20412
rect 22652 20356 22700 20412
rect 22756 20356 22784 20412
rect 22464 18844 22784 20356
rect 22464 18788 22492 18844
rect 22548 18788 22596 18844
rect 22652 18788 22700 18844
rect 22756 18788 22784 18844
rect 22464 17276 22784 18788
rect 22464 17220 22492 17276
rect 22548 17220 22596 17276
rect 22652 17220 22700 17276
rect 22756 17220 22784 17276
rect 22464 15708 22784 17220
rect 22464 15652 22492 15708
rect 22548 15652 22596 15708
rect 22652 15652 22700 15708
rect 22756 15652 22784 15708
rect 22464 14140 22784 15652
rect 22464 14084 22492 14140
rect 22548 14084 22596 14140
rect 22652 14084 22700 14140
rect 22756 14084 22784 14140
rect 22464 12572 22784 14084
rect 22464 12516 22492 12572
rect 22548 12516 22596 12572
rect 22652 12516 22700 12572
rect 22756 12516 22784 12572
rect 22464 11004 22784 12516
rect 22464 10948 22492 11004
rect 22548 10948 22596 11004
rect 22652 10948 22700 11004
rect 22756 10948 22784 11004
rect 22464 9436 22784 10948
rect 22464 9380 22492 9436
rect 22548 9380 22596 9436
rect 22652 9380 22700 9436
rect 22756 9380 22784 9436
rect 22464 7868 22784 9380
rect 22464 7812 22492 7868
rect 22548 7812 22596 7868
rect 22652 7812 22700 7868
rect 22756 7812 22784 7868
rect 22464 6300 22784 7812
rect 22464 6244 22492 6300
rect 22548 6244 22596 6300
rect 22652 6244 22700 6300
rect 22756 6244 22784 6300
rect 22464 4732 22784 6244
rect 22464 4676 22492 4732
rect 22548 4676 22596 4732
rect 22652 4676 22700 4732
rect 22756 4676 22784 4732
rect 22464 3164 22784 4676
rect 22464 3108 22492 3164
rect 22548 3108 22596 3164
rect 22652 3108 22700 3164
rect 22756 3108 22784 3164
rect 22464 3076 22784 3108
use gf180mcu_as_sc_mcu7t3v3__buff_2  _102_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751534193
transform -1 0 20944 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _103_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532043
transform 1 0 15120 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _104_
timestamp 1751534193
transform -1 0 4592 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _105_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751740063
transform -1 0 10192 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753182340
transform 1 0 7952 0 -1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _107_
timestamp 1751534193
transform 1 0 9072 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _108_
timestamp 1753182340
transform 1 0 14112 0 1 15680
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _109_
timestamp 1751534193
transform 1 0 15344 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _110_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751531619
transform -1 0 21392 0 -1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _111_
timestamp 1751534193
transform 1 0 17808 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751889808
transform 1 0 18592 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _113_
timestamp 1751740063
transform 1 0 18928 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _114_
timestamp 1751740063
transform 1 0 17472 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _115_
timestamp 1751534193
transform -1 0 11984 0 -1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _116_
timestamp 1753182340
transform 1 0 7952 0 -1 14112
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _117_
timestamp 1751534193
transform 1 0 9408 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _118_
timestamp 1751532043
transform -1 0 13776 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _119_
timestamp 1751532043
transform -1 0 17696 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1752345181
transform -1 0 16128 0 1 4704
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _121_
timestamp 1751534193
transform -1 0 9296 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _122_
timestamp 1751534193
transform -1 0 8176 0 -1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751889408
transform -1 0 20608 0 -1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _124_
timestamp 1751534193
transform 1 0 16800 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _125_
timestamp 1751740063
transform 1 0 19152 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _126_
timestamp 1751531619
transform 1 0 18368 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _127_
timestamp 1751889408
transform 1 0 13776 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _128_
timestamp 1751534193
transform -1 0 14560 0 -1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _129_
timestamp 1753182340
transform 1 0 16240 0 1 12544
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _130_
timestamp 1751534193
transform 1 0 17248 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _131_
timestamp 1751534193
transform -1 0 15456 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _132_
timestamp 1751889408
transform -1 0 14784 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _133_
timestamp 1751889808
transform -1 0 14112 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _134_
timestamp 1751740063
transform 1 0 8288 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _135_
timestamp 1751534193
transform -1 0 8736 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _136_
timestamp 1753182340
transform 1 0 11984 0 -1 15680
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _137_
timestamp 1751889808
transform 1 0 14112 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _138_
timestamp 1751889408
transform 1 0 13888 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _139_
timestamp 1751531619
transform 1 0 14000 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _140_
timestamp 1751532043
transform -1 0 5264 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _141_
timestamp 1751889808
transform 1 0 18816 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _142_
timestamp 1751740063
transform 1 0 18032 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _143_
timestamp 1751740063
transform -1 0 15456 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _144_
timestamp 1751889808
transform -1 0 14112 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _145_
timestamp 1751740063
transform -1 0 7952 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _146_
timestamp 1751889408
transform 1 0 4592 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _147_
timestamp 1751534193
transform -1 0 5264 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _148_
timestamp 1751534193
transform 1 0 20048 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _149_
timestamp 1751534193
transform -1 0 20944 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _150_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753441877
transform -1 0 22288 0 1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _151_
timestamp 1751740063
transform 1 0 19712 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _152_
timestamp 1751889408
transform -1 0 18928 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _153_
timestamp 1751534193
transform -1 0 18144 0 -1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _154_
timestamp 1751740063
transform 1 0 11088 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _155_
timestamp 1751740063
transform 1 0 12096 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _156_
timestamp 1751532043
transform 1 0 11872 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _157_
timestamp 1751534193
transform -1 0 18368 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _158_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753371985
transform -1 0 12880 0 -1 4704
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _159_
timestamp 1751740063
transform 1 0 11760 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _160_
timestamp 1753182340
transform 1 0 13104 0 -1 12544
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _161_
timestamp 1751534193
transform 1 0 17808 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _162_
timestamp 1751889808
transform -1 0 14112 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _163_
timestamp 1751740063
transform -1 0 8064 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _164_
timestamp 1751889408
transform -1 0 5264 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _165_
timestamp 1751740063
transform 1 0 3360 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _166_
timestamp 1751531619
transform -1 0 4928 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _167_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751905124
transform 1 0 2576 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _168_
timestamp 1753371985
transform 1 0 3696 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _169_
timestamp 1751889408
transform 1 0 13328 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _170_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753868718
transform -1 0 14560 0 -1 9408
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _171_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753891287
transform 1 0 11760 0 -1 17248
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _172_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1752061876
transform 1 0 4032 0 -1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _173_
timestamp 1751534193
transform -1 0 8624 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _174_
timestamp 1753371985
transform -1 0 5264 0 1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _175_
timestamp 1751532043
transform 1 0 4480 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _176_
timestamp 1753371985
transform -1 0 8624 0 1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _177_
timestamp 1751531619
transform 1 0 7280 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _178_
timestamp 1751532043
transform 1 0 8176 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _179_
timestamp 1751889808
transform 1 0 11984 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _180_
timestamp 1751905124
transform -1 0 13216 0 -1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _181_
timestamp 1751740063
transform -1 0 9184 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _182_
timestamp 1751889808
transform 1 0 10752 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _183_
timestamp 1753371985
transform 1 0 8064 0 -1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _184_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753960525
transform 1 0 8960 0 1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _185_
timestamp 1753960525
transform -1 0 10528 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _186_
timestamp 1752061876
transform 1 0 8624 0 1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _187_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751914308
transform 1 0 9408 0 -1 9408
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _188_
timestamp 1753441877
transform -1 0 7280 0 -1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _189_
timestamp 1751532043
transform -1 0 3584 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _190_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753277515
transform -1 0 4928 0 -1 6272
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _191_
timestamp 1753277515
transform 1 0 2912 0 -1 4704
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _192_
timestamp 1753277515
transform 1 0 3360 0 1 4704
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _193_
timestamp 1753182340
transform 1 0 11424 0 -1 14112
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _194_
timestamp 1753441877
transform 1 0 7504 0 1 4704
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _195_
timestamp 1753960525
transform -1 0 8736 0 -1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _196_
timestamp 1753371985
transform 1 0 6384 0 1 4704
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_2  _197_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753579406
transform -1 0 12096 0 1 4704
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _198_
timestamp 1751889408
transform -1 0 18816 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _199_
timestamp 1751534193
transform 1 0 18256 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _200_
timestamp 1753441877
transform -1 0 21952 0 -1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _201_
timestamp 1751740063
transform 1 0 18928 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _202_
timestamp 1751532043
transform -1 0 18592 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _203_
timestamp 1753182340
transform -1 0 18816 0 -1 9408
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _204_
timestamp 1753960525
transform 1 0 18816 0 -1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _205_
timestamp 1751534193
transform 1 0 20272 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _206_
timestamp 1751532043
transform -1 0 18144 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _207_
timestamp 1753371985
transform -1 0 19488 0 1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _208_
timestamp 1751532043
transform -1 0 19152 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _209_
timestamp 1751740063
transform 1 0 13440 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _210_
timestamp 1753441877
transform 1 0 14560 0 -1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _211_
timestamp 1753371985
transform 1 0 17248 0 1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _212_
timestamp 1753371985
transform -1 0 21280 0 -1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _213_
timestamp 1751889408
transform 1 0 19264 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _214_
timestamp 1751534193
transform -1 0 19824 0 -1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _215_
timestamp 1751740063
transform 1 0 17584 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _216_
timestamp 1751889408
transform -1 0 4032 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _217_
timestamp 1751534193
transform -1 0 3248 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _218_
timestamp 1752061876
transform -1 0 4144 0 1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _219_
timestamp 1751889408
transform 1 0 13328 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _220_
timestamp 1751534193
transform 1 0 14672 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _221_
timestamp 1751532043
transform -1 0 9632 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _222_
timestamp 1753441877
transform -1 0 9184 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _223_
timestamp 1751531619
transform -1 0 8176 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _224_
timestamp 1752061876
transform 1 0 7840 0 1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _225_
timestamp 1751740063
transform 1 0 7168 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _226_
timestamp 1751531619
transform 1 0 4592 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _227_
timestamp 1753371985
transform 1 0 5488 0 1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _228_
timestamp 1751914308
transform -1 0 4032 0 1 10976
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _229_
timestamp 1751534193
transform 1 0 3136 0 -1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _230_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753272495
transform 1 0 3136 0 -1 7840
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _231_
timestamp 1753441877
transform -1 0 4816 0 1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _232_
timestamp 1753182340
transform 1 0 4032 0 1 10976
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _233_
timestamp 1753371985
transform 1 0 3136 0 -1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _234_
timestamp 1751889808
transform -1 0 21168 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _235_
timestamp 1751889408
transform 1 0 19600 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _236_
timestamp 1751534193
transform 1 0 20048 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _237_
timestamp 1753182340
transform -1 0 21392 0 -1 15680
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _238_
timestamp 1753182340
transform 1 0 19600 0 -1 14112
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _239_
timestamp 1751534193
transform 1 0 21168 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _240_
timestamp 1751740063
transform -1 0 14896 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _241_
timestamp 1751889408
transform -1 0 11424 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _242_
timestamp 1751534193
transform 1 0 10640 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _243_
timestamp 1752061876
transform 1 0 18928 0 1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _244_
timestamp 1751534193
transform -1 0 3472 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _245_
timestamp 1751534193
transform -1 0 4144 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _246_
timestamp 1751534193
transform 1 0 4144 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _247_
timestamp 1751534193
transform 1 0 5488 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _248_
timestamp 1751534193
transform -1 0 11312 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _249_
timestamp 1751534193
transform -1 0 19376 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _250_
timestamp 1751534193
transform 1 0 14784 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _251_
timestamp 1751534193
transform 1 0 16016 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _252_
timestamp 1751534193
transform 1 0 18256 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _253_
timestamp 1751534193
transform 1 0 21168 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__110__A dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532392
transform 1 0 22064 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__111__A
timestamp 1751532392
transform 1 0 19376 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__123__A
timestamp 1751532392
transform 1 0 21616 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__127__A
timestamp 1751532392
transform 1 0 13552 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__139__A
timestamp 1751532392
transform 1 0 15680 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__146__A
timestamp 1751532392
transform 1 0 5600 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__158__C
timestamp 1751532392
transform 1 0 11536 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__164__A
timestamp 1751532392
transform 1 0 5712 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__171__B
timestamp 1751532392
transform 1 0 11536 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__175__A
timestamp 1751532392
transform 1 0 5152 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__191__A
timestamp 1751532392
transform 1 0 4704 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__194__B
timestamp 1751532392
transform -1 0 8848 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__194__C
timestamp 1751532392
transform 1 0 9520 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__219__A
timestamp 1751532392
transform -1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__223__A
timestamp 1751532392
transform 1 0 8400 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__226__B
timestamp 1751532392
transform 1 0 5600 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__227__C
timestamp 1751532392
transform 1 0 6832 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__231__A
timestamp 1751532392
transform 1 0 5712 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__231__B
timestamp 1751532392
transform 1 0 5040 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__238__B
timestamp 1751532392
transform 1 0 21392 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__241__B
timestamp 1751532392
transform -1 0 11648 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__244__A
timestamp 1751532392
transform 1 0 3472 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input1_A
timestamp 1751532392
transform -1 0 21728 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input2_A
timestamp 1751532392
transform -1 0 21728 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input3_A
timestamp 1751532392
transform -1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input4_A
timestamp 1751532392
transform -1 0 21728 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input5_A
timestamp 1751532392
transform -1 0 21728 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input6_A
timestamp 1751532392
transform -1 0 21728 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532351
transform 1 0 1568 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_18
timestamp 1751532351
transform 1 0 3360 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_36
timestamp 1751532351
transform 1 0 5376 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_52
timestamp 1751532351
transform 1 0 7168 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_70
timestamp 1751532351
transform 1 0 9184 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_86
timestamp 1751532351
transform 1 0 10976 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_104
timestamp 1751532351
transform 1 0 12992 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_120
timestamp 1751532351
transform 1 0 14784 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_138
timestamp 1751532351
transform 1 0 16800 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_154
timestamp 1751532351
transform 1 0 18592 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_172
timestamp 1751532351
transform 1 0 20608 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532312
transform 1 0 1568 0 -1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_10 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532246
transform 1 0 2464 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_28 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532440
transform 1 0 4480 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_32
timestamp 1751532351
transform 1 0 4928 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_48
timestamp 1751532246
transform 1 0 6720 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_52
timestamp 1751532440
transform 1 0 7168 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_54 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532423
transform 1 0 7392 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_61
timestamp 1751532246
transform 1 0 8176 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_67
timestamp 1751532440
transform 1 0 8848 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_69
timestamp 1751532423
transform 1 0 9072 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_72
timestamp 1751532351
transform 1 0 9408 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_88
timestamp 1751532440
transform 1 0 11200 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_90
timestamp 1751532423
transform 1 0 11424 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_103
timestamp 1751532246
transform 1 0 12880 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_107
timestamp 1751532440
transform 1 0 13328 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_111
timestamp 1751532423
transform 1 0 13776 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_118
timestamp 1751532351
transform 1 0 14560 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_134
timestamp 1751532246
transform 1 0 16352 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_138
timestamp 1751532440
transform 1 0 16800 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_1_146
timestamp 1751532312
transform 1 0 17696 0 -1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_154
timestamp 1751532246
transform 1 0 18592 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_158
timestamp 1751532423
transform 1 0 19040 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_179
timestamp 1751532440
transform 1 0 21392 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_183
timestamp 1751532440
transform 1 0 21840 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_187
timestamp 1751532423
transform 1 0 22288 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_2
timestamp 1751532351
transform 1 0 1568 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_32
timestamp 1751532440
transform 1 0 4928 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_34
timestamp 1751532423
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_2_37
timestamp 1751532312
transform 1 0 5488 0 1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_71
timestamp 1751532440
transform 1 0 9296 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_2_75
timestamp 1751532246
transform 1 0 9744 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_79
timestamp 1751532440
transform 1 0 10192 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_81
timestamp 1751532423
transform 1 0 10416 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_103
timestamp 1751532440
transform 1 0 12880 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_118
timestamp 1751532440
transform 1 0 14560 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_120
timestamp 1751532423
transform 1 0 14784 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_2_132
timestamp 1751532246
transform 1 0 16128 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_136
timestamp 1751532440
transform 1 0 16576 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_144
timestamp 1751532423
transform 1 0 17472 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_166
timestamp 1751532440
transform 1 0 19936 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_168
timestamp 1751532423
transform 1 0 20160 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_177
timestamp 1751532440
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_179
timestamp 1751532423
transform 1 0 21392 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_2
timestamp 1751532351
transform 1 0 1568 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_3_32
timestamp 1751532312
transform 1 0 4928 0 -1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_40
timestamp 1751532440
transform 1 0 5824 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_42
timestamp 1751532423
transform 1 0 6048 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_53
timestamp 1751532440
transform 1 0 7280 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_55
timestamp 1751532423
transform 1 0 7504 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_66
timestamp 1751532246
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_3_72
timestamp 1751532312
transform 1 0 9408 0 -1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_80
timestamp 1751532246
transform 1 0 10304 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_84
timestamp 1751532440
transform 1 0 10752 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_86
timestamp 1751532423
transform 1 0 10976 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_3_98
timestamp 1751532312
transform 1 0 12320 0 -1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_106
timestamp 1751532246
transform 1 0 13216 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_110
timestamp 1751532440
transform 1 0 13664 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_112
timestamp 1751532423
transform 1 0 13888 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_3_126
timestamp 1751532312
transform 1 0 15456 0 -1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_134
timestamp 1751532246
transform 1 0 16352 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_138
timestamp 1751532440
transform 1 0 16800 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_142
timestamp 1751532351
transform 1 0 17248 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_158
timestamp 1751532440
transform 1 0 19040 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_3_173
timestamp 1751532312
transform 1 0 20720 0 -1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_181
timestamp 1751532246
transform 1 0 21616 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_185
timestamp 1751532440
transform 1 0 22064 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_187
timestamp 1751532423
transform 1 0 22288 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_2
timestamp 1751532351
transform 1 0 1568 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_18
timestamp 1751532351
transform 1 0 3360 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_34
timestamp 1751532423
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_37
timestamp 1751532351
transform 1 0 5488 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_53
timestamp 1751532440
transform 1 0 7280 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_65
timestamp 1751532351
transform 1 0 8624 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_81
timestamp 1751532351
transform 1 0 10416 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_4_97
timestamp 1751532312
transform 1 0 12208 0 1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_107
timestamp 1751532351
transform 1 0 13328 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_123
timestamp 1751532351
transform 1 0 15120 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_139
timestamp 1751532351
transform 1 0 16912 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_155
timestamp 1751532351
transform 1 0 18704 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_4_171
timestamp 1751532246
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_4_177
timestamp 1751532312
transform 1 0 21168 0 1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_185
timestamp 1751532440
transform 1 0 22064 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_187
timestamp 1751532423
transform 1 0 22288 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_5_2
timestamp 1751532312
transform 1 0 1568 0 -1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_10
timestamp 1751532246
transform 1 0 2464 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_14
timestamp 1751532440
transform 1 0 2912 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_32
timestamp 1751532440
transform 1 0 4928 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_36
timestamp 1751532351
transform 1 0 5376 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_52
timestamp 1751532351
transform 1 0 7168 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_68
timestamp 1751532440
transform 1 0 8960 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_72
timestamp 1751532351
transform 1 0 9408 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_88
timestamp 1751532351
transform 1 0 11200 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_104
timestamp 1751532351
transform 1 0 12992 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_120
timestamp 1751532351
transform 1 0 14784 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_136
timestamp 1751532246
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_142
timestamp 1751532246
transform 1 0 17248 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_5_154
timestamp 1751532312
transform 1 0 18592 0 -1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_162
timestamp 1751532246
transform 1 0 19488 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_166
timestamp 1751532440
transform 1 0 19936 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_5_178
timestamp 1751532312
transform 1 0 21280 0 -1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_186
timestamp 1751532440
transform 1 0 22176 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_6_2
timestamp 1751532312
transform 1 0 1568 0 1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_10
timestamp 1751532246
transform 1 0 2464 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_14
timestamp 1751532440
transform 1 0 2912 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_20
timestamp 1751532423
transform 1 0 3584 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_31
timestamp 1751532440
transform 1 0 4816 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_37
timestamp 1751532440
transform 1 0 5488 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_41
timestamp 1751532351
transform 1 0 5936 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_57
timestamp 1751532440
transform 1 0 7728 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_65
timestamp 1751532440
transform 1 0 8624 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_67
timestamp 1751532423
transform 1 0 8848 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_78
timestamp 1751532351
transform 1 0 10080 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_6_94
timestamp 1751532312
transform 1 0 11872 0 1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_102
timestamp 1751532440
transform 1 0 12768 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_104
timestamp 1751532423
transform 1 0 12992 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_114
timestamp 1751532351
transform 1 0 14112 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_6_130
timestamp 1751532312
transform 1 0 15904 0 1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_138
timestamp 1751532246
transform 1 0 16800 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_6_162
timestamp 1751532312
transform 1 0 19488 0 1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_170
timestamp 1751532246
transform 1 0 20384 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_174
timestamp 1751532423
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_177
timestamp 1751532440
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_179
timestamp 1751532423
transform 1 0 21392 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_2
timestamp 1751532351
transform 1 0 1568 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_7_18
timestamp 1751532312
transform 1 0 3360 0 -1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_26
timestamp 1751532440
transform 1 0 4256 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_28
timestamp 1751532423
transform 1 0 4480 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_36
timestamp 1751532440
transform 1 0 5376 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_7_40
timestamp 1751532312
transform 1 0 5824 0 -1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_48
timestamp 1751532246
transform 1 0 6720 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_52
timestamp 1751532423
transform 1 0 7168 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_91
timestamp 1751532246
transform 1 0 11536 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_95
timestamp 1751532423
transform 1 0 11984 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_106
timestamp 1751532423
transform 1 0 13216 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_7_128
timestamp 1751532312
transform 1 0 15680 0 -1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_136
timestamp 1751532246
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_142
timestamp 1751532440
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_144
timestamp 1751532423
transform 1 0 17472 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_166
timestamp 1751532440
transform 1 0 19936 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_168
timestamp 1751532423
transform 1 0 20160 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_7_175
timestamp 1751532312
transform 1 0 20944 0 -1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_183
timestamp 1751532246
transform 1 0 21840 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_187
timestamp 1751532423
transform 1 0 22288 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_2
timestamp 1751532351
transform 1 0 1568 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_18
timestamp 1751532246
transform 1 0 3360 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_22
timestamp 1751532440
transform 1 0 3808 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_24
timestamp 1751532423
transform 1 0 4032 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_47
timestamp 1751532440
transform 1 0 6608 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_8_51
timestamp 1751532312
transform 1 0 7056 0 1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_59
timestamp 1751532440
transform 1 0 7952 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_75
timestamp 1751532351
transform 1 0 9744 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_8_91
timestamp 1751532312
transform 1 0 11536 0 1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_99
timestamp 1751532246
transform 1 0 12432 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_103
timestamp 1751532440
transform 1 0 12880 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_107
timestamp 1751532423
transform 1 0 13328 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_115
timestamp 1751532351
transform 1 0 14224 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_131
timestamp 1751532351
transform 1 0 16016 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_153
timestamp 1751532440
transform 1 0 18480 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_159
timestamp 1751532440
transform 1 0 19152 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_163
timestamp 1751532246
transform 1 0 19600 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_167
timestamp 1751532440
transform 1 0 20048 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_187
timestamp 1751532423
transform 1 0 22288 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_9_2
timestamp 1751532312
transform 1 0 1568 0 -1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_10
timestamp 1751532246
transform 1 0 2464 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_14
timestamp 1751532440
transform 1 0 2912 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_26
timestamp 1751532351
transform 1 0 4256 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_42
timestamp 1751532351
transform 1 0 6048 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_9_58
timestamp 1751532312
transform 1 0 7840 0 -1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_66
timestamp 1751532246
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_72
timestamp 1751532351
transform 1 0 9408 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_88
timestamp 1751532351
transform 1 0 11200 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_104
timestamp 1751532351
transform 1 0 12992 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_120
timestamp 1751532351
transform 1 0 14784 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_136
timestamp 1751532246
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_142
timestamp 1751532246
transform 1 0 17248 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_152
timestamp 1751532351
transform 1 0 18368 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_9_168
timestamp 1751532312
transform 1 0 20160 0 -1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_176
timestamp 1751532246
transform 1 0 21056 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_10_2
timestamp 1751532312
transform 1 0 1568 0 1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_10
timestamp 1751532440
transform 1 0 2464 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_37
timestamp 1751532351
transform 1 0 5488 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_53
timestamp 1751532351
transform 1 0 7280 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_69
timestamp 1751532351
transform 1 0 9072 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_85
timestamp 1751532351
transform 1 0 10864 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_101
timestamp 1751532246
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_107
timestamp 1751532351
transform 1 0 13328 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_123
timestamp 1751532351
transform 1 0 15120 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_10_139
timestamp 1751532312
transform 1 0 16912 0 1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_147
timestamp 1751532246
transform 1 0 17808 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_151
timestamp 1751532440
transform 1 0 18256 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_153
timestamp 1751532423
transform 1 0 18480 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_10_161
timestamp 1751532312
transform 1 0 19376 0 1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_169
timestamp 1751532246
transform 1 0 20272 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_173
timestamp 1751532440
transform 1 0 20720 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_10_177
timestamp 1751532312
transform 1 0 21168 0 1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_185
timestamp 1751532440
transform 1 0 22064 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_187
timestamp 1751532423
transform 1 0 22288 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_11_2
timestamp 1751532312
transform 1 0 1568 0 -1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_10
timestamp 1751532246
transform 1 0 2464 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_14
timestamp 1751532440
transform 1 0 2912 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_22
timestamp 1751532351
transform 1 0 3808 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_38
timestamp 1751532351
transform 1 0 5600 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_11_54
timestamp 1751532312
transform 1 0 7392 0 -1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_62
timestamp 1751532423
transform 1 0 8288 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_82
timestamp 1751532246
transform 1 0 10528 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_86
timestamp 1751532440
transform 1 0 10976 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_88
timestamp 1751532423
transform 1 0 11200 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_102
timestamp 1751532440
transform 1 0 12768 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_104
timestamp 1751532423
transform 1 0 12992 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_116
timestamp 1751532246
transform 1 0 14336 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_120
timestamp 1751532440
transform 1 0 14784 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_122
timestamp 1751532423
transform 1 0 15008 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_11_127
timestamp 1751532312
transform 1 0 15568 0 -1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_135
timestamp 1751532246
transform 1 0 16464 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_139
timestamp 1751532423
transform 1 0 16912 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_142
timestamp 1751532440
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_171
timestamp 1751532351
transform 1 0 20496 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_187
timestamp 1751532423
transform 1 0 22288 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_12_2
timestamp 1751532351
transform 1 0 1568 0 1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_18
timestamp 1751532312
transform 1 0 3360 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_26
timestamp 1751532440
transform 1 0 4256 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_28
timestamp 1751532423
transform 1 0 4480 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_12_37
timestamp 1751532351
transform 1 0 5488 0 1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_60
timestamp 1751532440
transform 1 0 8064 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_12_69
timestamp 1751532351
transform 1 0 9072 0 1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_85
timestamp 1751532312
transform 1 0 10864 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_100
timestamp 1751532246
transform 1 0 12544 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_104
timestamp 1751532423
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_121
timestamp 1751532312
transform 1 0 14896 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_129
timestamp 1751532246
transform 1 0 15792 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_12_151
timestamp 1751532351
transform 1 0 18256 0 1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_167
timestamp 1751532246
transform 1 0 20048 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_171
timestamp 1751532440
transform 1 0 20496 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_177
timestamp 1751532440
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_181
timestamp 1751532423
transform 1 0 21616 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_2
timestamp 1751532351
transform 1 0 1568 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_18
timestamp 1751532246
transform 1 0 3360 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_22
timestamp 1751532423
transform 1 0 3808 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_36
timestamp 1751532440
transform 1 0 5376 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_13_40
timestamp 1751532312
transform 1 0 5824 0 -1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_48
timestamp 1751532246
transform 1 0 6720 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_13_78
timestamp 1751532312
transform 1 0 10080 0 -1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_86
timestamp 1751532246
transform 1 0 10976 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_101
timestamp 1751532246
transform 1 0 12656 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_105
timestamp 1751532440
transform 1 0 13104 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_114
timestamp 1751532351
transform 1 0 14112 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_13_130
timestamp 1751532312
transform 1 0 15904 0 -1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_138
timestamp 1751532440
transform 1 0 16800 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_13_148
timestamp 1751532312
transform 1 0 17920 0 -1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_156
timestamp 1751532246
transform 1 0 18816 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_160
timestamp 1751532440
transform 1 0 19264 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_162
timestamp 1751532423
transform 1 0 19488 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_184
timestamp 1751532246
transform 1 0 21952 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_2
timestamp 1751532351
transform 1 0 1568 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_14_18
timestamp 1751532312
transform 1 0 3360 0 1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_26
timestamp 1751532440
transform 1 0 4256 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_37
timestamp 1751532440
transform 1 0 5488 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_41
timestamp 1751532351
transform 1 0 5936 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_57
timestamp 1751532440
transform 1 0 7728 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_59
timestamp 1751532423
transform 1 0 7952 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_66
timestamp 1751532351
transform 1 0 8736 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_82
timestamp 1751532351
transform 1 0 10528 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_98
timestamp 1751532246
transform 1 0 12320 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_102
timestamp 1751532440
transform 1 0 12768 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_104
timestamp 1751532423
transform 1 0 12992 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_114
timestamp 1751532351
transform 1 0 14112 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_130
timestamp 1751532351
transform 1 0 15904 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_146
timestamp 1751532351
transform 1 0 17696 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_14_162
timestamp 1751532312
transform 1 0 19488 0 1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_170
timestamp 1751532246
transform 1 0 20384 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_174
timestamp 1751532423
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_183
timestamp 1751532246
transform 1 0 21840 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_187
timestamp 1751532423
transform 1 0 22288 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_2
timestamp 1751532351
transform 1 0 1568 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_25
timestamp 1751532351
transform 1 0 4144 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_41
timestamp 1751532351
transform 1 0 5936 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_15_57
timestamp 1751532312
transform 1 0 7728 0 -1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_65
timestamp 1751532246
transform 1 0 8624 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_69
timestamp 1751532423
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_72
timestamp 1751532351
transform 1 0 9408 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_88
timestamp 1751532246
transform 1 0 11200 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_92
timestamp 1751532440
transform 1 0 11648 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_94
timestamp 1751532423
transform 1 0 11872 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_15_106
timestamp 1751532312
transform 1 0 13216 0 -1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_114
timestamp 1751532246
transform 1 0 14112 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_118
timestamp 1751532423
transform 1 0 14560 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_15_126
timestamp 1751532312
transform 1 0 15456 0 -1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_134
timestamp 1751532246
transform 1 0 16352 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_138
timestamp 1751532440
transform 1 0 16800 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_142
timestamp 1751532246
transform 1 0 17248 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_146
timestamp 1751532440
transform 1 0 17696 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_148
timestamp 1751532423
transform 1 0 17920 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_156
timestamp 1751532423
transform 1 0 18816 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_164
timestamp 1751532246
transform 1 0 19712 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_15_179
timestamp 1751532312
transform 1 0 21392 0 -1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_187
timestamp 1751532423
transform 1 0 22288 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_2
timestamp 1751532312
transform 1 0 1568 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_10
timestamp 1751532246
transform 1 0 2464 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_14
timestamp 1751532423
transform 1 0 2912 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_32
timestamp 1751532440
transform 1 0 4928 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_34
timestamp 1751532423
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_37
timestamp 1751532351
transform 1 0 5488 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_53
timestamp 1751532351
transform 1 0 7280 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_69
timestamp 1751532351
transform 1 0 9072 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_85
timestamp 1751532246
transform 1 0 10864 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_89
timestamp 1751532440
transform 1 0 11312 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_93
timestamp 1751532312
transform 1 0 11760 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_101
timestamp 1751532246
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_107
timestamp 1751532246
transform 1 0 13328 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_111
timestamp 1751532440
transform 1 0 13776 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_113
timestamp 1751532423
transform 1 0 14000 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_131
timestamp 1751532351
transform 1 0 16016 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_147
timestamp 1751532440
transform 1 0 17808 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_163
timestamp 1751532312
transform 1 0 19600 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_171
timestamp 1751532246
transform 1 0 20496 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_177
timestamp 1751532312
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_185
timestamp 1751532440
transform 1 0 22064 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_187
timestamp 1751532423
transform 1 0 22288 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_17_2
timestamp 1751532312
transform 1 0 1568 0 -1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_10
timestamp 1751532423
transform 1 0 2464 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_34
timestamp 1751532351
transform 1 0 5152 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_50
timestamp 1751532246
transform 1 0 6944 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_61
timestamp 1751532440
transform 1 0 8176 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_65
timestamp 1751532246
transform 1 0 8624 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_69
timestamp 1751532423
transform 1 0 9072 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_17_72
timestamp 1751532312
transform 1 0 9408 0 -1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_80
timestamp 1751532440
transform 1 0 10304 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_82
timestamp 1751532423
transform 1 0 10528 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_90
timestamp 1751532440
transform 1 0 11424 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_92
timestamp 1751532423
transform 1 0 11648 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_107
timestamp 1751532351
transform 1 0 13328 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_123
timestamp 1751532351
transform 1 0 15120 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_139
timestamp 1751532423
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_17_142
timestamp 1751532312
transform 1 0 17248 0 -1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_150
timestamp 1751532423
transform 1 0 18144 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_157
timestamp 1751532351
transform 1 0 18928 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_173
timestamp 1751532246
transform 1 0 20720 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_177
timestamp 1751532440
transform 1 0 21168 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_179
timestamp 1751532423
transform 1 0 21392 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_18_2
timestamp 1751532312
transform 1 0 1568 0 1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_10
timestamp 1751532423
transform 1 0 2464 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_31
timestamp 1751532246
transform 1 0 4816 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_37
timestamp 1751532351
transform 1 0 5488 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_53
timestamp 1751532246
transform 1 0 7280 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_57
timestamp 1751532440
transform 1 0 7728 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_59
timestamp 1751532423
transform 1 0 7952 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_74
timestamp 1751532351
transform 1 0 9632 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_18_92
timestamp 1751532312
transform 1 0 11648 0 1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_100
timestamp 1751532440
transform 1 0 12544 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_102
timestamp 1751532423
transform 1 0 12768 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_121
timestamp 1751532351
transform 1 0 14896 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_137
timestamp 1751532351
transform 1 0 16688 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_153
timestamp 1751532351
transform 1 0 18480 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_169
timestamp 1751532246
transform 1 0 20272 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_173
timestamp 1751532440
transform 1 0 20720 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_18_177
timestamp 1751532312
transform 1 0 21168 0 1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_185
timestamp 1751532440
transform 1 0 22064 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_187
timestamp 1751532423
transform 1 0 22288 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_19_2
timestamp 1751532351
transform 1 0 1568 0 -1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_18
timestamp 1751532423
transform 1 0 3360 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_19_21
timestamp 1751532351
transform 1 0 3696 0 -1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_19_37
timestamp 1751532312
transform 1 0 5488 0 -1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_45
timestamp 1751532246
transform 1 0 6384 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_49
timestamp 1751532440
transform 1 0 6832 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_51
timestamp 1751532423
transform 1 0 7056 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_79
timestamp 1751532246
transform 1 0 10192 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_19_89
timestamp 1751532351
transform 1 0 11312 0 -1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_105
timestamp 1751532246
transform 1 0 13104 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_109
timestamp 1751532440
transform 1 0 13552 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_111
timestamp 1751532423
transform 1 0 13776 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_19_125
timestamp 1751532312
transform 1 0 15344 0 -1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_133
timestamp 1751532246
transform 1 0 16240 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_137
timestamp 1751532440
transform 1 0 16688 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_139
timestamp 1751532423
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_142
timestamp 1751532246
transform 1 0 17248 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_146
timestamp 1751532423
transform 1 0 17696 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_153
timestamp 1751532440
transform 1 0 18480 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_161
timestamp 1751532440
transform 1 0 19376 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_177
timestamp 1751532440
transform 1 0 21168 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_179
timestamp 1751532423
transform 1 0 21392 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_20_2
timestamp 1751532312
transform 1 0 1568 0 1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_10
timestamp 1751532440
transform 1 0 2464 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_12
timestamp 1751532423
transform 1 0 2688 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_20_43
timestamp 1751532312
transform 1 0 6160 0 1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_51
timestamp 1751532246
transform 1 0 7056 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_55
timestamp 1751532440
transform 1 0 7504 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_57
timestamp 1751532423
transform 1 0 7728 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_68
timestamp 1751532423
transform 1 0 8960 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_20_75
timestamp 1751532312
transform 1 0 9744 0 1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_20_89
timestamp 1751532351
transform 1 0 11312 0 1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_107
timestamp 1751532246
transform 1 0 13328 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_111
timestamp 1751532440
transform 1 0 13776 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_126
timestamp 1751532440
transform 1 0 15456 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_130
timestamp 1751532423
transform 1 0 15904 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_20_137
timestamp 1751532312
transform 1 0 16688 0 1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_145
timestamp 1751532246
transform 1 0 17584 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_149
timestamp 1751532440
transform 1 0 18032 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_173
timestamp 1751532440
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_183
timestamp 1751532246
transform 1 0 21840 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_187
timestamp 1751532423
transform 1 0 22288 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_2
timestamp 1751532440
transform 1 0 1568 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_4
timestamp 1751532423
transform 1 0 1792 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_11
timestamp 1751532312
transform 1 0 2576 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_19
timestamp 1751532246
transform 1 0 3472 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_23
timestamp 1751532440
transform 1 0 3920 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_31
timestamp 1751532440
transform 1 0 4816 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_33
timestamp 1751532423
transform 1 0 5040 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_36
timestamp 1751532312
transform 1 0 5376 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_44
timestamp 1751532423
transform 1 0 6272 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_51
timestamp 1751532351
transform 1 0 7056 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_67
timestamp 1751532423
transform 1 0 8848 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_76
timestamp 1751532312
transform 1 0 9856 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_84
timestamp 1751532423
transform 1 0 10752 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_91
timestamp 1751532312
transform 1 0 11536 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_99
timestamp 1751532440
transform 1 0 12432 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_101
timestamp 1751532423
transform 1 0 12656 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_104
timestamp 1751532423
transform 1 0 12992 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_111
timestamp 1751532312
transform 1 0 13776 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_119
timestamp 1751532246
transform 1 0 14672 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_123
timestamp 1751532440
transform 1 0 15120 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_131
timestamp 1751532246
transform 1 0 16016 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_135
timestamp 1751532423
transform 1 0 16464 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_138
timestamp 1751532246
transform 1 0 16800 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_142
timestamp 1751532440
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_144
timestamp 1751532423
transform 1 0 17472 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_151
timestamp 1751532312
transform 1 0 18256 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_159
timestamp 1751532246
transform 1 0 19152 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_163
timestamp 1751532423
transform 1 0 19600 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_178
timestamp 1751532246
transform 1 0 21280 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input1
timestamp 1751534193
transform -1 0 22400 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input2
timestamp 1751534193
transform -1 0 22400 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input3
timestamp 1751534193
transform -1 0 22400 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input4
timestamp 1751534193
transform -1 0 22400 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input5
timestamp 1751534193
transform -1 0 22400 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input6
timestamp 1751534193
transform -1 0 22400 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  output7
timestamp 1751534193
transform 1 0 19712 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  output8
timestamp 1751534193
transform -1 0 2576 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  output9
timestamp 1751534193
transform 1 0 4144 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  output10
timestamp 1751534193
transform 1 0 6384 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  output11
timestamp 1751534193
transform 1 0 9184 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  output12
timestamp 1751534193
transform 1 0 10864 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  output13
timestamp 1751534193
transform -1 0 13776 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  output14
timestamp 1751534193
transform 1 0 15344 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  output15
timestamp 1751534193
transform 1 0 17584 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  output16
timestamp 1751534193
transform 1 0 20608 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  output17
timestamp 1751534193
transform 1 0 21728 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_0_Left_22 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532504
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_0_Right_0
timestamp 1751532504
transform -1 0 22624 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_1_Left_23
timestamp 1751532504
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_1_Right_1
timestamp 1751532504
transform -1 0 22624 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_2_Left_24
timestamp 1751532504
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_2_Right_2
timestamp 1751532504
transform -1 0 22624 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_3_Left_25
timestamp 1751532504
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_3_Right_3
timestamp 1751532504
transform -1 0 22624 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_4_Left_26
timestamp 1751532504
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_4_Right_4
timestamp 1751532504
transform -1 0 22624 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_5_Left_27
timestamp 1751532504
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_5_Right_5
timestamp 1751532504
transform -1 0 22624 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_6_Left_28
timestamp 1751532504
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_6_Right_6
timestamp 1751532504
transform -1 0 22624 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_7_Left_29
timestamp 1751532504
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_7_Right_7
timestamp 1751532504
transform -1 0 22624 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_8_Left_30
timestamp 1751532504
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_8_Right_8
timestamp 1751532504
transform -1 0 22624 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_9_Left_31
timestamp 1751532504
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_9_Right_9
timestamp 1751532504
transform -1 0 22624 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_10_Left_32
timestamp 1751532504
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_10_Right_10
timestamp 1751532504
transform -1 0 22624 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_11_Left_33
timestamp 1751532504
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_11_Right_11
timestamp 1751532504
transform -1 0 22624 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_12_Left_34
timestamp 1751532504
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_12_Right_12
timestamp 1751532504
transform -1 0 22624 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_13_Left_35
timestamp 1751532504
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_13_Right_13
timestamp 1751532504
transform -1 0 22624 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_14_Left_36
timestamp 1751532504
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_14_Right_14
timestamp 1751532504
transform -1 0 22624 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_15_Left_37
timestamp 1751532504
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_15_Right_15
timestamp 1751532504
transform -1 0 22624 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_16_Left_38
timestamp 1751532504
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_16_Right_16
timestamp 1751532504
transform -1 0 22624 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_17_Left_39
timestamp 1751532504
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_17_Right_17
timestamp 1751532504
transform -1 0 22624 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_18_Left_40
timestamp 1751532504
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_18_Right_18
timestamp 1751532504
transform -1 0 22624 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_19_Left_41
timestamp 1751532504
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_19_Right_19
timestamp 1751532504
transform -1 0 22624 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_20_Left_42
timestamp 1751532504
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_20_Right_20
timestamp 1751532504
transform -1 0 22624 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_21_Left_43
timestamp 1751532504
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_21_Right_21
timestamp 1751532504
transform -1 0 22624 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_44
timestamp 1751532504
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_45
timestamp 1751532504
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_46
timestamp 1751532504
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_47
timestamp 1751532504
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_48
timestamp 1751532504
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_49
timestamp 1751532504
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_50
timestamp 1751532504
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_51
timestamp 1751532504
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_52
timestamp 1751532504
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_53
timestamp 1751532504
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_54
timestamp 1751532504
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_55
timestamp 1751532504
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_56
timestamp 1751532504
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_57
timestamp 1751532504
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_58
timestamp 1751532504
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_59
timestamp 1751532504
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_60
timestamp 1751532504
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_61
timestamp 1751532504
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_62
timestamp 1751532504
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_63
timestamp 1751532504
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_64
timestamp 1751532504
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_65
timestamp 1751532504
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_66
timestamp 1751532504
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_67
timestamp 1751532504
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_68
timestamp 1751532504
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_69
timestamp 1751532504
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_70
timestamp 1751532504
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_71
timestamp 1751532504
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_72
timestamp 1751532504
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_73
timestamp 1751532504
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_74
timestamp 1751532504
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_75
timestamp 1751532504
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_76
timestamp 1751532504
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_77
timestamp 1751532504
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_78
timestamp 1751532504
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_79
timestamp 1751532504
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_80
timestamp 1751532504
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_81
timestamp 1751532504
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_82
timestamp 1751532504
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_83
timestamp 1751532504
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_84
timestamp 1751532504
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_85
timestamp 1751532504
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_86
timestamp 1751532504
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_87
timestamp 1751532504
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_88
timestamp 1751532504
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_89
timestamp 1751532504
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_90
timestamp 1751532504
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_91
timestamp 1751532504
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_92
timestamp 1751532504
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_93
timestamp 1751532504
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_94
timestamp 1751532504
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_95
timestamp 1751532504
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_96
timestamp 1751532504
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_97
timestamp 1751532504
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_98
timestamp 1751532504
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_99
timestamp 1751532504
transform 1 0 5152 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_100
timestamp 1751532504
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_101
timestamp 1751532504
transform 1 0 12768 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_102
timestamp 1751532504
transform 1 0 16576 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_103
timestamp 1751532504
transform 1 0 20384 0 -1 20384
box -86 -86 310 870
<< labels >>
flabel metal3 s 23200 1568 24000 1680 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 23200 7392 24000 7504 0 FreeSans 448 0 0 0 io_in[0]
port 1 nsew signal input
flabel metal3 s 23200 10304 24000 10416 0 FreeSans 448 0 0 0 io_in[1]
port 2 nsew signal input
flabel metal3 s 23200 13216 24000 13328 0 FreeSans 448 0 0 0 io_in[2]
port 3 nsew signal input
flabel metal3 s 23200 16128 24000 16240 0 FreeSans 448 0 0 0 io_in[3]
port 4 nsew signal input
flabel metal3 s 23200 19040 24000 19152 0 FreeSans 448 0 0 0 io_in[4]
port 5 nsew signal input
flabel metal3 s 23200 21952 24000 22064 0 FreeSans 448 0 0 0 io_oeb
port 6 nsew signal output
flabel metal2 s 1792 23200 1904 24000 0 FreeSans 448 90 0 0 io_out[0]
port 7 nsew signal output
flabel metal2 s 4032 23200 4144 24000 0 FreeSans 448 90 0 0 io_out[1]
port 8 nsew signal output
flabel metal2 s 6272 23200 6384 24000 0 FreeSans 448 90 0 0 io_out[2]
port 9 nsew signal output
flabel metal2 s 8512 23200 8624 24000 0 FreeSans 448 90 0 0 io_out[3]
port 10 nsew signal output
flabel metal2 s 10752 23200 10864 24000 0 FreeSans 448 90 0 0 io_out[4]
port 11 nsew signal output
flabel metal2 s 12992 23200 13104 24000 0 FreeSans 448 90 0 0 io_out[5]
port 12 nsew signal output
flabel metal2 s 15232 23200 15344 24000 0 FreeSans 448 90 0 0 io_out[6]
port 13 nsew signal output
flabel metal2 s 17472 23200 17584 24000 0 FreeSans 448 90 0 0 io_out[7]
port 14 nsew signal output
flabel metal2 s 19712 23200 19824 24000 0 FreeSans 448 90 0 0 io_out[8]
port 15 nsew signal output
flabel metal2 s 21952 23200 22064 24000 0 FreeSans 448 90 0 0 io_out[9]
port 16 nsew signal output
flabel metal3 s 23200 4480 24000 4592 0 FreeSans 448 0 0 0 rst_n
port 17 nsew signal input
flabel metal4 s 3844 3076 4164 20444 0 FreeSans 1280 90 0 0 vdd
port 18 nsew power bidirectional
flabel metal4 s 9164 3076 9484 20444 0 FreeSans 1280 90 0 0 vdd
port 18 nsew power bidirectional
flabel metal4 s 14484 3076 14804 20444 0 FreeSans 1280 90 0 0 vdd
port 18 nsew power bidirectional
flabel metal4 s 19804 3076 20124 20444 0 FreeSans 1280 90 0 0 vdd
port 18 nsew power bidirectional
flabel metal4 s 6504 3076 6824 20444 0 FreeSans 1280 90 0 0 vss
port 19 nsew ground bidirectional
flabel metal4 s 11824 3076 12144 20444 0 FreeSans 1280 90 0 0 vss
port 19 nsew ground bidirectional
flabel metal4 s 17144 3076 17464 20444 0 FreeSans 1280 90 0 0 vss
port 19 nsew ground bidirectional
flabel metal4 s 22464 3076 22784 20444 0 FreeSans 1280 90 0 0 vss
port 19 nsew ground bidirectional
rlabel metal1 11984 19600 11984 19600 0 vdd
rlabel via1 12064 20384 12064 20384 0 vss
rlabel metal2 15624 5432 15624 5432 0 _000_
rlabel metal2 8232 6048 8232 6048 0 _001_
rlabel metal2 13188 17416 13188 17416 0 _002_
rlabel metal2 16856 5264 16856 5264 0 _003_
rlabel metal2 18536 5320 18536 5320 0 _004_
rlabel metal3 18480 5096 18480 5096 0 _005_
rlabel metal2 18648 5292 18648 5292 0 _006_
rlabel metal2 14504 4648 14504 4648 0 _007_
rlabel metal2 17192 13244 17192 13244 0 _008_
rlabel via2 12040 16872 12040 16872 0 _009_
rlabel metal2 8008 16912 8008 16912 0 _010_
rlabel metal3 12992 12152 12992 12152 0 _011_
rlabel metal2 14336 16296 14336 16296 0 _012_
rlabel metal2 12096 12936 12096 12936 0 _013_
rlabel metal2 12712 16172 12712 16172 0 _014_
rlabel metal2 14532 17864 14532 17864 0 _015_
rlabel metal2 14476 18536 14476 18536 0 _016_
rlabel metal2 18536 16184 18536 16184 0 _017_
rlabel metal2 18648 15232 18648 15232 0 _018_
rlabel metal2 10024 12880 10024 12880 0 _019_
rlabel metal2 7336 13664 7336 13664 0 _020_
rlabel metal2 5180 12936 5180 12936 0 _021_
rlabel metal2 20664 6776 20664 6776 0 _022_
rlabel metal2 20244 7896 20244 7896 0 _023_
rlabel metal2 20216 12230 20216 12230 0 _024_
rlabel metal2 18228 12152 18228 12152 0 _025_
rlabel metal2 12124 5656 12124 5656 0 _026_
rlabel metal2 17752 4984 17752 4984 0 _027_
rlabel metal2 17864 15568 17864 15568 0 _028_
rlabel metal2 9912 12488 9912 12488 0 _029_
rlabel metal2 4984 9492 4984 9492 0 _030_
rlabel metal2 3976 15680 3976 15680 0 _031_
rlabel metal2 3640 15764 3640 15764 0 _032_
rlabel metal2 3976 16744 3976 16744 0 _033_
rlabel metal2 3528 17780 3528 17780 0 _034_
rlabel via2 13832 9030 13832 9030 0 _035_
rlabel metal2 13091 16296 13091 16296 0 _036_
rlabel metal2 4872 17248 4872 17248 0 _037_
rlabel metal2 4704 9016 4704 9016 0 _038_
rlabel metal2 6104 9408 6104 9408 0 _039_
rlabel metal3 7000 7672 7000 7672 0 _040_
rlabel metal2 7784 7840 7784 7840 0 _041_
rlabel metal2 7896 8932 7896 8932 0 _042_
rlabel metal2 9464 8344 9464 8344 0 _043_
rlabel metal2 13052 9091 13052 9091 0 _044_
rlabel metal2 9576 8344 9576 8344 0 _045_
rlabel metal2 8456 8918 8456 8918 0 _046_
rlabel metal2 9072 8932 9072 8932 0 _047_
rlabel metal2 9016 8232 9016 8232 0 _048_
rlabel metal2 9800 8456 9800 8456 0 _049_
rlabel metal2 9520 9800 9520 9800 0 _050_
rlabel metal2 9576 9380 9576 9380 0 _051_
rlabel metal2 11032 6776 11032 6776 0 _052_
rlabel metal2 6552 5404 6552 5404 0 _053_
rlabel metal2 3304 5264 3304 5264 0 _054_
rlabel metal2 3640 6739 3640 6739 0 _055_
rlabel metal2 4302 4424 4302 4424 0 _056_
rlabel via2 6776 5082 6776 5082 0 _057_
rlabel metal2 11536 17248 11536 17248 0 _058_
rlabel metal2 8568 5600 8568 5600 0 _059_
rlabel metal2 7392 5404 7392 5404 0 _060_
rlabel metal3 8960 5096 8960 5096 0 _061_
rlabel metal2 18256 16576 18256 16576 0 _062_
rlabel metal2 19432 14455 19432 14455 0 _063_
rlabel metal2 18872 8176 18872 8176 0 _064_
rlabel metal2 18284 8344 18284 8344 0 _065_
rlabel metal3 20020 9016 20020 9016 0 _066_
rlabel metal3 18508 7672 18508 7672 0 _067_
rlabel metal3 18396 9576 18396 9576 0 _068_
rlabel metal3 16464 8344 16464 8344 0 _069_
rlabel metal2 19544 6608 19544 6608 0 _070_
rlabel metal2 19824 4312 19824 4312 0 _071_
rlabel metal2 3332 16856 3332 16856 0 _072_
rlabel metal2 13888 18032 13888 18032 0 _073_
rlabel metal2 9212 17640 9212 17640 0 _074_
rlabel metal2 8176 19208 8176 19208 0 _075_
rlabel metal2 7672 18095 7672 18095 0 _076_
rlabel metal2 5208 9044 5208 9044 0 _077_
rlabel metal2 4872 10640 4872 10640 0 _078_
rlabel metal2 2950 11872 2950 11872 0 _079_
rlabel metal2 4200 7616 4200 7616 0 _080_
rlabel metal2 3584 10612 3584 10612 0 _081_
rlabel metal2 4144 10780 4144 10780 0 _082_
rlabel metal3 20244 18424 20244 18424 0 _083_
rlabel metal2 20132 18536 20132 18536 0 _084_
rlabel metal2 20440 14588 20440 14588 0 _085_
rlabel metal2 20552 14196 20552 14196 0 _086_
rlabel metal2 10836 16968 10836 16968 0 _087_
rlabel metal2 20328 6160 20328 6160 0 _088_
rlabel metal2 15344 12488 15344 12488 0 _089_
rlabel metal2 8120 17248 8120 17248 0 _090_
rlabel metal2 8792 18368 8792 18368 0 _091_
rlabel metal2 8904 18900 8904 18900 0 _092_
rlabel metal2 15064 15988 15064 15988 0 _093_
rlabel metal2 20216 13272 20216 13272 0 _094_
rlabel metal2 19096 12320 19096 12320 0 _095_
rlabel metal3 18900 11592 18900 11592 0 _096_
rlabel metal2 19544 12208 19544 12208 0 _097_
rlabel metal2 8904 12264 8904 12264 0 _098_
rlabel metal2 8904 13804 8904 13804 0 _099_
rlabel metal2 15400 5824 15400 5824 0 _100_
rlabel metal3 16380 4536 16380 4536 0 _101_
rlabel metal2 22176 3920 22176 3920 0 clk
rlabel metal2 22344 7840 22344 7840 0 io_in[0]
rlabel metal2 22344 10472 22344 10472 0 io_in[1]
rlabel metal2 22344 13104 22344 13104 0 io_in[2]
rlabel metal2 22344 16520 22344 16520 0 io_in[3]
rlabel metal2 22344 18760 22344 18760 0 io_in[4]
rlabel metal3 21658 22008 21658 22008 0 io_oeb
rlabel metal2 1848 21686 1848 21686 0 io_out[0]
rlabel metal2 4088 21686 4088 21686 0 io_out[1]
rlabel metal2 6328 21686 6328 21686 0 io_out[2]
rlabel metal2 9240 23240 9240 23240 0 io_out[3]
rlabel metal2 10808 21686 10808 21686 0 io_out[4]
rlabel metal2 13048 21686 13048 21686 0 io_out[5]
rlabel metal2 15288 21686 15288 21686 0 io_out[6]
rlabel metal2 17528 21686 17528 21686 0 io_out[7]
rlabel metal2 19768 21686 19768 21686 0 io_out[8]
rlabel metal2 22064 20104 22064 20104 0 io_out[9]
rlabel metal2 3696 16296 3696 16296 0 main.CAR
rlabel metal2 3080 4592 3080 4592 0 main.GATES_1.input1
rlabel metal2 20888 9520 20888 9520 0 main.GATES_100.input1
rlabel metal2 19096 18816 19096 18816 0 main.GATES_100.input2
rlabel metal2 16856 12972 16856 12972 0 main.GATES_102.input1
rlabel metal2 15288 15568 15288 15568 0 main.GATES_102.input2
rlabel metal3 12040 13048 12040 13048 0 main.GATES_102.input3
rlabel metal2 3192 16268 3192 16268 0 main.GATES_103.input2
rlabel metal2 3864 15366 3864 15366 0 main.GATES_105.input3
rlabel metal2 8568 18760 8568 18760 0 main.GATES_106.input2
rlabel metal2 14784 15176 14784 15176 0 main.GATES_107.input2
rlabel metal2 11592 5208 11592 5208 0 main.GATES_108.input1
rlabel metal3 15064 18424 15064 18424 0 main.GATES_109.input1
rlabel metal2 9688 18375 9688 18375 0 main.GATES_109.input2
rlabel metal2 13608 10989 13608 10989 0 main.GATES_11.input2
rlabel metal2 4984 15904 4984 15904 0 main.GATES_110.input1
rlabel metal2 4536 18144 4536 18144 0 main.GATES_111.input2
rlabel metal3 12152 5096 12152 5096 0 main.GATES_113.input1
rlabel metal2 4256 9884 4256 9884 0 main.GATES_114.input2
rlabel metal3 16912 16072 16912 16072 0 main.GATES_115.input2
rlabel metal2 17640 13216 17640 13216 0 main.GATES_116.input1
rlabel metal2 8624 14504 8624 14504 0 main.GATES_116.input3
rlabel metal2 11200 5880 11200 5880 0 main.GATES_119.result
rlabel metal2 17864 4620 17864 4620 0 main.GATES_124.input2
rlabel metal2 17640 10640 17640 10640 0 main.GATES_125.input2
rlabel metal2 17752 11648 17752 11648 0 main.GATES_127.result
rlabel via2 4536 11354 4536 11354 0 main.GATES_132.input1
rlabel metal2 18872 11704 18872 11704 0 main.GATES_15.input3
rlabel metal2 20888 18704 20888 18704 0 main.GATES_16.input1
rlabel metal2 18648 7784 18648 7784 0 main.GATES_18.result
rlabel metal2 20552 15456 20552 15456 0 main.GATES_19.input1
rlabel metal2 14280 13384 14280 13384 0 main.GATES_20.result
rlabel metal2 19432 4816 19432 4816 0 main.GATES_26.input3
rlabel metal2 19208 15764 19208 15764 0 main.GATES_29.input3
rlabel metal2 18088 7784 18088 7784 0 main.GATES_46.input3
rlabel metal2 15064 18928 15064 18928 0 main.GATES_65.result
rlabel metal2 11032 18928 11032 18928 0 main.GATES_8.result
rlabel metal2 19320 18592 19320 18592 0 main.NOPF
rlabel metal3 4564 19208 4564 19208 0 main.WRITE
rlabel metal3 21084 8232 21084 8232 0 net1
rlabel metal3 5488 19432 5488 19432 0 net10
rlabel metal2 5880 19712 5880 19712 0 net11
rlabel metal2 10920 19712 10920 19712 0 net12
rlabel metal3 16352 18312 16352 18312 0 net13
rlabel metal2 15176 19712 15176 19712 0 net14
rlabel metal3 17024 19432 17024 19432 0 net15
rlabel metal2 20664 19712 20664 19712 0 net16
rlabel metal2 21672 19432 21672 19432 0 net17
rlabel metal2 22008 10080 22008 10080 0 net2
rlabel metal3 21840 13160 21840 13160 0 net3
rlabel metal2 21224 16072 21224 16072 0 net4
rlabel metal3 21616 8008 21616 8008 0 net5
rlabel metal2 20888 5432 20888 5432 0 net6
rlabel metal2 14280 19292 14280 19292 0 net7
rlabel metal2 3080 19712 3080 19712 0 net8
rlabel metal2 3752 19712 3752 19712 0 net9
rlabel metal2 22344 4816 22344 4816 0 rst_n
<< properties >>
string FIXED_BBOX 0 0 24000 24000
<< end >>
