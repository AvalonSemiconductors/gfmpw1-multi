magic
tech gf180mcuD
magscale 1 5
timestamp 1753967996
<< nwell >>
rect 629 9585 11355 10015
rect 629 8801 11355 9231
rect 629 8017 11355 8447
rect 629 7233 11355 7663
rect 629 6449 11355 6879
rect 629 5665 11355 6095
rect 629 4881 11355 5311
rect 629 4097 11355 4527
rect 629 3313 11355 3743
rect 629 2529 11355 2959
rect 629 1745 11355 2175
<< pwell >>
rect 629 10015 11355 10235
rect 629 9231 11355 9585
rect 629 8447 11355 8801
rect 629 7663 11355 8017
rect 629 6879 11355 7233
rect 629 6095 11355 6449
rect 629 5311 11355 5665
rect 629 4527 11355 4881
rect 629 3743 11355 4097
rect 629 2959 11355 3313
rect 629 2175 11355 2529
rect 629 1525 11355 1745
<< obsm1 >>
rect 672 1538 11392 10222
<< metal2 >>
rect 896 11600 952 12000
rect 2016 11600 2072 12000
rect 3136 11600 3192 12000
rect 4256 11600 4312 12000
rect 5376 11600 5432 12000
rect 6496 11600 6552 12000
rect 7616 11600 7672 12000
rect 8736 11600 8792 12000
rect 9856 11600 9912 12000
rect 10976 11600 11032 12000
<< obsm2 >>
rect 982 11570 1986 11634
rect 2102 11570 3106 11634
rect 3222 11570 4226 11634
rect 4342 11570 5346 11634
rect 5462 11570 6466 11634
rect 6582 11570 7586 11634
rect 7702 11570 8706 11634
rect 8822 11570 9826 11634
rect 9942 11570 10946 11634
rect 11062 11570 11378 11634
rect 910 793 11378 11570
<< metal3 >>
rect 11600 10976 12000 11032
rect 11600 9520 12000 9576
rect 11600 8064 12000 8120
rect 11600 6608 12000 6664
rect 11600 5152 12000 5208
rect 11600 3696 12000 3752
rect 11600 2240 12000 2296
rect 11600 784 12000 840
<< obsm3 >>
rect 1409 10946 11570 11018
rect 1409 9606 11600 10946
rect 1409 9490 11570 9606
rect 1409 8150 11600 9490
rect 1409 8034 11570 8150
rect 1409 6694 11600 8034
rect 1409 6578 11570 6694
rect 1409 5238 11600 6578
rect 1409 5122 11570 5238
rect 1409 3782 11600 5122
rect 1409 3666 11570 3782
rect 1409 2326 11600 3666
rect 1409 2210 11570 2326
rect 1409 870 11600 2210
rect 1409 798 11570 870
<< metal4 >>
rect 1922 1538 2082 10222
rect 3252 1538 3412 10222
rect 4582 1538 4742 10222
rect 5912 1538 6072 10222
rect 7242 1538 7402 10222
rect 8572 1538 8732 10222
rect 9902 1538 10062 10222
rect 11232 1538 11392 10222
<< obsm4 >>
rect 5166 6113 5194 6543
<< labels >>
rlabel metal3 s 11600 784 12000 840 6 clk
port 1 nsew signal input
rlabel metal3 s 11600 3696 12000 3752 6 io_in[0]
port 2 nsew signal input
rlabel metal3 s 11600 5152 12000 5208 6 io_in[1]
port 3 nsew signal input
rlabel metal3 s 11600 6608 12000 6664 6 io_in[2]
port 4 nsew signal input
rlabel metal3 s 11600 8064 12000 8120 6 io_in[3]
port 5 nsew signal input
rlabel metal3 s 11600 9520 12000 9576 6 io_in[4]
port 6 nsew signal input
rlabel metal3 s 11600 10976 12000 11032 6 io_oeb
port 7 nsew signal output
rlabel metal2 s 896 11600 952 12000 6 io_out[0]
port 8 nsew signal output
rlabel metal2 s 2016 11600 2072 12000 6 io_out[1]
port 9 nsew signal output
rlabel metal2 s 3136 11600 3192 12000 6 io_out[2]
port 10 nsew signal output
rlabel metal2 s 4256 11600 4312 12000 6 io_out[3]
port 11 nsew signal output
rlabel metal2 s 5376 11600 5432 12000 6 io_out[4]
port 12 nsew signal output
rlabel metal2 s 6496 11600 6552 12000 6 io_out[5]
port 13 nsew signal output
rlabel metal2 s 7616 11600 7672 12000 6 io_out[6]
port 14 nsew signal output
rlabel metal2 s 8736 11600 8792 12000 6 io_out[7]
port 15 nsew signal output
rlabel metal2 s 9856 11600 9912 12000 6 io_out[8]
port 16 nsew signal output
rlabel metal2 s 10976 11600 11032 12000 6 io_out[9]
port 17 nsew signal output
rlabel metal3 s 11600 2240 12000 2296 6 rst_n
port 18 nsew signal input
rlabel metal4 s 1922 1538 2082 10222 6 vdd
port 19 nsew power bidirectional
rlabel metal4 s 4582 1538 4742 10222 6 vdd
port 19 nsew power bidirectional
rlabel metal4 s 7242 1538 7402 10222 6 vdd
port 19 nsew power bidirectional
rlabel metal4 s 9902 1538 10062 10222 6 vdd
port 19 nsew power bidirectional
rlabel metal4 s 3252 1538 3412 10222 6 vss
port 20 nsew ground bidirectional
rlabel metal4 s 5912 1538 6072 10222 6 vss
port 20 nsew ground bidirectional
rlabel metal4 s 8572 1538 8732 10222 6 vss
port 20 nsew ground bidirectional
rlabel metal4 s 11232 1538 11392 10222 6 vss
port 20 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 12000 12000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 429652
string GDS_FILE /home/lucah/gfmpw1-multi/openlane/ue1/runs/25_07_31_15_19/results/signoff/ue1.magic.gds
string GDS_START 123196
<< end >>

