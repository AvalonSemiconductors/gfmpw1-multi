VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_sid
  CLASS BLOCK ;
  FOREIGN wrapped_sid ;
  ORIGIN 0.000 0.000 ;
  SIZE 1150.000 BY 800.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    ANTENNADIFFAREA 0.877000 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 13.440 1150.000 14.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 159.040 1150.000 159.600 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 173.600 1150.000 174.160 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 188.160 1150.000 188.720 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    ANTENNADIFFAREA 0.877000 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 202.720 1150.000 203.280 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 217.280 1150.000 217.840 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 231.840 1150.000 232.400 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 246.400 1150.000 246.960 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 260.960 1150.000 261.520 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 275.520 1150.000 276.080 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 290.080 1150.000 290.640 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    ANTENNADIFFAREA 0.877000 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 28.000 1150.000 28.560 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 304.640 1150.000 305.200 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 319.200 1150.000 319.760 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 333.760 1150.000 334.320 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 348.320 1150.000 348.880 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 362.880 1150.000 363.440 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 377.440 1150.000 378.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 392.000 1150.000 392.560 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 406.560 1150.000 407.120 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 421.120 1150.000 421.680 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 435.680 1150.000 436.240 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    ANTENNADIFFAREA 0.877000 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 42.560 1150.000 43.120 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 450.240 1150.000 450.800 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 464.800 1150.000 465.360 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 479.360 1150.000 479.920 ;
    END
  END io_in[32]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.999200 ;
    ANTENNADIFFAREA 1.315500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 57.120 1150.000 57.680 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.999200 ;
    ANTENNADIFFAREA 1.315500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 71.680 1150.000 72.240 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.999200 ;
    ANTENNADIFFAREA 1.315500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 86.240 1150.000 86.800 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.999200 ;
    ANTENNADIFFAREA 1.315500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 100.800 1150.000 101.360 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.999200 ;
    ANTENNADIFFAREA 1.315500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 115.360 1150.000 115.920 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 129.920 1150.000 130.480 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 144.480 1150.000 145.040 ;
    END
  END io_in[9]
  PIN io_oeb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 574.560 796.000 575.120 800.000 ;
    END
  END io_oeb
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 493.920 1150.000 494.480 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 639.520 1150.000 640.080 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 654.080 1150.000 654.640 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 668.640 1150.000 669.200 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 683.200 1150.000 683.760 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 697.760 1150.000 698.320 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 712.320 1150.000 712.880 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 726.880 1150.000 727.440 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 741.440 1150.000 742.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 756.000 1150.000 756.560 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 770.560 1150.000 771.120 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 508.480 1150.000 509.040 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 785.120 1150.000 785.680 ;
    END
  END io_out[20]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 523.040 1150.000 523.600 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 537.600 1150.000 538.160 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 552.160 1150.000 552.720 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 566.720 1150.000 567.280 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 581.280 1150.000 581.840 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 595.840 1150.000 596.400 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 610.400 1150.000 610.960 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 624.960 1150.000 625.520 ;
    END
  END io_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 861.280 0.000 861.840 4.000 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 784.300 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 784.300 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.352000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 286.720 0.000 287.280 4.000 ;
    END
  END wb_clk_i
  OBS
      LAYER Pwell ;
        RECT 6.290 782.230 1143.390 784.430 ;
      LAYER Nwell ;
        RECT 6.290 777.930 1143.390 782.230 ;
      LAYER Pwell ;
        RECT 6.290 774.390 1143.390 777.930 ;
      LAYER Nwell ;
        RECT 6.290 770.090 1143.390 774.390 ;
      LAYER Pwell ;
        RECT 6.290 766.550 1143.390 770.090 ;
      LAYER Nwell ;
        RECT 6.290 762.250 1143.390 766.550 ;
      LAYER Pwell ;
        RECT 6.290 758.710 1143.390 762.250 ;
      LAYER Nwell ;
        RECT 6.290 754.410 1143.390 758.710 ;
      LAYER Pwell ;
        RECT 6.290 750.870 1143.390 754.410 ;
      LAYER Nwell ;
        RECT 6.290 746.570 1143.390 750.870 ;
      LAYER Pwell ;
        RECT 6.290 743.030 1143.390 746.570 ;
      LAYER Nwell ;
        RECT 6.290 738.730 1143.390 743.030 ;
      LAYER Pwell ;
        RECT 6.290 735.190 1143.390 738.730 ;
      LAYER Nwell ;
        RECT 6.290 730.890 1143.390 735.190 ;
      LAYER Pwell ;
        RECT 6.290 727.350 1143.390 730.890 ;
      LAYER Nwell ;
        RECT 6.290 723.050 1143.390 727.350 ;
      LAYER Pwell ;
        RECT 6.290 719.510 1143.390 723.050 ;
      LAYER Nwell ;
        RECT 6.290 715.210 1143.390 719.510 ;
      LAYER Pwell ;
        RECT 6.290 711.670 1143.390 715.210 ;
      LAYER Nwell ;
        RECT 6.290 707.370 1143.390 711.670 ;
      LAYER Pwell ;
        RECT 6.290 703.830 1143.390 707.370 ;
      LAYER Nwell ;
        RECT 6.290 699.530 1143.390 703.830 ;
      LAYER Pwell ;
        RECT 6.290 695.990 1143.390 699.530 ;
      LAYER Nwell ;
        RECT 6.290 691.690 1143.390 695.990 ;
      LAYER Pwell ;
        RECT 6.290 688.150 1143.390 691.690 ;
      LAYER Nwell ;
        RECT 6.290 683.850 1143.390 688.150 ;
      LAYER Pwell ;
        RECT 6.290 680.310 1143.390 683.850 ;
      LAYER Nwell ;
        RECT 6.290 676.010 1143.390 680.310 ;
      LAYER Pwell ;
        RECT 6.290 672.470 1143.390 676.010 ;
      LAYER Nwell ;
        RECT 6.290 668.170 1143.390 672.470 ;
      LAYER Pwell ;
        RECT 6.290 664.630 1143.390 668.170 ;
      LAYER Nwell ;
        RECT 6.290 660.330 1143.390 664.630 ;
      LAYER Pwell ;
        RECT 6.290 656.790 1143.390 660.330 ;
      LAYER Nwell ;
        RECT 6.290 652.490 1143.390 656.790 ;
      LAYER Pwell ;
        RECT 6.290 648.950 1143.390 652.490 ;
      LAYER Nwell ;
        RECT 6.290 644.650 1143.390 648.950 ;
      LAYER Pwell ;
        RECT 6.290 641.110 1143.390 644.650 ;
      LAYER Nwell ;
        RECT 6.290 636.810 1143.390 641.110 ;
      LAYER Pwell ;
        RECT 6.290 633.270 1143.390 636.810 ;
      LAYER Nwell ;
        RECT 6.290 628.970 1143.390 633.270 ;
      LAYER Pwell ;
        RECT 6.290 625.430 1143.390 628.970 ;
      LAYER Nwell ;
        RECT 6.290 621.130 1143.390 625.430 ;
      LAYER Pwell ;
        RECT 6.290 617.590 1143.390 621.130 ;
      LAYER Nwell ;
        RECT 6.290 613.290 1143.390 617.590 ;
      LAYER Pwell ;
        RECT 6.290 609.750 1143.390 613.290 ;
      LAYER Nwell ;
        RECT 6.290 605.450 1143.390 609.750 ;
      LAYER Pwell ;
        RECT 6.290 601.910 1143.390 605.450 ;
      LAYER Nwell ;
        RECT 6.290 597.610 1143.390 601.910 ;
      LAYER Pwell ;
        RECT 6.290 594.070 1143.390 597.610 ;
      LAYER Nwell ;
        RECT 6.290 589.770 1143.390 594.070 ;
      LAYER Pwell ;
        RECT 6.290 586.230 1143.390 589.770 ;
      LAYER Nwell ;
        RECT 6.290 581.930 1143.390 586.230 ;
      LAYER Pwell ;
        RECT 6.290 578.390 1143.390 581.930 ;
      LAYER Nwell ;
        RECT 6.290 574.090 1143.390 578.390 ;
      LAYER Pwell ;
        RECT 6.290 570.550 1143.390 574.090 ;
      LAYER Nwell ;
        RECT 6.290 566.250 1143.390 570.550 ;
      LAYER Pwell ;
        RECT 6.290 562.710 1143.390 566.250 ;
      LAYER Nwell ;
        RECT 6.290 558.410 1143.390 562.710 ;
      LAYER Pwell ;
        RECT 6.290 554.870 1143.390 558.410 ;
      LAYER Nwell ;
        RECT 6.290 550.570 1143.390 554.870 ;
      LAYER Pwell ;
        RECT 6.290 547.030 1143.390 550.570 ;
      LAYER Nwell ;
        RECT 6.290 542.730 1143.390 547.030 ;
      LAYER Pwell ;
        RECT 6.290 539.190 1143.390 542.730 ;
      LAYER Nwell ;
        RECT 6.290 534.890 1143.390 539.190 ;
      LAYER Pwell ;
        RECT 6.290 531.350 1143.390 534.890 ;
      LAYER Nwell ;
        RECT 6.290 527.050 1143.390 531.350 ;
      LAYER Pwell ;
        RECT 6.290 523.510 1143.390 527.050 ;
      LAYER Nwell ;
        RECT 6.290 519.210 1143.390 523.510 ;
      LAYER Pwell ;
        RECT 6.290 515.670 1143.390 519.210 ;
      LAYER Nwell ;
        RECT 6.290 511.370 1143.390 515.670 ;
      LAYER Pwell ;
        RECT 6.290 507.830 1143.390 511.370 ;
      LAYER Nwell ;
        RECT 6.290 503.530 1143.390 507.830 ;
      LAYER Pwell ;
        RECT 6.290 499.990 1143.390 503.530 ;
      LAYER Nwell ;
        RECT 6.290 495.690 1143.390 499.990 ;
      LAYER Pwell ;
        RECT 6.290 492.150 1143.390 495.690 ;
      LAYER Nwell ;
        RECT 6.290 487.850 1143.390 492.150 ;
      LAYER Pwell ;
        RECT 6.290 484.310 1143.390 487.850 ;
      LAYER Nwell ;
        RECT 6.290 480.010 1143.390 484.310 ;
      LAYER Pwell ;
        RECT 6.290 476.470 1143.390 480.010 ;
      LAYER Nwell ;
        RECT 6.290 472.170 1143.390 476.470 ;
      LAYER Pwell ;
        RECT 6.290 468.630 1143.390 472.170 ;
      LAYER Nwell ;
        RECT 6.290 464.330 1143.390 468.630 ;
      LAYER Pwell ;
        RECT 6.290 460.790 1143.390 464.330 ;
      LAYER Nwell ;
        RECT 6.290 456.490 1143.390 460.790 ;
      LAYER Pwell ;
        RECT 6.290 452.950 1143.390 456.490 ;
      LAYER Nwell ;
        RECT 6.290 448.650 1143.390 452.950 ;
      LAYER Pwell ;
        RECT 6.290 445.110 1143.390 448.650 ;
      LAYER Nwell ;
        RECT 6.290 440.810 1143.390 445.110 ;
      LAYER Pwell ;
        RECT 6.290 437.270 1143.390 440.810 ;
      LAYER Nwell ;
        RECT 6.290 432.970 1143.390 437.270 ;
      LAYER Pwell ;
        RECT 6.290 429.430 1143.390 432.970 ;
      LAYER Nwell ;
        RECT 6.290 425.130 1143.390 429.430 ;
      LAYER Pwell ;
        RECT 6.290 421.590 1143.390 425.130 ;
      LAYER Nwell ;
        RECT 6.290 417.290 1143.390 421.590 ;
      LAYER Pwell ;
        RECT 6.290 413.750 1143.390 417.290 ;
      LAYER Nwell ;
        RECT 6.290 409.450 1143.390 413.750 ;
      LAYER Pwell ;
        RECT 6.290 405.910 1143.390 409.450 ;
      LAYER Nwell ;
        RECT 6.290 401.610 1143.390 405.910 ;
      LAYER Pwell ;
        RECT 6.290 398.070 1143.390 401.610 ;
      LAYER Nwell ;
        RECT 6.290 393.770 1143.390 398.070 ;
      LAYER Pwell ;
        RECT 6.290 390.230 1143.390 393.770 ;
      LAYER Nwell ;
        RECT 6.290 385.930 1143.390 390.230 ;
      LAYER Pwell ;
        RECT 6.290 382.390 1143.390 385.930 ;
      LAYER Nwell ;
        RECT 6.290 378.090 1143.390 382.390 ;
      LAYER Pwell ;
        RECT 6.290 374.550 1143.390 378.090 ;
      LAYER Nwell ;
        RECT 6.290 370.250 1143.390 374.550 ;
      LAYER Pwell ;
        RECT 6.290 366.710 1143.390 370.250 ;
      LAYER Nwell ;
        RECT 6.290 362.410 1143.390 366.710 ;
      LAYER Pwell ;
        RECT 6.290 358.870 1143.390 362.410 ;
      LAYER Nwell ;
        RECT 6.290 354.570 1143.390 358.870 ;
      LAYER Pwell ;
        RECT 6.290 351.030 1143.390 354.570 ;
      LAYER Nwell ;
        RECT 6.290 346.730 1143.390 351.030 ;
      LAYER Pwell ;
        RECT 6.290 343.190 1143.390 346.730 ;
      LAYER Nwell ;
        RECT 6.290 338.890 1143.390 343.190 ;
      LAYER Pwell ;
        RECT 6.290 335.350 1143.390 338.890 ;
      LAYER Nwell ;
        RECT 6.290 331.050 1143.390 335.350 ;
      LAYER Pwell ;
        RECT 6.290 327.510 1143.390 331.050 ;
      LAYER Nwell ;
        RECT 6.290 323.210 1143.390 327.510 ;
      LAYER Pwell ;
        RECT 6.290 319.670 1143.390 323.210 ;
      LAYER Nwell ;
        RECT 6.290 315.370 1143.390 319.670 ;
      LAYER Pwell ;
        RECT 6.290 311.830 1143.390 315.370 ;
      LAYER Nwell ;
        RECT 6.290 307.530 1143.390 311.830 ;
      LAYER Pwell ;
        RECT 6.290 303.990 1143.390 307.530 ;
      LAYER Nwell ;
        RECT 6.290 299.690 1143.390 303.990 ;
      LAYER Pwell ;
        RECT 6.290 296.150 1143.390 299.690 ;
      LAYER Nwell ;
        RECT 6.290 291.850 1143.390 296.150 ;
      LAYER Pwell ;
        RECT 6.290 288.310 1143.390 291.850 ;
      LAYER Nwell ;
        RECT 6.290 284.010 1143.390 288.310 ;
      LAYER Pwell ;
        RECT 6.290 280.470 1143.390 284.010 ;
      LAYER Nwell ;
        RECT 6.290 276.170 1143.390 280.470 ;
      LAYER Pwell ;
        RECT 6.290 272.630 1143.390 276.170 ;
      LAYER Nwell ;
        RECT 6.290 268.330 1143.390 272.630 ;
      LAYER Pwell ;
        RECT 6.290 264.790 1143.390 268.330 ;
      LAYER Nwell ;
        RECT 6.290 260.490 1143.390 264.790 ;
      LAYER Pwell ;
        RECT 6.290 256.950 1143.390 260.490 ;
      LAYER Nwell ;
        RECT 6.290 252.650 1143.390 256.950 ;
      LAYER Pwell ;
        RECT 6.290 249.110 1143.390 252.650 ;
      LAYER Nwell ;
        RECT 6.290 244.810 1143.390 249.110 ;
      LAYER Pwell ;
        RECT 6.290 241.270 1143.390 244.810 ;
      LAYER Nwell ;
        RECT 6.290 236.970 1143.390 241.270 ;
      LAYER Pwell ;
        RECT 6.290 233.430 1143.390 236.970 ;
      LAYER Nwell ;
        RECT 6.290 229.130 1143.390 233.430 ;
      LAYER Pwell ;
        RECT 6.290 225.590 1143.390 229.130 ;
      LAYER Nwell ;
        RECT 6.290 221.290 1143.390 225.590 ;
      LAYER Pwell ;
        RECT 6.290 217.750 1143.390 221.290 ;
      LAYER Nwell ;
        RECT 6.290 213.450 1143.390 217.750 ;
      LAYER Pwell ;
        RECT 6.290 209.910 1143.390 213.450 ;
      LAYER Nwell ;
        RECT 6.290 205.610 1143.390 209.910 ;
      LAYER Pwell ;
        RECT 6.290 202.070 1143.390 205.610 ;
      LAYER Nwell ;
        RECT 6.290 197.770 1143.390 202.070 ;
      LAYER Pwell ;
        RECT 6.290 194.230 1143.390 197.770 ;
      LAYER Nwell ;
        RECT 6.290 189.930 1143.390 194.230 ;
      LAYER Pwell ;
        RECT 6.290 186.390 1143.390 189.930 ;
      LAYER Nwell ;
        RECT 6.290 182.090 1143.390 186.390 ;
      LAYER Pwell ;
        RECT 6.290 178.550 1143.390 182.090 ;
      LAYER Nwell ;
        RECT 6.290 174.250 1143.390 178.550 ;
      LAYER Pwell ;
        RECT 6.290 170.710 1143.390 174.250 ;
      LAYER Nwell ;
        RECT 6.290 166.410 1143.390 170.710 ;
      LAYER Pwell ;
        RECT 6.290 162.870 1143.390 166.410 ;
      LAYER Nwell ;
        RECT 6.290 158.570 1143.390 162.870 ;
      LAYER Pwell ;
        RECT 6.290 155.030 1143.390 158.570 ;
      LAYER Nwell ;
        RECT 6.290 150.730 1143.390 155.030 ;
      LAYER Pwell ;
        RECT 6.290 147.190 1143.390 150.730 ;
      LAYER Nwell ;
        RECT 6.290 142.890 1143.390 147.190 ;
      LAYER Pwell ;
        RECT 6.290 139.350 1143.390 142.890 ;
      LAYER Nwell ;
        RECT 6.290 135.050 1143.390 139.350 ;
      LAYER Pwell ;
        RECT 6.290 131.510 1143.390 135.050 ;
      LAYER Nwell ;
        RECT 6.290 127.210 1143.390 131.510 ;
      LAYER Pwell ;
        RECT 6.290 123.670 1143.390 127.210 ;
      LAYER Nwell ;
        RECT 6.290 119.370 1143.390 123.670 ;
      LAYER Pwell ;
        RECT 6.290 115.830 1143.390 119.370 ;
      LAYER Nwell ;
        RECT 6.290 111.530 1143.390 115.830 ;
      LAYER Pwell ;
        RECT 6.290 107.990 1143.390 111.530 ;
      LAYER Nwell ;
        RECT 6.290 103.690 1143.390 107.990 ;
      LAYER Pwell ;
        RECT 6.290 100.150 1143.390 103.690 ;
      LAYER Nwell ;
        RECT 6.290 95.850 1143.390 100.150 ;
      LAYER Pwell ;
        RECT 6.290 92.310 1143.390 95.850 ;
      LAYER Nwell ;
        RECT 6.290 88.010 1143.390 92.310 ;
      LAYER Pwell ;
        RECT 6.290 84.470 1143.390 88.010 ;
      LAYER Nwell ;
        RECT 6.290 80.170 1143.390 84.470 ;
      LAYER Pwell ;
        RECT 6.290 76.630 1143.390 80.170 ;
      LAYER Nwell ;
        RECT 6.290 72.330 1143.390 76.630 ;
      LAYER Pwell ;
        RECT 6.290 68.790 1143.390 72.330 ;
      LAYER Nwell ;
        RECT 6.290 64.490 1143.390 68.790 ;
      LAYER Pwell ;
        RECT 6.290 60.950 1143.390 64.490 ;
      LAYER Nwell ;
        RECT 6.290 56.650 1143.390 60.950 ;
      LAYER Pwell ;
        RECT 6.290 53.110 1143.390 56.650 ;
      LAYER Nwell ;
        RECT 6.290 48.810 1143.390 53.110 ;
      LAYER Pwell ;
        RECT 6.290 45.270 1143.390 48.810 ;
      LAYER Nwell ;
        RECT 6.290 40.970 1143.390 45.270 ;
      LAYER Pwell ;
        RECT 6.290 37.430 1143.390 40.970 ;
      LAYER Nwell ;
        RECT 6.290 33.130 1143.390 37.430 ;
      LAYER Pwell ;
        RECT 6.290 29.590 1143.390 33.130 ;
      LAYER Nwell ;
        RECT 6.290 25.290 1143.390 29.590 ;
      LAYER Pwell ;
        RECT 6.290 21.750 1143.390 25.290 ;
      LAYER Nwell ;
        RECT 6.290 17.450 1143.390 21.750 ;
      LAYER Pwell ;
        RECT 6.290 15.250 1143.390 17.450 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 1142.960 784.970 ;
      LAYER Metal2 ;
        RECT 7.980 795.700 574.260 796.000 ;
        RECT 575.420 795.700 1142.260 796.000 ;
        RECT 7.980 4.300 1142.260 795.700 ;
        RECT 7.980 4.000 286.420 4.300 ;
        RECT 287.580 4.000 860.980 4.300 ;
        RECT 862.140 4.000 1142.260 4.300 ;
      LAYER Metal3 ;
        RECT 7.930 785.980 1146.740 792.260 ;
        RECT 7.930 784.820 1145.700 785.980 ;
        RECT 7.930 771.420 1146.740 784.820 ;
        RECT 7.930 770.260 1145.700 771.420 ;
        RECT 7.930 756.860 1146.740 770.260 ;
        RECT 7.930 755.700 1145.700 756.860 ;
        RECT 7.930 742.300 1146.740 755.700 ;
        RECT 7.930 741.140 1145.700 742.300 ;
        RECT 7.930 727.740 1146.740 741.140 ;
        RECT 7.930 726.580 1145.700 727.740 ;
        RECT 7.930 713.180 1146.740 726.580 ;
        RECT 7.930 712.020 1145.700 713.180 ;
        RECT 7.930 698.620 1146.740 712.020 ;
        RECT 7.930 697.460 1145.700 698.620 ;
        RECT 7.930 684.060 1146.740 697.460 ;
        RECT 7.930 682.900 1145.700 684.060 ;
        RECT 7.930 669.500 1146.740 682.900 ;
        RECT 7.930 668.340 1145.700 669.500 ;
        RECT 7.930 654.940 1146.740 668.340 ;
        RECT 7.930 653.780 1145.700 654.940 ;
        RECT 7.930 640.380 1146.740 653.780 ;
        RECT 7.930 639.220 1145.700 640.380 ;
        RECT 7.930 625.820 1146.740 639.220 ;
        RECT 7.930 624.660 1145.700 625.820 ;
        RECT 7.930 611.260 1146.740 624.660 ;
        RECT 7.930 610.100 1145.700 611.260 ;
        RECT 7.930 596.700 1146.740 610.100 ;
        RECT 7.930 595.540 1145.700 596.700 ;
        RECT 7.930 582.140 1146.740 595.540 ;
        RECT 7.930 580.980 1145.700 582.140 ;
        RECT 7.930 567.580 1146.740 580.980 ;
        RECT 7.930 566.420 1145.700 567.580 ;
        RECT 7.930 553.020 1146.740 566.420 ;
        RECT 7.930 551.860 1145.700 553.020 ;
        RECT 7.930 538.460 1146.740 551.860 ;
        RECT 7.930 537.300 1145.700 538.460 ;
        RECT 7.930 523.900 1146.740 537.300 ;
        RECT 7.930 522.740 1145.700 523.900 ;
        RECT 7.930 509.340 1146.740 522.740 ;
        RECT 7.930 508.180 1145.700 509.340 ;
        RECT 7.930 494.780 1146.740 508.180 ;
        RECT 7.930 493.620 1145.700 494.780 ;
        RECT 7.930 480.220 1146.740 493.620 ;
        RECT 7.930 479.060 1145.700 480.220 ;
        RECT 7.930 465.660 1146.740 479.060 ;
        RECT 7.930 464.500 1145.700 465.660 ;
        RECT 7.930 451.100 1146.740 464.500 ;
        RECT 7.930 449.940 1145.700 451.100 ;
        RECT 7.930 436.540 1146.740 449.940 ;
        RECT 7.930 435.380 1145.700 436.540 ;
        RECT 7.930 421.980 1146.740 435.380 ;
        RECT 7.930 420.820 1145.700 421.980 ;
        RECT 7.930 407.420 1146.740 420.820 ;
        RECT 7.930 406.260 1145.700 407.420 ;
        RECT 7.930 392.860 1146.740 406.260 ;
        RECT 7.930 391.700 1145.700 392.860 ;
        RECT 7.930 378.300 1146.740 391.700 ;
        RECT 7.930 377.140 1145.700 378.300 ;
        RECT 7.930 363.740 1146.740 377.140 ;
        RECT 7.930 362.580 1145.700 363.740 ;
        RECT 7.930 349.180 1146.740 362.580 ;
        RECT 7.930 348.020 1145.700 349.180 ;
        RECT 7.930 334.620 1146.740 348.020 ;
        RECT 7.930 333.460 1145.700 334.620 ;
        RECT 7.930 320.060 1146.740 333.460 ;
        RECT 7.930 318.900 1145.700 320.060 ;
        RECT 7.930 305.500 1146.740 318.900 ;
        RECT 7.930 304.340 1145.700 305.500 ;
        RECT 7.930 290.940 1146.740 304.340 ;
        RECT 7.930 289.780 1145.700 290.940 ;
        RECT 7.930 276.380 1146.740 289.780 ;
        RECT 7.930 275.220 1145.700 276.380 ;
        RECT 7.930 261.820 1146.740 275.220 ;
        RECT 7.930 260.660 1145.700 261.820 ;
        RECT 7.930 247.260 1146.740 260.660 ;
        RECT 7.930 246.100 1145.700 247.260 ;
        RECT 7.930 232.700 1146.740 246.100 ;
        RECT 7.930 231.540 1145.700 232.700 ;
        RECT 7.930 218.140 1146.740 231.540 ;
        RECT 7.930 216.980 1145.700 218.140 ;
        RECT 7.930 203.580 1146.740 216.980 ;
        RECT 7.930 202.420 1145.700 203.580 ;
        RECT 7.930 189.020 1146.740 202.420 ;
        RECT 7.930 187.860 1145.700 189.020 ;
        RECT 7.930 174.460 1146.740 187.860 ;
        RECT 7.930 173.300 1145.700 174.460 ;
        RECT 7.930 159.900 1146.740 173.300 ;
        RECT 7.930 158.740 1145.700 159.900 ;
        RECT 7.930 145.340 1146.740 158.740 ;
        RECT 7.930 144.180 1145.700 145.340 ;
        RECT 7.930 130.780 1146.740 144.180 ;
        RECT 7.930 129.620 1145.700 130.780 ;
        RECT 7.930 116.220 1146.740 129.620 ;
        RECT 7.930 115.060 1145.700 116.220 ;
        RECT 7.930 101.660 1146.740 115.060 ;
        RECT 7.930 100.500 1145.700 101.660 ;
        RECT 7.930 87.100 1146.740 100.500 ;
        RECT 7.930 85.940 1145.700 87.100 ;
        RECT 7.930 72.540 1146.740 85.940 ;
        RECT 7.930 71.380 1145.700 72.540 ;
        RECT 7.930 57.980 1146.740 71.380 ;
        RECT 7.930 56.820 1145.700 57.980 ;
        RECT 7.930 43.420 1146.740 56.820 ;
        RECT 7.930 42.260 1145.700 43.420 ;
        RECT 7.930 28.860 1146.740 42.260 ;
        RECT 7.930 27.700 1145.700 28.860 ;
        RECT 7.930 14.300 1146.740 27.700 ;
        RECT 7.930 13.580 1145.700 14.300 ;
      LAYER Metal4 ;
        RECT 13.580 25.290 21.940 767.670 ;
        RECT 24.140 25.290 98.740 767.670 ;
        RECT 100.940 25.290 175.540 767.670 ;
        RECT 177.740 25.290 252.340 767.670 ;
        RECT 254.540 25.290 329.140 767.670 ;
        RECT 331.340 25.290 405.940 767.670 ;
        RECT 408.140 25.290 482.740 767.670 ;
        RECT 484.940 25.290 559.540 767.670 ;
        RECT 561.740 25.290 636.340 767.670 ;
        RECT 638.540 25.290 713.140 767.670 ;
        RECT 715.340 25.290 789.940 767.670 ;
        RECT 792.140 25.290 866.740 767.670 ;
        RECT 868.940 25.290 943.540 767.670 ;
        RECT 945.740 25.290 1020.340 767.670 ;
        RECT 1022.540 25.290 1097.140 767.670 ;
        RECT 1099.340 25.290 1133.860 767.670 ;
  END
END wrapped_sid
END LIBRARY

