* NGSPICE file created from wrapped_qcpu.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

.subckt wrapped_qcpu custom_settings[0] custom_settings[10] custom_settings[11] custom_settings[12]
+ custom_settings[13] custom_settings[14] custom_settings[15] custom_settings[16]
+ custom_settings[17] custom_settings[18] custom_settings[19] custom_settings[1] custom_settings[20]
+ custom_settings[21] custom_settings[22] custom_settings[23] custom_settings[24]
+ custom_settings[25] custom_settings[26] custom_settings[27] custom_settings[28]
+ custom_settings[29] custom_settings[2] custom_settings[30] custom_settings[31] custom_settings[3]
+ custom_settings[4] custom_settings[5] custom_settings[6] custom_settings[7] custom_settings[8]
+ custom_settings[9] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15]
+ io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23]
+ io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31]
+ io_in[32] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0]
+ io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17]
+ io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[24] io_oeb[25] io_oeb[26]
+ io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[3]
+ io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10]
+ io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18]
+ io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25]
+ io_out[27] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[3] io_out[4]
+ io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] rst_n sram_addr[0] sram_addr[1]
+ sram_addr[2] sram_addr[3] sram_addr[4] sram_addr[5] sram_gwe sram_in[0] sram_in[1]
+ sram_in[2] sram_in[3] sram_in[4] sram_in[5] sram_in[6] sram_in[7] sram_out[0] sram_out[1]
+ sram_out[2] sram_out[3] sram_out[4] sram_out[5] sram_out[6] sram_out[7] vdd vss
+ wb_clk_i io_oeb[23] io_oeb[22] io_out[28] io_out[26]
X_05903_ _01385_ cpu.uart.divisor\[9\] _01196_ _01386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09671_ _04204_ _04680_ _04681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06883_ _02041_ _02044_ _02359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_27_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05834_ _01302_ _01304_ _01318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08622_ _03750_ _03773_ _03774_ _00344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_89_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05765_ _01237_ _01240_ _01244_ _01248_ _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_08553_ cpu.toggle_top\[15\] _03717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09287__A1 cpu.PC\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08484_ _03045_ _03651_ _03663_ _03653_ _00317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07504_ _01360_ _02900_ _02902_ _00098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07435_ cpu.uart.receive_div_counter\[15\] _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_81_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05696_ _01126_ _01180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_49_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05848__A1 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07051__C _02518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07366_ _02783_ _02552_ _02784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06317_ _01788_ _01370_ _01794_ _01795_ _01489_ _01796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_09105_ _04152_ _00449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07297_ _02727_ _02719_ _02728_ _02724_ _00065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09036_ _01110_ _04069_ _04071_ _04098_ _04094_ _04099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_06248_ _01725_ _01728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06462__I _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09211__A1 _00950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05078__I _00571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06179_ _01643_ _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_92_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09938_ cpu.PORTB_DDR\[2\] _04892_ _04899_ _04897_ _04900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_5_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09869_ _04031_ _04845_ _04848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09278__A1 _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output37_I net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10644_ _00538_ clknet_leaf_60_wb_clk_i cpu.PORTB_DDR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_70_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10575_ _00469_ clknet_leaf_81_wb_clk_i cpu.last_addr\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer7 _00872_ net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_51_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06567__A2 _01001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05716__I _01199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_60_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_60_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10009_ net65 _04945_ _04947_ _04954_ _02620_ _04955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_05550_ _01027_ _01030_ _01033_ _01034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_19_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05481_ _00760_ _00967_ _00968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_58_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07220_ cpu.timer\[1\] _02666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07151_ _02606_ _02598_ _02607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06102_ _01583_ _01584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09992__A2 _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07082_ _02317_ _02318_ _02547_ _02548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06215__C _01121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06033_ cpu.timer_top\[2\] _01240_ _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07984_ cpu.spi.div_counter\[4\] _03264_ _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09723_ _04728_ _00491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06935_ _02150_ _02340_ _02408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08937__I _04002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09654_ _04382_ _04650_ _04664_ _04406_ _04665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06866_ _02338_ _02341_ _02342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_38_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08605_ _02882_ _03748_ _03762_ _03763_ _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_05817_ _01299_ _01300_ _01301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09585_ _04575_ _04592_ _04595_ _04598_ _04081_ _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_49_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06797_ _02269_ _02272_ _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_05748_ _01037_ _01061_ _01185_ _01232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_08536_ _03700_ _00332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06457__I _01934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08483__A2 _03609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08467_ cpu.orig_PC\[3\] _03636_ _03652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05679_ _01162_ _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08398_ _03598_ _03599_ _03600_ _00294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_108_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07418_ cpu.uart.receive_div_counter\[10\] _02829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07349_ _02767_ _02768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06246__A1 _00985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10360_ _00255_ clknet_leaf_36_wb_clk_i cpu.uart.div_counter\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06246__B2 _01336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09019_ cpu.orig_IO_addr_buff\[1\] _04075_ _04076_ _02668_ _04085_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10291_ _00186_ clknet_leaf_107_wb_clk_i cpu.regs\[2\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07746__A1 _01358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09008__I _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05472__S _00851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05080__S1 _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06485__A1 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10627_ _00521_ clknet_leaf_68_wb_clk_i net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07198__I _02646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10558_ _00452_ clknet_leaf_79_wb_clk_i cpu.ROM_addr_buff\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10489_ _00384_ clknet_leaf_27_wb_clk_i cpu.timer\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05446__I _00933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06720_ _02193_ _02195_ _02192_ _02196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06651_ _02100_ _02101_ _02127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05602_ _01083_ _01085_ _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09370_ _04387_ _04386_ _04389_ _04390_ _04391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06582_ _02049_ _02050_ _02057_ _02058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__05071__S1 _00575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08321_ _03515_ _02863_ _03538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05533_ _01016_ _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_46_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08252_ _03464_ _03486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05464_ _00951_ _00952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_47_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07203_ _01863_ _02651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_104_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08183_ _03344_ _03425_ _03430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05395_ cpu.regs\[0\]\[1\] cpu.regs\[1\]\[1\] cpu.regs\[2\]\[1\] cpu.regs\[3\]\[1\]
+ _00882_ _00884_ _00885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10024__A2 _02583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07134_ _02592_ _02587_ _02594_ _02589_ _00036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_42_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07065_ _02524_ _02525_ _02530_ _02531_ _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06016_ _01496_ _01497_ _01122_ _01498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_76_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08441__B _03633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05451__A2 _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09256__C _04270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07967_ _03250_ _03252_ _03254_ _03255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05203__A2 _00717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09706_ _04674_ _04714_ _04713_ _04715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06918_ _02391_ _02392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07898_ _03095_ _03195_ _03196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08153__A1 _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07571__I _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09637_ _02367_ cpu.PC\[13\] _04500_ _04648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06849_ _02265_ _02323_ _02324_ _02325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_87_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09568_ _04578_ _04581_ _04582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08519_ _02742_ _03680_ _03688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09653__A1 _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09499_ _04509_ _04513_ _04515_ _04516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07416__B1 cpu.uart.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10412_ _00307_ clknet_leaf_56_wb_clk_i cpu.orig_flags\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10343_ _00238_ clknet_leaf_62_wb_clk_i cpu.spi.counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10274_ _00169_ clknet_leaf_111_wb_clk_i cpu.regs\[5\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07719__A1 _01359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_14_Left_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_104_Right_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05180_ net71 _00696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07958__A1 _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09357__B _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Left_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08870_ _00967_ _03955_ _03966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07821_ cpu.timer_div_counter\[5\] _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07752_ _02241_ _02325_ _02326_ _03062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06703_ _02175_ _02176_ _02179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_32_Left_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07683_ _02985_ _03011_ _03015_ _00164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09820__B _03474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09422_ _04383_ _04423_ _04441_ _04407_ _04442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06634_ _00831_ _01287_ _02110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09353_ _04226_ _04375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08304_ cpu.uart.receive_buff\[1\] _03523_ _03526_ cpu.uart.receive_buff\[2\] _03528_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_4_5_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06565_ _02024_ _02040_ _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__09635__A1 _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06449__A1 _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09284_ _04303_ _04305_ _04306_ _04307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06496_ _01953_ _01971_ _01325_ _01973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05516_ _00849_ _01001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08235_ cpu.uart.counter\[0\] cpu.uart.counter\[1\] _03456_ cpu.uart.counter\[3\]
+ _03472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_62_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05447_ _00934_ _00935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_34_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08166_ _03415_ _03416_ _00246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05378_ _00863_ _00866_ _00867_ _00868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_31_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07117_ _02499_ _02580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_42_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_41_Left_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08097_ cpu.uart.data_buff\[0\] _03360_ _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07048_ _00683_ _02516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_30_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_89_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08999_ _04058_ _04065_ _02609_ _04066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08397__I _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05814__I cpu.base_address\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05283__S1 _00786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09874__A1 _04851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_117_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_117_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_66_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08062__B1 _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10326_ _00221_ clknet_leaf_50_wb_clk_i cpu.spi.data_in_buff\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05415__A2 _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10257_ _00152_ clknet_leaf_117_wb_clk_i cpu.regs\[7\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08365__A1 _02830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10188_ _00083_ clknet_leaf_14_wb_clk_i _00001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05724__I _01207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05351__A1 net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06350_ _01818_ _01828_ _01829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06281_ _01633_ _00977_ _01761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05301_ cpu.regs\[8\]\[1\] cpu.regs\[9\]\[1\] cpu.regs\[10\]\[1\] cpu.regs\[11\]\[1\]
+ _00568_ _00573_ _00811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08020_ _03289_ _03295_ _00221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_72_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05232_ _00701_ _00745_ _00746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_21_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05163_ _00671_ _00679_ _00680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09971_ _03231_ _04916_ _04924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_73_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05094_ _00613_ net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_0_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08922_ _04004_ _00414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08853_ _03952_ _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07804_ _01510_ _03102_ _03108_ _00192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08784_ _03131_ _03894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05996_ _01478_ _01479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07735_ _03045_ _02058_ _03046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_67_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07666_ _01857_ _03004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09405_ cpu.PC\[3\] _01134_ _04424_ _04425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_62_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06617_ _00831_ _02093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07597_ _01584_ _02961_ _00132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06548_ _00682_ _00688_ _02024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_75_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09336_ _04061_ _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09267_ _02511_ _04291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_51_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08218_ cpu.uart.counter\[3\] _03456_ _03359_ _03457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06479_ _01955_ _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05645__A2 _01128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09198_ _00926_ _04218_ _04223_ _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08149_ _03325_ _03397_ _03403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_95_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07642__I0 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10111_ _05043_ _00564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10042_ _04965_ _04982_ _04984_ _02762_ _00554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_output67_I net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_10_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05581__A1 _01035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08855__I _03942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_85_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_85_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_108_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_14_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_14_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06833__A1 _02270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10309_ _00204_ clknet_leaf_59_wb_clk_i cpu.spi.data_out_buff\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07010__A1 cpu.ROM_addr_buff\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05850_ _00969_ _00715_ _01334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_107_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09838__A1 _03288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05572__A1 _01054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05781_ _01264_ _01265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07520_ _01109_ _01130_ _02911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07451_ _02840_ _02853_ _02858_ _02861_ _02862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_9_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06402_ cpu.timer_div\[6\] _01801_ _01880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07382_ _02557_ _02575_ _02798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06218__C _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09121_ _03672_ _04136_ _04163_ _04164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06333_ cpu.toggle_top\[13\] _01257_ _01812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09052_ cpu.IO_addr_buff\[7\] _04097_ _04111_ _04100_ _04112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_60_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06264_ _01660_ _01662_ _01744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08003_ cpu.spi.div_counter\[7\] _03280_ _03283_ _03279_ _03284_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05215_ _00696_ net18 _00730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_13_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06195_ _01529_ _01633_ _01675_ _01676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05146_ cpu.startup_cycle\[6\] cpu.startup_cycle\[5\] cpu.startup_cycle\[4\] _00663_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__06052__A2 _00923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09954_ _04911_ _00539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05077_ _00597_ net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_110_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09885_ _04045_ _04857_ _04860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08905_ cpu.spi.divisor\[5\] _03990_ _03992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08836_ _03936_ _03937_ _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_79_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08767_ cpu.timer\[3\] _03879_ _03880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_56_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05979_ _01443_ _01451_ _01453_ _01456_ _01461_ _01462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08698_ _03827_ _03828_ _00366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_0_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07718_ cpu.regs\[3\]\[0\] _03036_ _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07649_ cpu.regs\[7\]\[7\] _02979_ _02993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10660_ _00554_ clknet_leaf_74_wb_clk_i net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_36_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09319_ _04273_ _04341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10591_ _00485_ clknet_leaf_84_wb_clk_i cpu.PC\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05618__A2 _01101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput42 net42 io_oeb[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput64 net64 io_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput75 net75 io_out[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput53 net53 io_oeb[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput97 net97 sram_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput86 net86 sram_addr[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10025_ _04670_ _02034_ _04968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07690__S _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05609__A2 _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05449__I _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07231__A1 _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06951_ cpu.startup_cycle\[5\] _02422_ _02423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_118_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05902_ _01370_ _01382_ _01384_ _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09670_ cpu.last_addr\[9\] cpu.last_addr\[8\] _04679_ _04680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06882_ _02017_ _02023_ _02357_ _02358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08621_ cpu.toggle_ctr\[11\] _03703_ _03771_ _03774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XPHY_EDGE_ROW_6_Left_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05833_ _01315_ _01316_ _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05764_ cpu.timer_top\[0\] _01245_ _01247_ _01248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08552_ cpu.toggle_ctr\[14\] _03714_ _03715_ _03716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08483_ cpu.orig_PC\[8\] _03609_ _03663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07332__C _02753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07503_ cpu.regs\[13\]\[0\] _02901_ _02902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07434_ cpu.uart.divisor\[15\] _02845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_81_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05695_ _01118_ _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_64_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05848__A2 _00878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07365_ _02782_ _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06316_ net11 _01372_ _01200_ _01795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09104_ _04151_ cpu.ROM_addr_buff\[7\] _04148_ _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07296_ cpu.timer_top\[7\] _02720_ _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08798__A1 _03170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09035_ cpu.orig_IO_addr_buff\[4\] _04091_ _04092_ _00967_ _04098_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06247_ _00596_ _00985_ _01727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06178_ _01655_ _01657_ _01658_ _01659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_92_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05129_ _00644_ _00645_ _00646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09275__B _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09937_ _04851_ _04893_ _04899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_5_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09868_ _04847_ _00517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08722__A1 cpu.timer_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09799_ _04791_ _04773_ _04779_ _04792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08819_ _01591_ _03866_ _03923_ _03920_ _00392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_68_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09278__A2 _00757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10643_ _00537_ clknet_leaf_69_wb_clk_i cpu.PORTB_DDR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10574_ _00468_ clknet_leaf_81_wb_clk_i cpu.last_addr\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08789__A1 _02697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer8 _00862_ net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08961__A1 _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06567__A3 _01296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_79_Left_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10008_ _04949_ _04951_ _04953_ _04954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05527__A1 _00711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05732__I _01034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05480_ _00966_ _00967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_27_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_30_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07150_ _01018_ _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09441__A2 _01774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07081_ _02391_ _02319_ _02547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06101_ _01582_ _01583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_112_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06032_ _01486_ _01402_ _01512_ _01513_ _01245_ _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__08711__C _03201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09722_ _03116_ _04727_ _04728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07983_ _03267_ _00212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05310__S0 _00569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06934_ _02406_ _02407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09653_ _00742_ _04390_ _04661_ _04663_ _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06865_ _02339_ _02340_ _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_38_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09584_ _04368_ _04577_ _04597_ _04547_ _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08604_ _03730_ _03760_ _03725_ _03763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05816_ cpu.base_address\[3\] _00714_ _01300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_118_Right_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09114__I _04022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08535_ cpu.toggle_top\[7\] _03690_ _03699_ _03697_ _03700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06796_ _02271_ _00899_ _02267_ _02268_ _02272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_05747_ _01184_ _01229_ _01230_ _01231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08953__I _04025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08466_ _03621_ _03651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05678_ _01161_ _01162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08397_ _03311_ _03600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07417_ cpu.uart.divisor\[10\] _02828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06494__A2 _01957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07348_ _02766_ _02767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07279_ _02624_ _02711_ _02714_ _02716_ _00059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09018_ _03551_ _04084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10290_ _00185_ clknet_leaf_112_wb_clk_i cpu.regs\[3\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08943__A1 _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08349__B _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09959__I _04914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06485__A2 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10626_ _00520_ clknet_leaf_67_wb_clk_i net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_70_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10557_ _00451_ clknet_leaf_87_wb_clk_i cpu.ROM_addr_buff\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_114_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10488_ _00383_ clknet_leaf_24_wb_clk_i cpu.timer\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05727__I _01210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_87_Left_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_4_12_0_wb_clk_i clknet_0_wb_clk_i clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_06650_ _02123_ _02124_ _02125_ _02126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05601_ _01078_ _01084_ _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05462__I _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06581_ cpu.PC\[5\] _02056_ _02057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08320_ cpu.uart.receive_div_counter\[0\] _03537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_96_Left_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05532_ _00745_ _01016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08251_ _03481_ _03483_ _03485_ _00262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_74_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05463_ _00950_ _00951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07202_ cpu.uart.divisor\[7\] _02650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_7_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08182_ _03392_ _03428_ _03429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06226__C _01183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05394_ _00883_ _00884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07133_ _02593_ _02585_ _02594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07064_ _02520_ _02531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06015_ cpu.PORTB_DDR\[2\] _01211_ _01497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_11_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07966_ _03250_ _03253_ _03254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input29_I sram_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09705_ _02461_ _02581_ _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06917_ _02360_ _02391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07897_ _03178_ _03179_ _03186_ _03194_ _03195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_0_69_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09636_ _03674_ _04550_ _04647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09350__A1 _02796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07361__B1 _02668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06848_ _02238_ _02239_ _02324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_87_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09567_ _04557_ _04579_ _04580_ _04581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06779_ _02252_ _02254_ _02255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_38_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09498_ _04388_ _04502_ _04514_ _04362_ _04515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08518_ _03687_ _00327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_38_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08449_ cpu.orig_flags\[2\] _03627_ _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_13_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10411_ _00306_ clknet_leaf_92_wb_clk_i cpu.orig_flags\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output97_I net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10342_ _00237_ clknet_leaf_49_wb_clk_i cpu.spi.counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08916__A1 _03822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10273_ _00168_ clknet_leaf_117_wb_clk_i cpu.regs\[5\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_39_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_39_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09463__B _04273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06155__A1 net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05505__I1 cpu.regs\[9\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10609_ _00503_ clknet_leaf_75_wb_clk_i cpu.ROM_spi_dat_out\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05969__A1 _01298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07820_ cpu.timer_div_counter\[1\] _03119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08768__I _03864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07751_ _03060_ _02059_ _03061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06702_ _02159_ _02160_ _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06146__B2 _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07682_ cpu.regs\[5\]\[2\] _03012_ _03015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09421_ _04429_ _04436_ _04440_ _04441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06633_ _02105_ _02108_ _02109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06941__I0 cpu.regs\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06564_ cpu.rom_data_dist _02039_ _02040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_75_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09352_ _04373_ _04374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08303_ _03519_ _03527_ _00272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05515_ _01000_ net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09283_ _01015_ _04277_ _04270_ _04306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06495_ _01953_ _01971_ _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07340__C _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08234_ _03470_ _03471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05446_ _00933_ _00934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_28_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08165_ _03335_ _03413_ _03276_ _03416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05377_ _00007_ _00867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07116_ _02544_ _02578_ _02579_ _00033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08096_ _03359_ _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05504__S0 _00956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07047_ _02497_ _02514_ _02515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09283__B _04270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08998_ _04059_ _04064_ _04065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07949_ cpu.spi.data_out_buff\[5\] _03230_ _03239_ _03240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_46_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06198__I _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09619_ cpu.PC\[11\] _01155_ _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06688__A2 cpu.regs\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09626__A2 _00763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08062__B2 _02630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10325_ _00220_ clknet_leaf_48_wb_clk_i cpu.spi.data_in_buff\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05415__A3 _00904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10256_ _00151_ clknet_leaf_115_wb_clk_i cpu.regs\[7\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10187_ _00082_ clknet_leaf_13_wb_clk_i _00000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_89_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09617__A2 _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05351__A2 cpu.ROM_spi_mode vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06280_ _01757_ _01759_ _01760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05300_ _00586_ _00809_ _00810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05231_ cpu.br_rel_dest\[4\] _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_4_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05162_ _00673_ _00678_ _00679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_110_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09970_ _04923_ _00543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_73_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05187__I _00701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05093_ _00612_ _00613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_12_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08921_ cpu.timer_div\[1\] _04000_ _04001_ _04003_ _04004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_0_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08852_ cpu.timer_capture\[8\] _03943_ _03950_ _03951_ _03952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07803_ cpu.spi.data_in_buff\[2\] _03107_ _03105_ _03108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08783_ _03892_ _03893_ _00386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07335__C _02753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05995_ _01150_ _01478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__06119__A1 _01598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07734_ _02048_ _03045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07665_ _03003_ _00158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06616_ _02090_ _02091_ _02092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06914__I0 _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09404_ _02802_ _01586_ _04339_ _04393_ _04424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_84_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07596_ _01482_ _02961_ _00131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09335_ _04347_ _04356_ _04357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_23_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06547_ _02022_ _02023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_117_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09266_ _02772_ _04288_ _04289_ _04284_ _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_06478_ _01954_ _01955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08217_ cpu.uart.counter\[2\] _03456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05429_ cpu.regs\[8\]\[2\] cpu.regs\[9\]\[2\] cpu.regs\[10\]\[2\] cpu.regs\[11\]\[2\]
+ _00881_ _00883_ _00918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_105_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09197_ cpu.orig_flags\[2\] _04218_ _04223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08148_ _03401_ _03402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08079_ _03340_ _02650_ _02630_ _03325_ _03342_ _03343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XTAP_TAPCELL_ROW_95_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10110_ _01934_ cpu.regs\[15\]\[6\] _05033_ _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05097__I _00575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10041_ _04759_ _04983_ _04982_ _02475_ _04984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_clkbuf_leaf_123_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_6_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07688__S _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06833__A2 _00908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_54_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_54_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10308_ _00203_ clknet_leaf_58_wb_clk_i cpu.spi.data_out_buff\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_60_Left_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10239_ _00134_ clknet_4_2_0_wb_clk_i cpu.regs\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05780_ _01262_ _01263_ _01264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05572__A2 _01055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07450_ _02859_ cpu.uart.receive_div_counter\[15\] _02822_ _02630_ _02860_ _02861_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__06521__A1 cpu.timer_capture\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06566__I _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06401_ _01865_ _01608_ _01877_ _01878_ _01801_ _01879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_8_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07381_ _02797_ _00080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09120_ _04137_ cpu.regs\[3\]\[4\] _04163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06332_ cpu.toggle_top\[5\] _01178_ _01810_ _01367_ _01811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_29_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09051_ _01133_ _04069_ _04071_ _04110_ _04094_ _04111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__10081__A1 _01734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06515__B _01081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08002_ cpu.spi.div_counter\[7\] _03203_ _03283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06263_ _00597_ _01742_ _01743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05214_ _00668_ _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06194_ _01315_ _01649_ _01665_ _01674_ _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_05145_ cpu.startup_cycle\[1\] cpu.startup_cycle\[0\] _00662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09953_ cpu.PORTB_DDR\[6\] _04903_ _04910_ _04908_ _04911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05260__A1 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05076_ _00596_ _00597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09884_ _04859_ _00521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08904_ _02635_ _03989_ _03991_ _00409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08835_ cpu.timer_capture\[14\] _03913_ _03914_ _03937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08766_ cpu.timer\[2\] cpu.timer\[1\] cpu.timer\[0\] _03879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA_input11_I io_in[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05563__A2 _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07717_ _03033_ _03036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05978_ _01457_ _01458_ _01460_ _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08697_ _03121_ cpu.timer_div_counter\[1\] _03828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_0_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08501__A2 _03626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05380__I _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07560__I0 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07648_ _02013_ _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07579_ _02920_ _02947_ _02951_ _00124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_36_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09318_ _04338_ _04339_ _04340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10590_ _00484_ clknet_leaf_95_wb_clk_i cpu.PC\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_97_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09249_ _00928_ _04272_ _04273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__06815__A2 _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08568__A2 cpu.toggle_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput43 net43 io_oeb[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_31_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06579__A1 _02052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput76 net76 io_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput65 net65 io_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput54 net54 io_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_8_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput87 net87 sram_addr[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10024_ _04940_ _02583_ _04966_ _04670_ _04967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__09027__I _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_101_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_101_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_67_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10063__B2 _01170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06950_ cpu.startup_cycle\[4\] _02422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input3_I io_in[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05901_ cpu.uart.divisor\[1\] _01383_ _01384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_68_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06881_ _02022_ _02356_ _02357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05832_ _01168_ _01305_ _01311_ _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08620_ _03703_ _03771_ cpu.toggle_ctr\[11\] _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06742__A1 _00829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05763_ _01246_ _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08551_ _03711_ cpu.toggle_top\[13\] _03715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08482_ _03661_ _03662_ _03650_ _00316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07298__A2 _00757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05694_ _01177_ _01178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07502_ _02898_ _02901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07433_ _02843_ cpu.uart.receive_div_counter\[12\] cpu.uart.receive_div_counter\[8\]
+ _02831_ _02844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_81_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_77_Right_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_33_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08247__A1 _02707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09103_ cpu.regs\[2\]\[7\] _02570_ _04150_ _04151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_61_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07364_ _02781_ _02782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06315_ net3 _01114_ _01089_ _01793_ _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_07295_ _02726_ _02727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09034_ _04066_ _04097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06246_ _00985_ _01339_ _01725_ _01336_ _01341_ _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_32_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_107_Left_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09747__A1 _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08460__B _03633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09211__A3 _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06177_ _01637_ _01656_ _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_92_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05128_ cpu.IO_addr_buff\[0\] _00645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09936_ _04898_ _00534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_86_Right_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_5_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05059_ _00579_ _00580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09867_ net59 _04844_ _04846_ _04788_ _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_116_Left_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09798_ _04750_ _04764_ _04791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08818_ _03921_ _03825_ _03857_ _03922_ _03865_ _03923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07590__I _01128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08749_ _03864_ _03865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08486__A1 _03664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_95_Right_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10642_ _00536_ clknet_leaf_68_wb_clk_i cpu.PORTB_DDR\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_101_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10573_ _00467_ clknet_leaf_78_wb_clk_i cpu.last_addr\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09986__A1 _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer9 _00854_ net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06567__A4 _01071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10007_ _04952_ _04953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05527__A2 _01010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_67_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09977__A1 cpu.PORTA_DDR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07080_ net12 _02361_ _02045_ _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06100_ _01484_ _01527_ _01581_ _01479_ _01582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_89_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06031_ cpu.timer_capture\[2\] _01235_ _01402_ _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_2_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08280__B _03505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07675__I _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07982_ _02882_ _03265_ _03266_ _03267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_1_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09721_ _04713_ _04710_ _04726_ _04727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06933_ _02405_ _02020_ _02406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05310__S1 _00574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09652_ _04388_ _04650_ _04662_ _04362_ _04663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06864_ _00619_ _01956_ _02340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_38_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09583_ _00818_ _04596_ _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08603_ cpu.toggle_ctr\[5\] cpu.toggle_ctr\[4\] cpu.toggle_ctr\[3\] _03757_ _03762_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_06795_ _00830_ _02271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07343__C _02763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05815_ _01298_ _00712_ _01299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05746_ cpu.timer_div\[0\] _01184_ _01230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08534_ _02652_ _03691_ _03699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08465_ _03647_ _03648_ _03650_ _00311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05677_ _01111_ _01161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08396_ _03593_ _03596_ _03599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07416_ _02821_ _02650_ cpu.uart.divisor\[3\] _02822_ _02826_ _02827_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_80_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09968__A1 _04851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07347_ _02765_ _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07278_ _02715_ _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09017_ _03781_ _04083_ _00430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06229_ cpu.timer_capture\[4\] _01690_ _01706_ _01708_ _01242_ _01709_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09919_ net56 _04880_ _04884_ _04885_ _04886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_output42_I net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09120__A2 cpu.regs\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06485__A3 _01757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07682__A2 _03012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10625_ _00519_ clknet_leaf_67_wb_clk_i net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__10018__A1 cpu.ROM_addr_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09975__I _04914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10556_ _00450_ clknet_leaf_87_wb_clk_i cpu.ROM_addr_buff\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_114_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10487_ _00382_ clknet_leaf_27_wb_clk_i cpu.timer\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09187__A2 _04213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07163__C _02518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05056__S0 _00572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09215__I _02796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05600_ _01058_ _00672_ _01084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06580_ _02051_ _02055_ _02056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_115_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05531_ cpu.br_rel_dest\[1\] _01015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08250_ cpu.uart.data_buff\[2\] _03484_ _03245_ _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08870__A1 _00967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07673__A2 _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05462_ _00949_ _00950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__10009__A1 net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10009__B2 _04954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08181_ _03344_ _03425_ _03428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07201_ _02649_ _00048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_9_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_9_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05393_ _00859_ _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07132_ _01151_ _02593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_70_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07063_ _02526_ _02527_ _02528_ _02529_ _02530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_30_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06014_ _01493_ _01495_ _01211_ _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05918__I cpu.timer_capture\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07965_ _03202_ _03253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09704_ _04672_ _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06916_ _02390_ _00022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07896_ cpu.spi.div_counter\[1\] _03187_ _03188_ cpu.spi.div_counter\[5\] _03193_
+ _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_09635_ _04222_ _04646_ _00485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07361__A1 _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06847_ _02285_ _02321_ _02322_ _02323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09566_ cpu.PC\[9\] _00843_ _04580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06778_ _02253_ _00973_ _02254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05729_ _01068_ _01213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09497_ cpu.orig_PC\[7\] _04074_ _04514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08517_ cpu.toggle_top\[2\] _03679_ _03685_ _03686_ _03687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_38_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08448_ _00779_ _03622_ _03638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08861__A1 _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08379_ cpu.uart.receive_div_counter\[11\] _03585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10410_ _00305_ clknet_leaf_92_wb_clk_i cpu.orig_flags\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10341_ _00236_ clknet_leaf_48_wb_clk_i cpu.spi.counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10272_ _00167_ clknet_leaf_115_wb_clk_i cpu.regs\[5\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_79_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_79_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_79_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_69_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06155__A2 _00976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07352__A1 _01358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08852__A1 cpu.timer_capture\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07655__A2 _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10608_ _00502_ clknet_leaf_76_wb_clk_i cpu.ROM_spi_dat_out\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10539_ _00433_ clknet_leaf_17_wb_clk_i cpu.IO_addr_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06394__A2 _01114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07750_ cpu.PC\[9\] _03060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06701_ _02175_ _02176_ _02177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07343__A1 _02592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07681_ _02983_ _03011_ _03014_ _00163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09420_ _04358_ _04423_ _04438_ _04439_ _04440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06632_ _02106_ _02107_ _02108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06563_ _02027_ _02030_ _02034_ _02038_ _02039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_09351_ _00753_ _04373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08302_ cpu.uart.receive_buff\[0\] _03523_ _03526_ cpu.uart.receive_buff\[1\] _03527_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05514_ _00764_ _00989_ _00999_ _01000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09282_ _02782_ _00762_ _04304_ _04305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08233_ _03364_ _03358_ _03470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06494_ _01895_ _01957_ _01911_ _01971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05445_ _00914_ _00916_ _00921_ _00919_ _00933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_08164_ _03335_ _03405_ _03414_ _03408_ _03415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09548__C _04432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09399__A2 _04379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05376_ cpu.regs\[4\]\[0\] cpu.regs\[5\]\[0\] cpu.regs\[6\]\[0\] cpu.regs\[7\]\[0\]
+ _00864_ _00865_ _00866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_08095_ _03358_ _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_70_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07115_ _02375_ _02544_ _02579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07046_ net20 _02498_ _02514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_42_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05504__S1 _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06082__A1 _01447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09020__A1 _01365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09571__A2 _04484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08997_ _04061_ _04063_ _04064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06479__I _01955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07948_ _02642_ _03225_ _03239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07879_ _03116_ _00698_ _03177_ _00198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07334__A1 _02652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09618_ _04061_ _04626_ _04629_ _04361_ _04630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05896__A1 _01070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09087__A1 _02803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09549_ _00847_ _04430_ _04563_ _04434_ _04564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_66_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05648__A1 _01109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07637__A2 _02981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_126_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_126_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_104_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10324_ _00219_ clknet_leaf_51_wb_clk_i cpu.spi.data_in_buff\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08869__I _03942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10255_ _00150_ clknet_leaf_118_wb_clk_i cpu.regs\[7\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10186_ _00081_ clknet_leaf_100_wb_clk_i cpu.regs\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06376__A2 _01854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07325__A1 _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05431__S0 _00856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05230_ _00657_ cpu.br_rel_dest\[6\] _00744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_114_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05161_ _00674_ _00677_ _00678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09250__A1 _01162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05092_ _00567_ _00606_ _00611_ _00612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08920_ _04002_ _04003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05811__A1 _01170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08851_ _03808_ _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07802_ _03103_ _03107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10042__C _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08782_ cpu.timer_capture\[5\] _03888_ _03889_ _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05994_ _01425_ _01475_ _01476_ _01477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_07733_ _02014_ _03036_ _03044_ _00185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07664_ _03002_ cpu.regs\[6\]\[4\] _02995_ _03003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_94_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09403_ _04422_ _04423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06615_ _02070_ _02071_ _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_48_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07595_ _01360_ _02961_ _00130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09334_ _02593_ _04349_ _04354_ _04355_ _04356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06546_ _02021_ _02022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_23_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09559__B _04523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09265_ _02767_ _04288_ _04289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06477_ _01781_ _01778_ _00871_ _01954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08216_ _03452_ _03360_ _03455_ _03365_ _00257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09196_ _02870_ _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05428_ _00914_ _00916_ _00917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08147_ _02872_ _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09092__I1 cpu.ROM_addr_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09241__A1 _04234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05359_ _00848_ _00849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08078_ _02823_ cpu.uart.div_counter\[9\] _03341_ _02825_ _03342_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_3_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08689__I _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07029_ _02497_ _02499_ _02500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10040_ _04952_ _04967_ _04979_ _04983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07555__A1 cpu.regs\[11\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08638__B _03505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06530__A2 _01784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09232__A1 _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10307_ _00202_ clknet_leaf_57_wb_clk_i cpu.spi.data_out_buff\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_94_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_94_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10238_ _00133_ clknet_leaf_119_wb_clk_i cpu.regs\[0\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_23_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_23_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10169_ _00068_ clknet_leaf_11_wb_clk_i cpu.toggle_top\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06400_ cpu.spi.divisor\[6\] _01606_ _01190_ _01878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_9_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07380_ _02795_ _02796_ _02775_ _02797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06331_ _01808_ _01809_ _01810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09050_ cpu.orig_IO_addr_buff\[7\] _04091_ _04092_ _01291_ _04110_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06262_ _01741_ _01645_ _01642_ _01742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_115_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08001_ _02874_ _03282_ _00215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05213_ _00727_ _00728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09074__I1 cpu.ROM_addr_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06193_ _01468_ _01668_ _01669_ _01671_ _01673_ _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_25_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09223__A1 _01162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05144_ cpu.ROM_spi_cycle\[4\] cpu.ROM_spi_cycle\[1\] cpu.ROM_spi_cycle\[0\] _00660_
+ _00661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
X_09952_ _04048_ _04904_ _04910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05075_ _00567_ _00582_ _00595_ _00596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_08903_ cpu.spi.divisor\[4\] _03990_ _03991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09883_ net63 _04856_ _04858_ _04849_ _04859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08834_ _03933_ _03825_ _03904_ _03935_ _03865_ _03936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08765_ _03874_ _03878_ _03868_ _00383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_56_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07716_ _03034_ _03035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05977_ _00901_ _01338_ _01459_ _01330_ _01147_ _01460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_95_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08696_ cpu.timer_div_counter\[0\] _03827_ _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_0_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06512__A2 _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07647_ _02991_ _00152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07578_ cpu.regs\[10\]\[2\] _02948_ _02951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_36_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06529_ _02005_ _02006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09317_ _02053_ _01151_ _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08193__B _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09248_ _01169_ _00705_ _04271_ _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_23_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09179_ cpu.ROM_addr_buff\[12\] _04185_ _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07776__A1 _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput55 net55 io_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput66 net66 io_out[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_output72_I net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput44 net44 io_oeb[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput77 net77 io_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput88 net88 sram_addr[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10023_ _02027_ _02450_ _02445_ _04966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_53_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08815__C _03920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05314__I0 cpu.regs\[8\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05900_ _01205_ _01383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06880_ _02042_ _02354_ _02355_ _02356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05831_ _01314_ _01315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06742__A2 _00933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05762_ _01102_ _01246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08550_ cpu.toggle_top\[14\] _03714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08481_ cpu.orig_PC\[7\] _03659_ _03662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05693_ _01097_ _01177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07501_ _02899_ _02900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07432_ _02842_ _02843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_81_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09102_ _00727_ _04150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_61_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07363_ _02054_ _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06314_ _01378_ _01791_ _01792_ _01793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_07294_ _02651_ _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09033_ _04084_ _04096_ _00433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06245_ _00596_ _00985_ _01725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__05481__A2 _00967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06176_ _01650_ _01656_ _01657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05127_ cpu.IO_addr_buff\[1\] _00644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09211__A4 _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09935_ cpu.PORTB_DDR\[1\] _04892_ _04896_ _04897_ _04898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_5_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06430__A1 _01435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05058_ _00002_ _00579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09866_ _04027_ _04845_ _04846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08817_ _03921_ _03916_ _03922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09797_ _02489_ _04790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09291__C _04313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08748_ _01042_ _02730_ _03864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08679_ _02746_ _03811_ _03815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06497__A1 _01441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10641_ _00535_ clknet_leaf_69_wb_clk_i cpu.PORTB_DDR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10572_ _00466_ clknet_leaf_80_wb_clk_i cpu.last_addr\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10138__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06421__A1 _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10006_ _00665_ _04952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10108__I0 _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09657__B _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06030_ cpu.timer_div\[2\] _01397_ _01509_ _01511_ _01182_ _01512_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_42_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07981_ _03181_ _03261_ _03184_ _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05215__A2 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06412__A1 _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09720_ _04723_ _04725_ _04726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06932_ _02019_ _02405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08165__A1 _03335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07912__A1 _03207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09651_ cpu.orig_PC\[13\] _04074_ _04662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06715__A2 _00907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06863_ _00634_ _00999_ _02339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_38_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09582_ _04593_ _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08602_ _03751_ _03761_ _00337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05814_ cpu.base_address\[1\] _01298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_06794_ _00805_ _02270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05745_ cpu.spi.dout\[0\] _01187_ _01191_ _01228_ _01229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08533_ _03698_ _00331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_18_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08464_ _03649_ _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05676_ _01159_ _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08395_ _02850_ _03597_ _03598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07415_ _02823_ cpu.uart.receive_div_counter\[9\] _02824_ _02825_ _02826_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_57_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07346_ cpu.PC\[0\] _02765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_116_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07277_ _00776_ _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09016_ _01077_ _04067_ _04080_ _04082_ _04083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06100__B1 _01581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06228_ _01612_ _01707_ _01708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06159_ _01301_ _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05386__I _00875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09918_ _04861_ _04885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_69_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08156__A1 _03333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07815__B _03112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09849_ cpu.pwm_top\[2\] _04831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_output35_I net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10624_ _00518_ clknet_leaf_67_wb_clk_i net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08092__B1 _03335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10555_ _00449_ clknet_leaf_80_wb_clk_i cpu.ROM_addr_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10486_ _00381_ clknet_leaf_26_wb_clk_i cpu.timer\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07690__I0 _03006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_14_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05056__S1 _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09647__A1 _03674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07122__A2 _02583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05530_ _01013_ _01014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_43_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05461_ _00940_ _00943_ _00948_ _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_08180_ _03401_ _03427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07200_ cpu.uart.divisor\[6\] _02623_ _02648_ _02640_ _02649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_43_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05392_ _00881_ _00882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_27_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07131_ _02508_ _02592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07062_ net1 _02361_ _02351_ _02529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_30_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06013_ net81 _01074_ _00677_ _01494_ _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_2_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_103_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07964_ _03251_ _03252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09703_ _04712_ _00487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07895_ _03180_ cpu.spi.divisor\[2\] _03188_ cpu.spi.div_counter\[5\] _03192_ _03193_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_06915_ _00604_ _02389_ _02363_ _02390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_69_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09634_ _04623_ _04296_ _04628_ _04645_ _04646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06846_ _02242_ _02264_ _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06777_ _00817_ _02253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09565_ cpu.PC\[9\] _00844_ _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05728_ cpu.PORTB_DDR\[0\] _01211_ _01212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_81_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08516_ _02752_ _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09496_ _04347_ _04512_ _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08447_ _03635_ _03618_ _03637_ _03620_ _00306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05659_ _01142_ _01143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_37_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05675__A2 _01158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08378_ _03580_ _03584_ _00290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09110__I0 cpu.regs\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08074__B1 _03337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07329_ _02754_ _00071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_104_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10340_ _00235_ clknet_leaf_61_wb_clk_i cpu.spi.counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10271_ _00166_ clknet_leaf_117_wb_clk_i cpu.regs\[5\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09877__A1 _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09629__A1 _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_48_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_48_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_83_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06863__A1 _00634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10607_ _00501_ clknet_leaf_73_wb_clk_i cpu.ROM_spi_dat_out\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10538_ _00432_ clknet_leaf_18_wb_clk_i cpu.IO_addr_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10469_ _00364_ clknet_leaf_19_wb_clk_i cpu.pwm_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07591__A2 _01145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06700_ _02129_ _02132_ _02176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07680_ cpu.regs\[5\]\[1\] _03012_ _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06631_ _02063_ _02064_ _02107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06562_ _02036_ _02037_ _02038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_87_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_86_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09350_ _02796_ _04369_ _04371_ _04372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08301_ _03525_ _03526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09281_ _00762_ _04299_ _04304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05513_ _00998_ _00999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_19_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08232_ _03468_ _03469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05657__A2 _00929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06493_ _01959_ _01961_ _01969_ _01970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05444_ _00931_ _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08163_ cpu.uart.div_counter\[6\] _03413_ _03414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05375_ _00858_ _00865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08094_ _03331_ _03357_ _03358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_43_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06606__A1 _00590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07114_ _02013_ _02577_ _02521_ _02578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_113_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07045_ _02512_ _02513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10056__B _04226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08996_ _00755_ _04062_ _04063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07947_ _03235_ _03237_ _03238_ _00205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_89_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08975__I _02692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07878_ _02620_ _03176_ cpu.needs_timer_interrupt _03177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09617_ cpu.orig_PC\[12\] _04239_ _04629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06829_ _02287_ _02304_ _02305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09548_ _04057_ _04554_ _04562_ _04432_ _04563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_66_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09479_ _02559_ _04297_ _04497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_54_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10323_ _00218_ clknet_leaf_48_wb_clk_i cpu.spi.data_in_buff\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10254_ _00149_ clknet_leaf_118_wb_clk_i cpu.regs\[7\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10185_ _00080_ clknet_leaf_103_wb_clk_i cpu.regs\[1\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08770__A1 cpu.timer_capture\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05431__S1 _00860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05160_ _00675_ _00676_ _00677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_24_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07261__A1 cpu.timer_capture\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09250__A2 _04273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05091_ _00567_ _00608_ _00610_ _00611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_0_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07013__A1 cpu.ROM_addr_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08850_ _03944_ _03949_ _03950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07801_ _01392_ _03102_ _03106_ _00191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05484__I _00970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08781_ _02691_ _03836_ _03858_ _03891_ _03881_ _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05993_ net27 _01425_ _01476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07732_ cpu.regs\[3\]\[7\] _03034_ _03044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07663_ _01771_ _03002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09402_ _04418_ _04420_ _04421_ _04422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06614_ _02088_ _02089_ _02086_ _02090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__07204__I _02651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09333_ _04313_ _04355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07594_ _02960_ _02961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_23_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06545_ _02019_ _02020_ _02021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09264_ _04287_ _04288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06476_ _01944_ _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08215_ _03452_ _03453_ _03454_ _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09195_ _04102_ _04221_ _00470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05427_ _00863_ _00915_ _00867_ _00916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_105_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08146_ _02813_ _03399_ _03400_ _00242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09241__A2 _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05358_ _00712_ _00848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08077_ cpu.uart.div_counter\[2\] _03341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05289_ _00799_ _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_07028_ net1 _02498_ _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_87_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08979_ _02698_ _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_59_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10306_ _00201_ clknet_leaf_57_wb_clk_i cpu.spi.data_out_buff\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08991__A1 _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10237_ _00132_ clknet_leaf_2_wb_clk_i cpu.regs\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08743__A1 _01395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05101__S0 _00615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10168_ _00067_ clknet_leaf_12_wb_clk_i cpu.toggle_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_89_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10099_ _01359_ _05035_ _05037_ _00558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_63_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_63_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_89_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06330_ cpu.pwm_top\[5\] _01619_ _01408_ _01809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09471__A2 _04359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06261_ _01134_ net93 _01741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08000_ _03190_ _03280_ _03281_ _03282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05212_ net71 _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06192_ _01574_ _01672_ _01673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05143_ cpu.ROM_spi_cycle\[3\] cpu.ROM_spi_cycle\[2\] _00660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_114_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07908__B net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08982__A1 cpu.uart.divisor\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09951_ _04909_ _00538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05074_ _00585_ _00594_ _00595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_110_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08902_ _03982_ _03990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09882_ _04041_ _04857_ _04858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08734__A1 _02643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08833_ _03933_ _03934_ _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08764_ _03860_ _03876_ _03877_ _03878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05976_ _01454_ _00901_ _01459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_56_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07715_ _03033_ _03034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08695_ _03826_ _03827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07646_ _02942_ cpu.regs\[7\]\[6\] _02978_ _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07577_ _02918_ _02947_ _02950_ _00123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_36_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06528_ _01264_ _01979_ _01717_ _02005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09316_ cpu.PC\[2\] cpu.br_rel_dest\[2\] _04338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_91_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09247_ cpu.Z _00705_ _04271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06459_ _01936_ _00019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09178_ _04201_ _04206_ _04207_ _00467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_102_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08129_ _00722_ _01395_ _03209_ _00756_ _03386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_31_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput34 net34 io_oeb[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput67 net67 io_out[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput56 net56 io_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_101_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput45 net45 io_oeb[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_12_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput78 net78 io_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_output65_I net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput89 net89 sram_gwe vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__08725__A1 _02627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10022_ net78 _04965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_113_Right_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_110_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_110_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_117_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06019__A2 _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07767__A2 _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_9_0_wb_clk_i clknet_0_wb_clk_i clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08716__A1 _01090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06858__I _00590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05830_ _01155_ _01313_ _01314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05761_ _01238_ _01245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07500_ _02898_ _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05950__A1 _01426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08480_ _02570_ _03657_ _03661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05692_ cpu.toggle_top\[0\] _01176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_49_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07431_ cpu.uart.divisor\[12\] _02842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_18_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07362_ _02526_ _02777_ _02779_ _02546_ _02780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_33_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06313_ net64 _01213_ _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09101_ _04149_ _00448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_61_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07293_ _02647_ _02719_ _02725_ _02724_ _00064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06258__A2 _00977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09032_ _00674_ _04067_ _04095_ _04082_ _04096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06244_ _00596_ _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06175_ _01531_ _00936_ _01563_ _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05126_ _00643_ net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_13_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09934_ _04861_ _04897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05057_ cpu.regs\[8\]\[4\] cpu.regs\[9\]\[4\] cpu.regs\[10\]\[4\] cpu.regs\[11\]\[4\]
+ _00572_ _00576_ _00578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09865_ _04843_ _04845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_59_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08816_ cpu.timer\[11\] _03921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09380__A1 _02052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09796_ _04789_ _00503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06194__A1 _01315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09132__A1 cpu.ROM_addr_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08747_ cpu.timer\[0\] _03858_ _03860_ _03862_ _03863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05959_ net90 _01340_ _01442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08678_ _03800_ _03814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07629_ _02979_ _02980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10640_ _00534_ clknet_leaf_69_wb_clk_i cpu.PORTB_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_101_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10571_ _00465_ clknet_leaf_80_wb_clk_i cpu.last_addr\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_75_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09199__A1 _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_98_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08946__A1 _02638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09319__I _04273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06452__B _01929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_2_Left_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_39_Left_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06421__A2 _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10005_ cpu.ROM_addr_buff\[0\] _04950_ _02483_ cpu.ROM_addr_buff\[4\] cpu.ROM_addr_buff\[8\]
+ _02484_ _04951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__07921__A2 _03195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_48_Left_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07302__I _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_57_Left_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_10_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07980_ _03184_ _03103_ _03214_ _03264_ _03203_ _03265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_10_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06931_ _02402_ _02403_ _02404_ _00023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09650_ _04656_ _04657_ _04660_ _04661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_38_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_66_Left_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08601_ cpu.toggle_ctr\[4\] _03760_ _03761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06862_ _02077_ _02078_ _02075_ _02338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05923__A1 cpu.timer_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09581_ _04594_ _04577_ _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06793_ _00899_ _02267_ _02268_ _02269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_05813_ _01296_ _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_38_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05744_ _01192_ _01226_ _01227_ _01228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08532_ cpu.toggle_top\[6\] _03690_ _03696_ _03697_ _03698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08463_ _00685_ _03649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07414_ cpu.uart.divisor\[2\] _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_18_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05675_ _01132_ _01158_ _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08394_ _03542_ _03596_ _03597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_57_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07345_ _02542_ _02764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_92_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_75_Left_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07276_ cpu.timer_top\[1\] _02712_ _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06227_ cpu.timer_div\[4\] _01183_ _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08471__C _03653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09015_ _04081_ _04082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08043__I _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06158_ _01637_ _01638_ _01639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05109_ _00614_ _00622_ _00627_ _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__07600__A1 _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06089_ _01455_ _01471_ _01571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09917_ _04045_ _04881_ _04884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09848_ _04824_ _04825_ _04828_ _04829_ _04830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__06167__A1 _01426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09779_ _02479_ _04774_ _04775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05142__A2 _00653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10623_ _00517_ clknet_leaf_67_wb_clk_i net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_36_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10554_ _00448_ clknet_leaf_83_wb_clk_i cpu.ROM_addr_buff\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10485_ _00380_ clknet_leaf_10_wb_clk_i cpu.timer_top\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_114_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05453__I0 cpu.regs\[12\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09647__A2 _00763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05460_ _00940_ _00945_ _00947_ _00948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_55_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05391_ _00855_ _00881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_70_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07130_ _02590_ _02587_ _02591_ _02589_ _00035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_40_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07061_ _02314_ net120 _02528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06012_ _01044_ _01041_ _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_2_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09583__A1 _00818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06397__A1 cpu.uart.divisor\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07963_ _03100_ _03211_ _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09702_ _04670_ _04673_ _04711_ _04124_ _04712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07894_ _03183_ cpu.spi.divisor\[3\] _03189_ _03190_ _03191_ _03192_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__06149__A1 _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06914_ _02365_ _02388_ _02022_ _02389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06111__I cpu.uart.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09633_ _02513_ _04626_ _04644_ _04227_ _04645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_4_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06845_ _02305_ _02319_ _02320_ _02321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_09564_ cpu.PC\[10\] _00929_ _04578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08515_ _02739_ _03680_ _03685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06776_ _02249_ _02251_ _02252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05727_ _01210_ _01211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09495_ _02606_ _04349_ _04511_ _04355_ _04512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_19_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08446_ cpu.orig_flags\[1\] _03636_ _03637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05658_ _00843_ _00848_ _01142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08377_ cpu.uart.receive_div_counter\[10\] _03518_ _03583_ _03584_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_83_Left_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09110__I1 _03664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05589_ _01070_ _01072_ _01073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07328_ cpu.toggle_top\[13\] _02745_ _02751_ _02753_ _02754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08074__A1 _02816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07259_ _02697_ _02686_ _02699_ _02700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10270_ _00165_ clknet_leaf_111_wb_clk_i cpu.regs\[5\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08377__A2 _03518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_92_Left_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08129__A2 _01395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07117__I _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05899__B1 _01379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05860__I _00712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06312__A1 cpu.PORTB_DDR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06863__A2 _00999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10606_ _00500_ clknet_leaf_73_wb_clk_i cpu.spi_clkdiv vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_88_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_88_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10537_ _00431_ clknet_leaf_55_wb_clk_i cpu.IO_addr_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_17_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_17_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10468_ _00363_ clknet_leaf_10_wb_clk_i cpu.pwm_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10399_ _00294_ clknet_leaf_38_wb_clk_i cpu.uart.receive_div_counter\[14\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07040__A2 _02508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07879__A1 _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07027__I _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06630_ _02103_ _02104_ _02106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08286__C _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06561_ cpu.mem_cycle\[2\] _02037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_86_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08300_ _03515_ _03524_ _03525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_87_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09280_ _04277_ _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06303__A1 _00982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05512_ _00997_ _00998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06492_ _01439_ _01949_ _01963_ _01321_ _01968_ _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08231_ _03464_ _03468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05443_ _00930_ _00931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07697__I _03021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08162_ cpu.uart.div_counter\[5\] cpu.uart.div_counter\[4\] _03406_ _03413_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_7_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05374_ _00854_ _00864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07103__I0 _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08093_ _03332_ _03334_ _03353_ _03356_ _03357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_15_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07113_ _02524_ _02572_ _02576_ _02577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07044_ _02511_ _02512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06106__I _01586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09556__A1 _00806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09417__I _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08995_ _00703_ _01110_ _04062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07946_ cpu.spi.data_out_buff\[3\] _03223_ _03228_ _03238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input27_I sram_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07877_ _03131_ _03175_ _03176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09616_ _04594_ _04626_ _04627_ _04413_ _04628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06828_ _02297_ _02303_ _02304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05680__I _01106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09547_ _03664_ _04351_ _04562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06759_ _02207_ _02208_ _02235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_93_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09478_ _04328_ _04492_ _04495_ _04496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08429_ _00670_ _03624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_4_11_0_wb_clk_i clknet_0_wb_clk_i clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_80_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10322_ _00217_ clknet_leaf_48_wb_clk_i cpu.spi.data_in_buff\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output95_I net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07270__A2 _02610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09547__A1 _03664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10253_ _00148_ clknet_leaf_110_wb_clk_i cpu.regs\[7\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07275__C _00778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10184_ _00079_ clknet_leaf_107_wb_clk_i cpu.regs\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05590__I _00671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06533__A1 _01115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07310__I _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05090_ _00583_ _00609_ _00610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07800_ cpu.spi.data_in_buff\[1\] _03104_ _03105_ _03106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08780_ _02691_ _03884_ _03891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07731_ _03043_ _00184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05992_ _01297_ net91 _01474_ _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__09710__A1 _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07662_ _02987_ _02996_ _03001_ _00157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09401_ _02767_ _02056_ _04421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06613_ _00830_ _01955_ _02089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07593_ _02959_ _02912_ _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09332_ _04350_ _04331_ _04352_ _04353_ _04354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06544_ _01137_ _01157_ _02020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_87_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09263_ _01298_ _01002_ _01528_ _04287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06475_ _01940_ _01951_ _01952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08214_ _03359_ _03454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09194_ cpu.TIE _04216_ _04217_ _04220_ _04221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09077__I0 _00806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05426_ cpu.regs\[4\]\[2\] cpu.regs\[5\]\[2\] cpu.regs\[6\]\[2\] cpu.regs\[7\]\[2\]
+ _00856_ _00860_ _00915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_08145_ _03348_ _03350_ _03341_ _03400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05357_ _00846_ _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_102_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08076_ cpu.uart.div_counter\[7\] _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_05288_ _00793_ _00798_ _00799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_07027_ _00729_ _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08201__A1 _03383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08978_ _04047_ _00427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07929_ cpu.spi.data_out_buff\[0\] _03223_ _03112_ _03224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_59_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05624__B _01107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10075__A1 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06455__B _01932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08226__I _03386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_20_Left_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10305_ _00200_ clknet_leaf_49_wb_clk_i cpu.spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__08991__A2 _01734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05585__I _01068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10236_ _00131_ clknet_leaf_2_wb_clk_i cpu.regs\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09940__A1 _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10167_ _00066_ clknet_leaf_12_wb_clk_i cpu.toggle_top\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10098_ cpu.regs\[15\]\[0\] _05036_ _05037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06506__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07305__I _00903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08259__A1 _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_32_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_32_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_84_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06260_ _01655_ _01739_ _01740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09759__A1 _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05211_ _00694_ _00721_ _00725_ _00726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05493__A1 _00928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06191_ _01660_ _01670_ _01672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05142_ _00650_ _00653_ _00656_ _00658_ _00659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_40_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09950_ cpu.PORTB_DDR\[5\] _04903_ _04907_ _04908_ _04909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05073_ _00587_ _00592_ _00593_ _00594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_49_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08901_ _03982_ _03989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09881_ _04843_ _04857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09931__A1 cpu.PORTB_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08832_ _03929_ _03924_ _03934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08763_ _02667_ _03862_ _02673_ _03877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05975_ net91 _00907_ _01458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08498__A1 _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07714_ _02020_ _02929_ _03033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08694_ _02619_ _03825_ _03826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07645_ _02990_ _00151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_0_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07576_ cpu.regs\[10\]\[1\] _02948_ _02950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_36_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06527_ cpu.toggle_top\[15\] _01257_ _01979_ _02003_ _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09315_ _04335_ _04310_ _04336_ _04337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_106_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09246_ _00706_ _00765_ _04270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06458_ _01935_ cpu.regs\[9\]\[6\] _01159_ _01936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05409_ _00892_ _00898_ _00899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06389_ cpu.PORTA_DDR\[6\] net57 _01207_ _01867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09177_ cpu.last_addr\[11\] _04176_ _04207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_88_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09586__B _04523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08128_ _03345_ _03384_ _03385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08059_ cpu.uart.div_counter\[12\] _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05236__A1 _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput57 net57 io_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput46 net46 io_oeb[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput35 net35 io_oeb[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput79 net79 io_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput68 net68 io_out[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10021_ _00778_ _04964_ _00553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_8_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09922__A1 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output58_I net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05314__I2 cpu.regs\[10\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05227__A1 _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05529__B _01012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10219_ _00114_ clknet_leaf_4_wb_clk_i cpu.regs\[11\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05760_ cpu.timer_capture\[8\] _01243_ _01244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_89_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07152__A1 _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05691_ _01174_ _01175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07430_ cpu.uart.receive_div_counter\[4\] cpu.uart.divisor\[4\] _02841_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07361_ _02778_ _01003_ _02668_ _02772_ _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_122_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06312_ cpu.PORTB_DDR\[5\] _01595_ _01790_ _01121_ _01791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_09100_ _04146_ _04147_ _04148_ _04149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07292_ cpu.timer_top\[6\] _02720_ _02725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09031_ _01587_ _04070_ _04072_ _04093_ _04094_ _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_45_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06243_ _01683_ _01164_ _01720_ _01722_ _01723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_115_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08404__A1 _03514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06174_ _01447_ _01655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05218__A1 _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_5_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05125_ _00642_ _00643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09933_ _04031_ _04893_ _04896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06114__I _01091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05056_ cpu.regs\[12\]\[4\] cpu.regs\[13\]\[4\] cpu.regs\[14\]\[4\] cpu.regs\[15\]\[4\]
+ _00572_ _00576_ _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09864_ _04843_ _04844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06718__A1 _00590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08469__C _03653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08815_ _01486_ _03866_ _03919_ _03920_ _00391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09380__A2 _04068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09795_ cpu.ROM_spi_dat_out\[2\] _04778_ _04787_ _04788_ _04789_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08746_ cpu.timer\[0\] _03861_ _03862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05958_ _01347_ _01441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05889_ _01371_ _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08677_ _03813_ _00360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07628_ _02978_ _02979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07559_ _01771_ _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_101_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10570_ _00464_ clknet_leaf_80_wb_clk_i cpu.last_addr\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08643__A1 _03514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09229_ _02334_ _02370_ _02373_ _02375_ _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_17_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09763__C _03474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_112_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10004_ _02025_ _04670_ _02445_ _02446_ _04950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XPHY_EDGE_ROW_73_Right_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07283__C _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06185__A2 _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_103_Left_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07134__A1 _02592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07685__A2 _03011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_80_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_82_Right_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_30_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_112_Left_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_91_Right_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05620__A1 _01100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06930_ _01934_ _02023_ _02363_ cpu.regs\[2\]\[6\] _02404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_38_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I io_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05773__I _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07748__I0 _00790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08600_ cpu.toggle_ctr\[3\] _03757_ _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06861_ _00603_ _01288_ _02337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07373__A1 _02789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09580_ _04593_ _04594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06792_ _00830_ _00877_ _02268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05812_ _00654_ _01296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_38_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05743_ cpu.uart.busy _01079_ _01076_ _01227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08531_ _02752_ _03697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07125__A1 _01111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08462_ cpu.orig_PC\[2\] _03643_ _03648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05674_ _01138_ _01157_ _01158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_07413_ cpu.uart.receive_div_counter\[2\] _02824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08873__A1 cpu.timer_capture\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08393_ _02850_ _03593_ _03539_ _03596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07344_ _02595_ _02760_ _02596_ _02763_ _00077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_73_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07275_ _02708_ _02711_ _02713_ _00778_ _00058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_61_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06226_ _01691_ _01608_ _01704_ _01705_ _01183_ _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_09014_ _02609_ _04081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_61_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09050__B2 _01291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06157_ _01532_ _01537_ _01534_ _01638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__06939__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05108_ _00614_ _00624_ _00626_ _00627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06088_ _01560_ _01568_ _01326_ _01570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09916_ _04883_ _00529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09847_ cpu.pwm_top\[5\] cpu.pwm_counter\[5\] _04829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09778_ _04765_ _04773_ _04774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08729_ _03840_ _03849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07403__I cpu.uart.divisor\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05142__A3 _00656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10622_ _00516_ clknet_leaf_88_wb_clk_i net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_63_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10553_ _00447_ clknet_leaf_83_wb_clk_i cpu.ROM_addr_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10484_ _00379_ clknet_leaf_23_wb_clk_i cpu.timer_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09041__B2 _00999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05390_ _00852_ _00880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_82_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07060_ _02314_ net120 _02527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06011_ _01027_ _01030_ _01046_ cpu.PORTA_DDR\[2\] _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_42_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05841__A1 _00970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09701_ _04672_ _04675_ _04710_ _04711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07962_ cpu.spi.div_counter\[0\] _03250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07893_ cpu.spi.div_counter\[1\] _03187_ _03189_ cpu.spi.div_counter\[6\] _03191_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06913_ _02042_ _02386_ _02387_ _02388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09632_ _04327_ _04643_ _04644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06844_ _02266_ _02284_ _02320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_09563_ _04576_ _04577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08514_ _03684_ _00326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06775_ _02244_ _02245_ _02250_ _02251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05726_ _01026_ _01029_ _01101_ _01210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_65_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09494_ _04350_ _04501_ _04510_ _04353_ _04511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09859__B net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08445_ _03608_ _03636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05657_ _00969_ _00929_ _01141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08376_ _03570_ _03581_ _03582_ _03583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_108_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05588_ _00702_ _00717_ _00755_ _01071_ _01072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_61_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07327_ _02752_ _02753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_6_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07258_ _02680_ _02698_ _02699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07189_ _02639_ _02640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06209_ cpu.timer_top\[4\] _01689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09023__B2 _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07888__A2 cpu.spi.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output40_I net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09637__I0 _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10605_ _00499_ clknet_leaf_78_wb_clk_i cpu.startup_cycle\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09262__A1 _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06076__A1 _01336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10536_ _00430_ clknet_leaf_18_wb_clk_i cpu.IO_addr_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_108_Right_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10467_ _00362_ clknet_leaf_15_wb_clk_i cpu.pwm_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_75_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09565__A2 _00844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10398_ _00293_ clknet_leaf_36_wb_clk_i cpu.uart.receive_div_counter\[13\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_57_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_57_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07576__A1 cpu.regs\[10\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06212__I cpu.uart.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07328__A1 cpu.toggle_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06000__A1 cpu.regs\[9\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06560_ _02035_ _02036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_59_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05511_ _00996_ _00997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06491_ _01457_ _01943_ _01964_ _01967_ _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_08230_ _03365_ _03467_ _00259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_51_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05442_ _00929_ _00930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06303__A2 _01781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08161_ _03402_ _03412_ _00245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_70_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05373_ _00006_ _00863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08092_ _02842_ _03354_ _03335_ _02815_ _03355_ _03356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_43_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07112_ _02392_ _02574_ _02575_ _02534_ _02576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07043_ _00707_ _02511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08994_ _04060_ _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07945_ cpu.spi.data_out_buff\[4\] _03230_ _03236_ _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07876_ _03174_ _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09615_ _00591_ _04596_ _04627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06827_ _02297_ _02298_ _02302_ _02303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_78_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08819__A1 _01591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09546_ _04334_ _04554_ _04560_ _04345_ _04561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_06758_ _02231_ _02232_ _02233_ _02234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05709_ _00681_ _01193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09477_ _04368_ _04474_ _04494_ _04374_ _04375_ _04495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_109_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08428_ cpu.IO_addr_buff\[5\] _03622_ _03623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09492__A1 _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06689_ _02163_ _02164_ _02165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_93_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08359_ _03568_ _03569_ _00286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_80_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09095__I1 cpu.ROM_addr_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10321_ _00216_ clknet_leaf_49_wb_clk_i cpu.spi.div_counter\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10252_ _00147_ clknet_leaf_13_wb_clk_i cpu.regs\[7\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10183_ _00078_ clknet_leaf_107_wb_clk_i cpu.regs\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06230__A1 cpu.timer_capture\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07128__I _02505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05584__A3 _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07291__C _02724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10519_ _00414_ clknet_leaf_30_wb_clk_i cpu.timer_div\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_39_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08422__I _03609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07730_ _03006_ cpu.regs\[3\]\[6\] _03033_ _03043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05991_ _01434_ _01437_ _01464_ _01473_ _01474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_88_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07661_ cpu.regs\[6\]\[3\] _02995_ _03001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07721__A1 _01481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06612_ _02086_ _02087_ _02088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07592_ _01137_ _02958_ _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09400_ _02802_ _04384_ _04420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09331_ _04303_ _04353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06543_ _02018_ _01130_ _02019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06288__A1 _01012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09262_ _00758_ _04283_ _04285_ _04286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06474_ _01941_ _01947_ _01950_ _01951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_clkbuf_leaf_78_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08213_ _00724_ _01395_ _03209_ _00758_ _03453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_09193_ _03231_ _04218_ _04219_ _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09077__I1 _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05425_ _00853_ _00913_ _00914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_99_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08144_ _03341_ _03388_ _03397_ _03398_ _03399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_16_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07088__I0 _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05356_ _00845_ _00846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08075_ _02814_ cpu.uart.div_counter\[13\] _03335_ _02815_ _03338_ _03339_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__05956__I _01438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05287_ _00003_ _00795_ _00797_ _00798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_07026_ _02495_ _02497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08977_ cpu.uart.divisor\[13\] _04040_ _04046_ _04035_ _04047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xclkbuf_leaf_2_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_2_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07928_ _03217_ _03223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07859_ _03155_ _03156_ _03157_ _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_3_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05624__C _00844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09529_ _04410_ _04527_ _04545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09465__A1 _04456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06279__A1 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08507__I _03678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10075__A2 _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09217__A1 _01587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10304_ _00199_ clknet_leaf_48_wb_clk_i net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_72_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10235_ _00130_ clknet_leaf_109_wb_clk_i cpu.regs\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08398__B _03600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10166_ _00065_ clknet_leaf_22_wb_clk_i cpu.timer_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10097_ _05033_ _05036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_88_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_112_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10066__A2 _04213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09208__A1 _01854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05210_ _00724_ _00725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05493__A2 _00951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06690__A1 cpu.regs\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06190_ _01660_ _01670_ _01671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_72_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_72_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_106_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05141_ _00657_ cpu.br_rel_dest\[6\] cpu.br_rel_dest\[4\] _00658_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_80_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05245__A2 _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05072_ _00003_ _00593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_09880_ _04843_ _04856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_94_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08900_ _02631_ _03983_ _03988_ _00408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08831_ cpu.timer\[14\] _03933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08762_ _03174_ _03875_ _03861_ _03876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05974_ _01143_ _01334_ _01457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08693_ _03131_ _03825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07713_ _02992_ _03024_ _03032_ _00177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07644_ _02940_ cpu.regs\[7\]\[5\] _02978_ _02990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_0_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07575_ _02910_ _02947_ _02949_ _00122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_36_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09998__A2 _00692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06526_ _02000_ _02001_ _02002_ _01625_ _02003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09314_ _02054_ cpu.br_rel_dest\[1\] _04336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09245_ cpu.orig_PC\[0\] _04267_ _04268_ _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06457_ _01934_ _01935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05408_ _00894_ _00897_ _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06388_ cpu.uart.divisor\[6\] _01866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_09176_ cpu.ROM_addr_buff\[11\] _04194_ _04206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08127_ _03383_ _03384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05339_ cpu.PORTB_DDR\[5\] net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__05686__I _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08058_ net68 _03322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput58 net58 io_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_07009_ _02470_ _02481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput47 net47 io_oeb[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput36 net36 io_oeb[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_31_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput69 net69 io_out[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10020_ net76 _04945_ _04947_ _04963_ _04964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_8_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06197__B1 _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07406__I cpu.uart.receive_div_counter\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08237__I _02619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05797__S _00852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05314__I3 cpu.regs\[11\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07924__A1 _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10218_ _00113_ clknet_leaf_126_wb_clk_i cpu.regs\[12\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10149_ _00048_ clknet_leaf_31_wb_clk_i cpu.uart.divisor\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06220__I _01195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05690_ _01100_ _01174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05163__A1 _00671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09429__A1 _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08147__I _02872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07360_ _02270_ _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08101__A1 _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06311_ net36 _01593_ _01789_ _01595_ _01790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_61_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07291_ _02643_ _02719_ _02722_ _02724_ _00063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09030_ _04078_ _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06242_ _00951_ _01278_ _01721_ _01722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06663__A1 _00619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06890__I _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06173_ _01451_ _01651_ _01646_ _01439_ _01653_ _01654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__06415__A1 _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05124_ _00614_ _00636_ _00641_ _00642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_110_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09932_ _04895_ _00533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05055_ _00575_ _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09863_ _01067_ _04842_ _04843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_5_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09794_ _04123_ _04788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_99_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08814_ _02761_ _03920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08745_ _03855_ _03861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05957_ _01439_ _01440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05888_ _01203_ _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08676_ cpu.pwm_top\[3\] _03801_ _03812_ _03809_ _03813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07627_ _02929_ _02977_ _02978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_64_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07558_ _02922_ _02932_ _02937_ _00117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06509_ net67 _01070_ _01216_ _01986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09840__A1 _03207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07489_ cpu.regs\[14\]\[3\] _02887_ _02893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09228_ _04252_ _04253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09159_ _04171_ _04194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06305__I _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output70_I net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08159__A1 _03337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10003_ cpu.ROM_addr_buff\[12\] _02465_ _04948_ _04949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07906__A1 _03201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08331__A1 _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09831__A1 _03288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06860_ _02333_ _02335_ _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05811_ _01170_ _01171_ _01173_ _01294_ _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_54_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06791_ _00805_ _00934_ _02267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_38_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05742_ _01194_ _01222_ _01225_ _01226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_54_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08530_ _02755_ _03691_ _03696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06885__I _02360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08461_ _02789_ _03641_ _03647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05673_ _01139_ _01145_ _01156_ _01157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_07412_ _02816_ _02823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_18_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08392_ _03580_ _03595_ _00293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07710__S _03021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07343_ _02592_ _02760_ _02594_ _02763_ _00076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_07274_ cpu.timer_top\[0\] _02712_ _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09210__B _00711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06225_ cpu.spi.divisor\[4\] _01606_ _01190_ _01705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_72_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09013_ _01163_ _04070_ _04072_ _04077_ _04079_ _04080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_14_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09637__S _04500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06125__I _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06156_ _01635_ _01636_ _01637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05107_ _00621_ _00625_ _00626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05964__I _01446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06087_ _01559_ _01568_ _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09915_ net55 _04880_ _04882_ _04874_ _04883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05611__A2 _01094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09846_ cpu.pwm_top\[1\] _04826_ _03782_ _04827_ _04828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_09777_ _04767_ _04773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06989_ _02448_ _02461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08728_ _03840_ _03848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08659_ _03781_ _03799_ _00356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_83_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09113__I0 cpu.regs\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07620__S _02963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10621_ _00515_ clknet_leaf_17_wb_clk_i net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_48_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10552_ _00446_ clknet_leaf_83_wb_clk_i cpu.ROM_addr_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_63_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10483_ _00378_ clknet_leaf_10_wb_clk_i cpu.timer_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_114_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05850__A2 _00715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09081__I _04022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05508__I3 cpu.regs\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_43_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07291__A1 _02643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06010_ net23 _01492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_23_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05841__A2 _00930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07961_ _03235_ _03248_ _03249_ _00208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09700_ _04709_ _04710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06912_ net12 _02041_ _02387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07892_ cpu.spi.div_counter\[6\] _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09631_ _04301_ _04626_ _04642_ _04365_ _04643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06843_ _02317_ _02318_ _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_09562_ _03070_ _04553_ _04576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06774_ _00589_ _00906_ _02250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05725_ cpu.PORTA_DDR\[0\] net79 _01208_ _01209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08513_ cpu.toggle_top\[1\] _03679_ _03683_ _03461_ _03684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09493_ _02569_ _04484_ _04510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05656_ _00652_ _00710_ _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08444_ cpu.Z _03635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08375_ _03576_ _03577_ cpu.uart.receive_div_counter\[10\] _03582_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_86_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05587_ _00649_ _00653_ _01008_ _01071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_46_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07326_ _02638_ _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07257_ _01785_ _02698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07188_ _02638_ _02639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06208_ _01687_ _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_14_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06139_ cpu.timer_top\[11\] _01118_ _01615_ _01618_ _01619_ _01620_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__08782__A1 cpu.timer_capture\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05596__A1 _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08129__A4 _00756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08534__A1 _02652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09829_ _04809_ _04807_ _04811_ _04815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_69_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05520__A1 _01002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10604_ _00498_ clknet_leaf_78_wb_clk_i cpu.startup_cycle\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05371__I1 cpu.regs\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10535_ _00429_ clknet_leaf_40_wb_clk_i cpu.uart.divisor\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10466_ _00361_ clknet_leaf_15_wb_clk_i cpu.pwm_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_29_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10397_ _00292_ clknet_leaf_36_wb_clk_i cpu.uart.receive_div_counter\[12\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_26_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_26_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08525__A1 cpu.toggle_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07324__I _02692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05510_ _00992_ _00995_ _00870_ _00996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06490_ _01450_ _01945_ _01966_ _01452_ _01967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_28_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05441_ cpu.base_address\[2\] _00929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_117_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_68_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08160_ _03337_ _03389_ _03411_ _03384_ _03412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_27_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08155__I _03383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05372_ _00861_ _00853_ _00862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07111_ net20 _02535_ _02575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08091_ cpu.uart.div_counter\[7\] _02856_ _02622_ _03349_ _03355_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_42_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07042_ _02510_ _00028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08993_ _01133_ _01146_ _00746_ _04060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_07944_ _02634_ _03225_ _03236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08758__C _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07875_ _03132_ _03173_ _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09614_ _04625_ _04626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06826_ _00907_ _02300_ _02301_ _02302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06757_ _02229_ _02230_ _02233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09545_ _04557_ _04558_ _04559_ _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05708_ _01079_ _01192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09476_ _02373_ _04369_ _04493_ _04494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06688_ _00997_ cpu.regs\[1\]\[1\] _02164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_93_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08427_ _03621_ _03622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05639_ _01086_ _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_93_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08358_ _02855_ _03566_ _03437_ _03569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08289_ cpu.uart.receiving _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_07309_ _02738_ _00067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06058__A2 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10320_ _00215_ clknet_leaf_49_wb_clk_i cpu.spi.div_counter\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10251_ _00146_ clknet_leaf_12_wb_clk_i cpu.regs\[7\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10182_ _00077_ clknet_leaf_109_wb_clk_i _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_70_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07144__I _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_102_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10518_ _00413_ clknet_leaf_21_wb_clk_i cpu.timer_div\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07319__I _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10449_ _00344_ clknet_leaf_6_wb_clk_i cpu.toggle_ctr\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05104__S0 _00615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05990_ _01467_ _01470_ _01472_ _01322_ _01473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_88_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07660_ _02985_ _02996_ _03000_ _00156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06611_ _02084_ _02085_ _02087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07591_ _02957_ _01145_ _01156_ _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09330_ _02788_ _04351_ _04352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06542_ _01109_ _02018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09261_ _00758_ _04283_ _04284_ _04285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08212_ cpu.uart.counter\[0\] _03452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06473_ _01941_ _01949_ _01950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09192_ cpu.orig_flags\[3\] _04218_ _04219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05424_ cpu.regs\[0\]\[2\] cpu.regs\[1\]\[2\] cpu.regs\[2\]\[2\] cpu.regs\[3\]\[2\]
+ _00881_ _00883_ _00913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_99_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08143_ _03383_ _03398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07237__A1 _00978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05355_ _00844_ _00845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08985__A1 _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08074_ _02816_ _03336_ _03337_ _02818_ _03338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_43_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07025_ _02495_ _02496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05286_ _00579_ _00796_ _00797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07229__I _02655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input32_I sram_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08976_ _04045_ _04042_ _04046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07927_ cpu.spi.data_out_buff\[1\] _03212_ _03221_ _03222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09162__A1 _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06289__B _01478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07858_ cpu.timer_top\[3\] _02679_ _02672_ cpu.timer_top\[2\] _03157_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_07789_ cpu.spi.dout\[0\] _03095_ _03096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_97_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06809_ _02266_ _02284_ _02285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_94_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09528_ _04383_ _04527_ _04543_ _04407_ _04544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_66_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09459_ _04475_ _04476_ _04477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05212__I net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09217__A2 _02093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08976__A1 _04045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10303_ _00198_ clknet_leaf_57_wb_clk_i cpu.needs_timer_interrupt vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08523__I _03678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10234_ _00129_ clknet_leaf_126_wb_clk_i cpu.regs\[10\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10165_ _00064_ clknet_leaf_23_wb_clk_i cpu.timer_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07400__A1 _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05882__I _01364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10096_ _05034_ _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08900__A1 _02631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08967__A1 cpu.uart.divisor\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05140_ cpu.br_rel_dest\[7\] _00657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_107_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05325__S0 _00570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05071_ cpu.regs\[0\]\[4\] _00590_ _00591_ cpu.regs\[3\]\[4\] _00571_ _00575_ _00592_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_40_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_41_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_41_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_94_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07049__I _02516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08830_ _03931_ _03932_ _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08761_ _02673_ _02667_ _02657_ _03875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_05973_ _01304_ _01455_ _01456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08692_ _03822_ _03824_ _00364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07712_ cpu.regs\[4\]\[7\] _03022_ _03032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09695__A2 cpu.ROM_addr_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07643_ _02989_ _00150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05800__S1 _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07574_ cpu.regs\[10\]\[0\] _02948_ _02949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09313_ cpu.PC\[1\] cpu.br_rel_dest\[1\] _04335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06525_ cpu.toggle_top\[7\] _01252_ _02002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_36_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09244_ _02766_ _04267_ _04268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06456_ _01933_ _01934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_29_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09867__C _04788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09175_ _04204_ _04172_ _04205_ _04006_ _00466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_63_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05407_ _00887_ _00895_ _00896_ _00897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08126_ _03362_ _03363_ _03359_ _03383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__08958__A1 _04031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06387_ cpu.spi.dout\[6\] _01865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_44_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05338_ cpu.PORTA_DDR\[4\] net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08057_ _03319_ _03320_ _03321_ _00232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05269_ _00694_ _00699_ _00781_ _00782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07008_ cpu.ROM_spi_dat_out\[7\] _02479_ _02480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_101_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput48 net48 io_oeb[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_12_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput37 net37 io_oeb[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput59 net59 io_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08959_ _02816_ _04026_ _04032_ _04015_ _04033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09686__A2 cpu.ROM_addr_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09438__A2 _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07449__A1 cpu.uart.divisor\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05877__I _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07297__C _02724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10217_ _00112_ clknet_leaf_122_wb_clk_i cpu.regs\[12\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09374__A1 _02803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10148_ _00047_ clknet_leaf_31_wb_clk_i cpu.uart.divisor\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10079_ _01938_ _01965_ _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09677__A2 cpu.ROM_addr_buff\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09429__A2 _04379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08101__A2 _03364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06310_ net56 _01208_ _01789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07290_ _02723_ _02724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_33_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06241_ _01024_ _01172_ _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06172_ _01457_ _01636_ _01652_ _01653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05123_ _00614_ _00638_ _00640_ _00641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07612__A1 cpu.regs\[8\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09931_ cpu.PORTB_DDR\[0\] _04892_ _04894_ _04885_ _04895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_68_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07708__S _03021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05054_ _00574_ _00575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09862_ _00677_ _02729_ _04842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_5_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09793_ _04780_ _04786_ _04787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08813_ _03143_ _03825_ _03857_ _03918_ _03865_ _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08744_ _03859_ _03860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05956_ _01438_ _01439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05887_ _01205_ _01370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_95_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08675_ _02742_ _03811_ _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08338__I _03551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07626_ _02976_ _02977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_76_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07557_ cpu.regs\[11\]\[3\] _02931_ _02937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06508_ cpu.PORTB_DDR\[7\] _01092_ _01984_ _01122_ _01985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_101_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07488_ _01584_ _02888_ _02892_ _00092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09169__I _03201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09227_ _00740_ _01267_ _04251_ _04252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06654__A2 _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06439_ _01338_ _01784_ _01899_ _01336_ _01917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_91_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09158_ _04187_ _04191_ _04193_ _00461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08109_ _03216_ cpu.spi.counter\[1\] _03370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09089_ _04140_ _00445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07618__S _02963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09356__A1 _02789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10002_ _02445_ _02446_ _02461_ _04948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_98_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06590__A1 cpu.regs\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_17_Left_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_26_Left_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07755__C _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05810_ _01275_ _01278_ _01291_ _01292_ _01293_ _01294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_89_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06790_ _02261_ _02262_ _02266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_38_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05741_ _01223_ _01224_ _01225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08460_ _03645_ _03646_ _03633_ _00310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06333__A1 cpu.toggle_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05672_ _01146_ _01150_ _01154_ _01155_ _01156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_07411_ cpu.uart.receive_div_counter\[3\] _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_08391_ cpu.uart.receive_div_counter\[13\] _03557_ _03592_ _03594_ _03595_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_35_Left_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09122__I1 cpu.ROM_addr_buff\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07342_ _02590_ _02760_ _02591_ _02763_ _00075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_73_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07273_ _02710_ _02712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06224_ cpu.uart.dout\[4\] _01194_ _01701_ _01703_ _01080_ _01704_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_73_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09012_ _04078_ _04079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06155_ net93 _00976_ _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_4_1_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_44_Left_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05106_ cpu.regs\[8\]\[6\] cpu.regs\[9\]\[6\] cpu.regs\[10\]\[6\] cpu.regs\[11\]\[6\]
+ _00615_ _00616_ _00625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06086_ _01469_ _01561_ _01568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09914_ _04041_ _04881_ _04882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09845_ cpu.pwm_top\[0\] _04827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09776_ _04770_ _04772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06988_ _02457_ _02459_ _02460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08727_ _02631_ _03841_ _03847_ _03844_ _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05939_ cpu.Z _01171_ _01422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_53_Left_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08658_ cpu.pwm_counter\[7\] _03797_ _03799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_49_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07609_ _02910_ _02965_ _02967_ _00138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_4_8_0_wb_clk_i clknet_0_wb_clk_i clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_95_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09113__I1 _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08589_ _03751_ _03752_ _00333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10620_ _00514_ clknet_leaf_73_wb_clk_i net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07824__B2 cpu.timer_div\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10551_ _00445_ clknet_leaf_83_wb_clk_i cpu.ROM_addr_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10482_ _00377_ clknet_leaf_23_wb_clk_i cpu.timer_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_19_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_62_Left_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_114_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_71_Left_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_115_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08068__A1 cpu.uart.divisor\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_58_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05429__I0 cpu.regs\[8\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07960_ cpu.spi.data_out_buff\[6\] _03218_ _03245_ _03249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06911_ _02045_ _02367_ _02383_ _02385_ _02386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07891_ cpu.spi.divisor\[6\] _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09740__A1 _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09630_ _04630_ _04641_ _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06842_ _02304_ _02287_ _02318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09561_ _04373_ _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06773_ _00899_ _02244_ _02245_ _02249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_05724_ _01207_ _01208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08512_ _02735_ _03680_ _03683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09492_ _00767_ _04507_ _04508_ _04509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__05305__I _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08443_ _01170_ _03618_ _03634_ _03620_ _00305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05655_ _01023_ _01065_ _01073_ _01105_ _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_08374_ cpu.uart.receive_div_counter\[10\] _03576_ _03577_ _03581_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and3_1
X_05586_ _01069_ _01070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_73_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07325_ _02750_ _02747_ _02751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07256_ cpu.timer\[6\] _02697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10086__C _04327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06207_ _01686_ _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07187_ _00683_ _02638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_14_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08351__I _03517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06138_ _01126_ _01619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_14_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06069_ _01303_ _01455_ _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05596__A2 _01079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06793__A1 _00899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09828_ _04809_ _04807_ _04814_ _02762_ _00510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09759_ _03789_ _04756_ _04757_ _00498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_69_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05520__A2 _01004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10603_ _00497_ clknet_leaf_76_wb_clk_i cpu.startup_cycle\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_92_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10534_ _00428_ clknet_leaf_40_wb_clk_i cpu.uart.divisor\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10465_ _00360_ clknet_leaf_15_wb_clk_i cpu.pwm_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_20_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10396_ _00291_ clknet_leaf_36_wb_clk_i cpu.uart.receive_div_counter\[11\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_75_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05587__A2 _00653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09722__A1 _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07605__I _02963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05326__S _00581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_66_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_66_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_99_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07541__S _02913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05125__I _00642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_86_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05440_ _00713_ _00928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_55_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05061__S _00581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05371_ cpu.regs\[0\]\[0\] cpu.regs\[1\]\[0\] cpu.regs\[2\]\[0\] cpu.regs\[3\]\[0\]
+ _00856_ _00860_ _00861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07110_ _02573_ _02322_ _02574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08090_ cpu.uart.div_counter\[12\] _03354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__07264__A2 _01291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08461__A1 _02789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07041_ _00735_ _02496_ _02509_ _02503_ _02510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_42_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08213__A1 _00724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10020__B2 _04963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10020__A1 net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09961__A1 _02707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08992_ _00748_ _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07943_ _03217_ _03235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07874_ _03153_ _03154_ _03165_ _03172_ _03173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06527__A1 cpu.toggle_top\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09613_ _02062_ _04499_ _04624_ _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06825_ _02292_ _02294_ _02301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09544_ _04557_ _04558_ _04341_ _04559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06756_ _02223_ _02224_ _02232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05707_ _01188_ _01189_ _01190_ _01191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09475_ _04370_ _04474_ _04493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10087__A1 _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06687_ _00816_ _00963_ _02163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05638_ _01121_ _01122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08426_ _03607_ _03621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_108_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07250__I _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08357_ _02855_ _03557_ _03558_ _03567_ _03568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05569_ _00678_ _01051_ _01044_ _01052_ _01049_ _01053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_61_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08288_ _02812_ _03514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_73_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08452__A1 _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07308_ cpu.toggle_top\[9\] _02732_ _02736_ _02737_ _02738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_18_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07239_ cpu.timer_capture\[3\] _02656_ _02682_ _02664_ _02683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_6_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10250_ _00145_ clknet_leaf_126_wb_clk_i cpu.regs\[8\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09952__A1 _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10181_ _00076_ clknet_leaf_109_wb_clk_i _00006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08030__B _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10078__A1 _01322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07160__I _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08443__A1 _01170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10517_ _00412_ clknet_leaf_53_wb_clk_i cpu.spi.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08205__B _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10448_ _00343_ clknet_leaf_4_wb_clk_i cpu.toggle_ctr\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10379_ _00274_ clknet_leaf_45_wb_clk_i cpu.uart.receive_buff\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05280__I1 _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06509__A1 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_9_Left_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06610_ _02084_ _02085_ _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07590_ _01128_ _02957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_88_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06541_ _01770_ _02017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09260_ _00753_ _04284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06472_ _01937_ _01948_ _01949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08211_ _03301_ _03451_ _03321_ _00256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08682__A1 _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05423_ _00879_ _00910_ _00911_ _00912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_7_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09191_ _04213_ _04218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_99_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08142_ cpu.uart.div_counter\[2\] cpu.uart.div_counter\[1\] cpu.uart.div_counter\[0\]
+ _03397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_7_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05354_ _00843_ _00844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_102_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08073_ cpu.uart.div_counter\[5\] _03337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_70_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05285_ cpu.regs\[8\]\[0\] cpu.regs\[9\]\[0\] cpu.regs\[10\]\[0\] cpu.regs\[11\]\[0\]
+ _00785_ _00573_ _00796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_101_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07024_ _02493_ _02494_ _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_101_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06748__A1 _00831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08975_ _02692_ _04045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07926_ _00904_ _03214_ _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input25_I rst_n vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07173__A1 _02621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07857_ cpu.timer_top\[2\] _02673_ _02666_ cpu.timer_top\[1\] _03156_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07788_ cpu.spi.counter\[3\] cpu.spi.counter\[2\] cpu.spi.counter\[4\] _03094_ _03095_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_3_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06808_ _02275_ _02282_ _02283_ _02284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_94_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09527_ _04536_ _04540_ _04542_ _04543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06739_ _02184_ _02162_ _02215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_39_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09458_ cpu.PC\[5\] _00701_ _04459_ _04476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08009__C _03288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08409_ _03608_ _03609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_50_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09389_ _04319_ _04410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05239__A1 _00711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output93_I net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10302_ _00197_ clknet_leaf_52_wb_clk_i cpu.spi.dout\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09925__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10233_ _00128_ clknet_leaf_121_wb_clk_i cpu.regs\[10\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10164_ _00063_ clknet_leaf_22_wb_clk_i cpu.timer_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05098__S0 _00615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10095_ _05033_ _05034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09303__C _04124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05325__S1 _00827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05070_ cpu.regs\[2\]\[4\] _00591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_110_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_94_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_6_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05089__S0 _00572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_10_0_wb_clk_i clknet_0_wb_clk_i clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xclkbuf_leaf_81_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_81_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08760_ cpu.timer_capture\[2\] _03866_ _03874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05972_ _01015_ _01454_ _01455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_73_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08691_ cpu.pwm_top\[7\] _03814_ _03823_ _03824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_10_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_10_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07711_ _03031_ _00176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07642_ _02938_ cpu.regs\[7\]\[4\] _02979_ _02989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_88_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09280__I _04277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09312_ _04333_ _04334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07573_ _02945_ _02948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06524_ cpu.pwm_top\[7\] _01180_ _01408_ _02001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_36_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09243_ _00704_ _01016_ _04251_ _04267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06455_ _01357_ _01894_ _01932_ _01933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_90_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09174_ cpu.ROM_addr_buff\[10\] _04171_ _04205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06386_ cpu.timer_top\[6\] _01864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_8_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05406_ _00871_ _00896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05337_ cpu.PORTB_DDR\[4\] net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_08125_ _03378_ _03381_ _03382_ _00238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_16_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08056_ _03311_ _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_102_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05268_ _00779_ cpu.needs_interrupt _00780_ _00781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06144__I _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09907__A1 net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07007_ _02419_ _02479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05199_ cpu.base_address\[2\] _00714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput49 net49 io_oeb[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput38 net38 io_oeb[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08958_ _04031_ _04028_ _04032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05944__A2 _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07909_ _03199_ _03204_ _03205_ _03206_ _00199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_08889_ _03981_ _00404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07146__A1 _01774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08894__A1 _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09071__A1 _00971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_117_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10216_ _00111_ clknet_leaf_124_wb_clk_i cpu.regs\[12\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09374__A2 _01587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10147_ _00046_ clknet_leaf_31_wb_clk_i cpu.uart.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10078_ _01322_ _05018_ _05019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07137__A1 _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05699__A1 _01054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_99_Left_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06240_ _01688_ _01416_ _01589_ _01719_ _01720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_111_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08444__I cpu.Z vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05871__A1 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09062__A1 _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06171_ _00950_ _01339_ _01635_ _01330_ _01341_ _01652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_80_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05122_ _00621_ _00639_ _00640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09930_ _04027_ _04893_ _04894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05053_ _00573_ _00574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09861_ _04840_ _04841_ _00516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_5_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09792_ cpu.ROM_spi_dat_out\[1\] _02489_ _04784_ _04785_ _04786_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_08812_ _03916_ _03917_ _03918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08743_ _01395_ _01041_ _02709_ _03859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_05955_ _00844_ _00849_ _01320_ _01438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_108_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05886_ _01193_ _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08674_ _03800_ _03811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07679__A2 _03011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07523__I _02913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07625_ _01137_ _01156_ _02884_ _02976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_07556_ _02920_ _02932_ _02936_ _00116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06507_ net38 _01593_ _01983_ _01595_ _01984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_75_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07300__A1 _01202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09226_ _00657_ _01146_ _04251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07487_ cpu.regs\[14\]\[2\] _02889_ _02892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06438_ _01898_ _01900_ _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_90_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09157_ cpu.last_addr\[5\] _04192_ _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06369_ _01847_ _01829_ _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08108_ cpu.spi.counter\[1\] _03367_ _03369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09088_ _04139_ cpu.ROM_addr_buff\[3\] _04134_ _04140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08800__A1 cpu.timer_capture\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07603__A2 _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08039_ cpu.uart.receive_buff\[3\] _03307_ _03308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05614__A1 _01093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_112_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10001_ _04946_ _04944_ _04947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09913__I _04868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05473__S0 _00956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_48_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09788__C _04721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_80_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05888__I _01203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_78_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_87_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_38_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05740_ _01193_ _01224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05671_ _00930_ _01155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07410_ cpu.uart.receive_div_counter\[7\] _02821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08390_ _03570_ _03593_ _03594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_18_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07341_ _02761_ _02763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_58_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09283__A1 _01015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07272_ _02710_ _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06223_ _01224_ _01702_ _01703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09035__B2 _00967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09011_ _04059_ _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05844__A1 _00928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06154_ _01633_ _00949_ _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_103_Right_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05105_ _00587_ _00623_ _00624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06085_ _01555_ _01558_ _01564_ _01566_ _01567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_111_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09913_ _04868_ _04881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09338__A2 _04359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09844_ cpu.pwm_counter\[1\] _04826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09775_ _04770_ _04771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06987_ _00690_ _02458_ _02459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08726_ cpu.timer_top\[11\] _03842_ _03847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08849__A1 _03170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05938_ _01415_ _01418_ _01420_ _01421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_96_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08657_ _03796_ _03798_ _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09510__A2 _04500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05869_ _01312_ _01317_ _01324_ _01352_ _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_07608_ cpu.regs\[8\]\[0\] _02966_ _02967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05383__I0 cpu.regs\[8\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08588_ _03677_ cpu.toggle_ctr\[0\] _03752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09274__A1 _02768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07539_ _01858_ cpu.regs\[12\]\[5\] _02913_ _02925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_36_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10550_ _00444_ clknet_leaf_84_wb_clk_i cpu.ROM_addr_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10481_ _00376_ clknet_leaf_18_wb_clk_i cpu.timer_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_63_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05835__A1 _01170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09209_ _04228_ _04229_ _04230_ _04233_ _01976_ _04234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_0_32_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_121_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08687__C _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07355__A4 _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_4_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06315__A2 _01114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05411__I _00900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07539__S _02913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09981__C _04931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07338__I _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06910_ _02384_ _02045_ _02385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07890_ cpu.spi.divisor\[5\] _03188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06841_ _02306_ _02311_ _02316_ _02317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_65_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09560_ _03083_ _04550_ _04574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06772_ _02228_ _02227_ _02248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_78_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05723_ _01025_ _01028_ _01045_ _01207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_08511_ _03682_ _00325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09491_ _04456_ _04501_ _04508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08442_ cpu.orig_flags\[0\] _03615_ _03634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05654_ _01137_ _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_08373_ _03551_ _03580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05585_ _01068_ _01069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_81_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09256__A1 _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07324_ _02692_ _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10110__I0 _01934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06417__I _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07255_ _02696_ _00055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06490__A1 _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06206_ _01685_ _01686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_103_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07186_ _02635_ _02636_ _02637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06490__B2 _01452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06137_ _01118_ _01617_ _01618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06242__A1 _00951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06152__I _00840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06068_ _01364_ net91 _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09827_ _04807_ _04813_ _04809_ _04814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09758_ _04755_ _04740_ _04751_ _04757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_08709_ _03826_ _03834_ _03835_ _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_69_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09689_ _04169_ _04697_ _04698_ _04699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09495__A1 _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08807__I _03275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09247__A1 cpu.Z vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10602_ _00496_ clknet_leaf_76_wb_clk_i cpu.startup_cycle\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_12_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05371__I3 cpu.regs\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10533_ _00427_ clknet_leaf_40_wb_clk_i cpu.uart.divisor\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08470__A2 _03636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10464_ _00359_ clknet_leaf_14_wb_clk_i cpu.pwm_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_20_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10395_ _00290_ clknet_leaf_36_wb_clk_i cpu.uart.receive_div_counter\[10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07158__I _02612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05587__A3 _01008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07733__A1 _02014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06536__A2 _01977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06011__B cpu.PORTA_DDR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05406__I _00871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08717__I _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05370_ _00859_ _00860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_28_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_35_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_35_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_83_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07040_ _02497_ _02508_ _02509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08213__A2 _01395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08991_ _04057_ _01734_ _04058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08401__B _03600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07942_ _03220_ _03233_ _03234_ _00204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_76_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07873_ _03135_ _03149_ _03169_ _03171_ _03172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_09612_ _03672_ _04499_ _04624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07724__A1 cpu.regs\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06824_ _02299_ _02244_ _02300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09543_ _03060_ _00846_ _04558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06755_ _02229_ _02230_ _02231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05706_ _01186_ _01190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09474_ _04329_ _04474_ _04491_ _04366_ _04492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10087__A2 _05009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06686_ _02159_ _02160_ _02161_ _02162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__07531__I _01583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05637_ _01087_ _01120_ _01121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_08425_ _00675_ _03618_ _03619_ _03620_ _00301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09229__A1 _02334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08356_ _02855_ _03566_ _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05568_ _00677_ _01032_ _01052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07307_ _02639_ _02737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05051__I _00571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08287_ _03513_ _00270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05499_ _00982_ _00962_ _00984_ _00985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_07238_ _02679_ _02659_ _02674_ _02681_ _02682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_61_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07169_ _02612_ _02623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10180_ _00075_ clknet_leaf_101_wb_clk_i _00005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_70_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08537__I cpu.toggle_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05329__I0 cpu.regs\[8\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05670__B _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10516_ _00411_ clknet_leaf_53_wb_clk_i cpu.spi.divisor\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06454__A1 net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05257__A2 _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10447_ _00342_ clknet_leaf_5_wb_clk_i cpu.toggle_ctr\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10378_ _00273_ clknet_leaf_45_wb_clk_i cpu.uart.receive_buff\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06301__S1 _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05280__I2 _00790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06509__A2 _01070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06540_ _01361_ _02015_ _02016_ _00020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06471_ _01895_ _01896_ _01948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08210_ cpu.uart.has_byte _03450_ _03451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05422_ _00845_ _00908_ _00911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09190_ _01006_ _04216_ _04217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08141_ _03296_ _03396_ _00241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_71_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05353_ cpu.base_address\[1\] _00843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08072_ cpu.uart.div_counter\[9\] _03336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_71_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05284_ _00002_ _00794_ _00795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07023_ _00693_ _02039_ _02040_ _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08974_ _04044_ _00426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_89_Right_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07925_ _03217_ _03220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07856_ cpu.timer_top\[1\] _02667_ _02657_ cpu.timer_top\[0\] _03155_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_input18_I io_in[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07787_ cpu.spi.counter\[0\] cpu.spi.counter\[1\] _03094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06807_ _02280_ _02281_ _02283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09526_ _04358_ _04527_ _04541_ _04439_ _04542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06738_ _02196_ _02212_ _02213_ _02214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09457_ cpu.PC\[5\] _00701_ _04475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_98_Right_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08408_ _03607_ _03608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06684__A1 _00603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06669_ _02143_ _02144_ _02145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_50_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09388_ _04288_ _04409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_22_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08339_ _03544_ _03553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09622__A1 _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05239__A2 _00656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06436__A1 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10301_ _00196_ clknet_leaf_52_wb_clk_i cpu.spi.dout\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10232_ _00127_ clknet_leaf_116_wb_clk_i cpu.regs\[10\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10163_ _00062_ clknet_leaf_22_wb_clk_i cpu.timer_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05665__B _01148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07436__I cpu.uart.divisor\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09689__A1 _04169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10094_ _02885_ _02929_ _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_89_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06496__B _01325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06911__A2 _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06675__A1 _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09613__A1 _02062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_94_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05089__S1 _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07346__I cpu.PC\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07710_ _03006_ cpu.regs\[4\]\[6\] _03021_ _03031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05971_ _00814_ _01454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07155__A2 _00756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08690_ _02727_ _03802_ _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07641_ _02987_ _02980_ _02988_ _00149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07572_ _02946_ _02947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_50_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_50_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06523_ cpu.timer_top\[15\] _01404_ _01251_ _01999_ _02000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_09311_ _04309_ _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09242_ _03635_ _04227_ _04266_ _03920_ _00472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06454_ net32 _01580_ _01478_ _01931_ _01932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_106_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09173_ cpu.last_addr\[10\] _04204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_56_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06385_ _01862_ _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05405_ cpu.regs\[12\]\[1\] cpu.regs\[13\]\[1\] cpu.regs\[14\]\[1\] cpu.regs\[15\]\[1\]
+ _00888_ _00889_ _00895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_05336_ cpu.PORTA_DDR\[3\] net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
X_08124_ _03195_ _03212_ _03382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06418__A1 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08055_ cpu.uart.dout\[7\] _03300_ _03320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05267_ _00697_ net18 _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07006_ net54 _02477_ _02478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05198_ cpu.base_address\[3\] _00713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_12_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput39 net39 io_oeb[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07256__I cpu.timer\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08957_ _00903_ _04031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07908_ _03199_ _03204_ net70 _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08888_ cpu.timer_capture\[15\] _03965_ _03980_ _03968_ _03981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07839_ cpu.timer_top\[12\] _03136_ _03137_ cpu.timer_top\[11\] _03138_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_55_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_38_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09509_ _04524_ _04379_ _04525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_117_Right_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06409__A1 cpu.toggle_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05632__A2 _01100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10215_ _00110_ clknet_leaf_125_wb_clk_i cpu.regs\[12\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07166__I _02619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10146_ _00045_ clknet_leaf_41_wb_clk_i cpu.uart.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05396__A1 _00880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_77_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10077_ _01938_ _01962_ _05018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06196__I0 net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08885__A2 _02651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06896__A1 _02370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05414__I _00903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10179__D _00074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_96_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09984__C _04931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05871__A2 _01012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06170_ _01650_ _01651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05121_ cpu.regs\[8\]\[7\] cpu.regs\[9\]\[7\] cpu.regs\[10\]\[7\] cpu.regs\[11\]\[7\]
+ _00630_ _00631_ _00639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_110_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05052_ _00001_ _00573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09860_ _02503_ _00738_ _04841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_5_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09791_ _02488_ _04773_ _04785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_84_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08811_ _03909_ _03910_ _03143_ _03917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08742_ _03857_ _03858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05954_ _01435_ _01436_ _01437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08673_ _03810_ _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05139__A1 _00654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05885_ _00680_ _01066_ _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_07624_ _01358_ _02975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_88_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07555_ cpu.regs\[11\]\[2\] _02933_ _02936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06506_ net58 _01593_ _01983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09240__B _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07486_ _01482_ _02888_ _02891_ _00091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06437_ net96 _01914_ _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09225_ _04246_ _04249_ _04250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_60_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09156_ _04175_ _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06368_ _01426_ _01847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08107_ _03366_ _03220_ _03368_ _00234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09087_ _02803_ _04136_ _04138_ _04139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06299_ _01776_ _01777_ _00851_ _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05319_ _00802_ _00827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08038_ _02880_ _03307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_111_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10000_ _02441_ _04946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09989_ _04790_ _02425_ _02428_ cpu.ROM_spi_mode _04937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_99_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05473__S1 _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_67_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07055__A1 _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06802__A1 _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06014__B _01211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10129_ _00028_ clknet_leaf_85_wb_clk_i cpu.instr_buff\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_89_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07624__I _01358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05670_ _01153_ _01139_ _01149_ _01154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_18_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08455__I _03626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07340_ _02580_ _02760_ _02588_ _02762_ _00074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_72_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09283__A2 _04277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07271_ _01494_ _02709_ _02710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09010_ cpu.orig_IO_addr_buff\[0\] _04075_ _04076_ _01004_ _04077_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06222_ cpu.uart.divisor\[12\] _01700_ _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05844__A2 cpu.base_address\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07046__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06153_ _01436_ _01546_ _01634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08794__A1 cpu.timer_capture\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05104_ cpu.regs\[12\]\[6\] cpu.regs\[13\]\[6\] cpu.regs\[14\]\[6\] cpu.regs\[15\]\[6\]
+ _00615_ _00616_ _00623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_110_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06084_ _01144_ _01538_ _01565_ _01440_ _01566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09912_ _04868_ _04880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09843_ cpu.pwm_top\[7\] cpu.pwm_counter\[7\] _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09774_ _02476_ _04769_ _04770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06986_ _02026_ _02028_ _02458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07534__I _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08725_ _02627_ _03841_ _03846_ _03844_ _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05780__A1 _01262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05937_ _01419_ _01292_ _01293_ _01420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10105__A1 _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08656_ _02882_ _03797_ _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05054__I _00574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05868_ _01326_ _01327_ _01351_ _01352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08587_ _03750_ _03751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07607_ _02963_ _02966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07538_ _02924_ _00110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05799_ cpu.regs\[4\]\[7\] cpu.regs\[5\]\[7\] cpu.regs\[6\]\[7\] cpu.regs\[7\]\[7\]
+ _00855_ _01282_ _01283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_9_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07469_ cpu.uart.receive_counter\[3\] _02877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10480_ _00375_ clknet_leaf_18_wb_clk_i cpu.timer_top\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_63_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09208_ _01854_ _01930_ _04232_ _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_17_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09139_ _04171_ _04179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08785__A1 cpu.timer\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05771__A1 _01176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_107_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_107_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08275__I _00776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06079__A2 _00908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05826__A2 _01309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07028__A1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05848__B _01331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05429__I2 cpu.regs\[10\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06840_ _02314_ _02315_ _02316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06771_ _02243_ _00966_ net128 _02247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_05722_ _01201_ _01204_ _01205_ _01206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08510_ cpu.toggle_top\[0\] _03679_ _03681_ _03461_ _03682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09490_ _04504_ _04505_ _04506_ _04507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08441_ _03631_ _03632_ _03633_ _00304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05653_ _01133_ _01014_ _01136_ _01137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08372_ _03552_ _03579_ _00289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05584_ _01026_ _01029_ _01067_ _01068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_73_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09256__A2 _04277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05117__I1 _00634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07323_ _02749_ _00070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08913__I _03995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07254_ cpu.timer_capture\[5\] _02684_ _02695_ _02689_ _02696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_73_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06205_ _00983_ _00995_ _01684_ _01685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_6_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08134__B _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07185_ _02612_ _02636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06136_ cpu.timer_top\[3\] _01616_ _01617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06067_ _01541_ _01549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_111_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08519__A1 _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05049__I _00569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09826_ _02415_ _04812_ _04813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06969_ _02436_ _02437_ _02440_ _02441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XPHY_EDGE_ROW_100_Left_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09757_ _04740_ _04751_ _04755_ _04756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_5_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_5_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08708_ cpu.timer_div_counter\[5\] _03832_ _03835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09688_ _04174_ cpu.ROM_addr_buff\[0\] _04698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09495__A2 _04349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08639_ _03784_ _03783_ _03785_ _00350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08095__I _03358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10601_ _00495_ clknet_leaf_75_wb_clk_i cpu.startup_cycle\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10532_ _00426_ clknet_leaf_40_wb_clk_i cpu.uart.divisor\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05808__A2 _01115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10463_ _00358_ clknet_leaf_15_wb_clk_i cpu.pwm_top\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06481__A2 _01957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10394_ _00289_ clknet_leaf_37_wb_clk_i cpu.uart.receive_div_counter\[9\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_75_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07174__I _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08930__A1 _02746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10187__D _00082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08997__A1 _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_75_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_75_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_70_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08990_ _04056_ _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07941_ cpu.spi.data_out_buff\[2\] _03223_ _03228_ _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07872_ _03140_ _03170_ _03152_ _03154_ _03171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08921__A1 cpu.timer_div\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09611_ cpu.PC\[12\] _04623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06823_ _02151_ _02299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06754_ _02201_ _02203_ _02230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09542_ _04530_ _04531_ _04556_ _04557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_92_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05705_ _01076_ _01189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09473_ _04483_ _04488_ _04490_ _04491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06685_ _02156_ _02158_ _02161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05636_ _00674_ _00672_ _01119_ _01120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_08424_ _02602_ _03620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09229__A2 _02370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06160__A1 _01586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08355_ _02835_ _03556_ _03559_ _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_74_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05567_ _01050_ _01051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07306_ _02735_ _02733_ _02736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08286_ cpu.uart.data_buff\[9\] _03469_ _03484_ _03461_ _03513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05498_ _00983_ _00959_ _00984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_18_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07237_ _00978_ _02680_ _02681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07168_ cpu.uart.divisor\[1\] _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06119_ _01598_ _01599_ _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07099_ net19 _02361_ _02351_ _02564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09809_ _04771_ _04798_ _04799_ _00506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_70_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08553__I cpu.toggle_top\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10515_ _00410_ clknet_leaf_53_wb_clk_i cpu.spi.divisor\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07169__I _02612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10446_ _00341_ clknet_leaf_6_wb_clk_i cpu.toggle_ctr\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10377_ _00272_ clknet_leaf_46_wb_clk_i cpu.uart.receive_buff\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05280__I3 cpu.regs\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_122_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_122_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06390__A1 net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08728__I _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06470_ _01945_ _01946_ _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09987__C _04931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05421_ _00845_ _00909_ _00910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08140_ _03348_ _03394_ _03395_ _03384_ _03396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05352_ _00842_ net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08071_ cpu.uart.div_counter\[6\] _03335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_43_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05283_ cpu.regs\[12\]\[0\] cpu.regs\[13\]\[0\] cpu.regs\[14\]\[0\] cpu.regs\[15\]\[0\]
+ _00785_ _00786_ _00794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07022_ _00732_ _02492_ _02493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_71_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08973_ _02842_ _04040_ _04043_ _04035_ _04044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07924_ _02708_ _03212_ _03215_ _03219_ _00201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07855_ _03151_ cpu.timer\[15\] _03154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_108_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07786_ cpu.spi.data_in_buff\[0\] _03093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06806_ _02280_ _02281_ _02282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09525_ cpu.orig_PC\[8\] _04359_ _04541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06737_ _02210_ _02211_ _02213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_94_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06133__A1 cpu.timer_capture\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09456_ _04473_ _04474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06668_ _02115_ _02116_ _02144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08407_ _00670_ _03606_ _03607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05619_ _01096_ _01067_ _01103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05062__I _00581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09387_ _04383_ _04386_ _04405_ _04407_ _04408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06599_ _02073_ _02074_ _02075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_19_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08373__I _03551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08338_ _03551_ _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08269_ _02634_ _03486_ _03500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06436__A2 _01757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10300_ _00195_ clknet_leaf_51_wb_clk_i cpu.spi.dout\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10231_ _00126_ clknet_leaf_125_wb_clk_i cpu.regs\[10\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07717__I _03033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10162_ _00061_ clknet_leaf_18_wb_clk_i cpu.timer_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05947__A1 _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_67_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10093_ _05030_ _05031_ _05032_ _00557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09138__A1 _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05237__I _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06675__A2 _00875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05700__I _01183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09613__A2 _04499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06017__B _01216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_94_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10429_ _00324_ clknet_leaf_8_wb_clk_i cpu.toggle_clkdiv vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05970_ _01452_ _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07563__S _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07640_ cpu.regs\[7\]\[3\] _02979_ _02988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07571_ _02945_ _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06522_ _01980_ _01245_ _01997_ _01998_ _01247_ _01999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__09301__A1 _00724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09310_ _04331_ _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06115__A1 net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09241_ _04234_ _04235_ _04265_ _04227_ _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06453_ _01424_ _01930_ _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09172_ _04201_ _04202_ _04203_ _00465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_leaf_90_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_90_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06384_ _00983_ _01285_ _01861_ _01862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_05404_ _00880_ _00893_ _00894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05874__B1 _01356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05335_ cpu.PORTB_DDR\[3\] net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_08123_ cpu.spi.counter\[4\] _03380_ _03381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08054_ cpu.uart.receive_buff\[7\] _02880_ _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07005_ _02469_ _02474_ _02476_ _02477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_98_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05266_ cpu.IE _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_101_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05197_ cpu.base_address\[0\] _00712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05929__A1 cpu.toggle_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input30_I sram_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08956_ _04030_ _00422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_98_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07907_ cpu.spi.data_out_buff\[7\] _03101_ _03205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08887_ _03944_ _03979_ _03980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08368__I cpu.uart.receive_div_counter\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07838_ cpu.timer\[11\] _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06354__A1 _01446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07769_ net19 _03053_ _03077_ _03078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09508_ cpu.PC\[8\] _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_109_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09439_ cpu.PC\[4\] _00745_ _04458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_35_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05632__A3 _01115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09359__A1 _02052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06290__B1 _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10214_ _00109_ clknet_leaf_0_wb_clk_i cpu.regs\[12\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10145_ _00044_ clknet_leaf_42_wb_clk_i cpu.uart.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10076_ _01938_ _01291_ _01960_ _05017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_clkbuf_4_10_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06345__A1 _01326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06896__A2 _01290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05120_ _00587_ _00637_ _00638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05051_ _00571_ _00572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__05474__I3 cpu.regs\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08810_ _03143_ _03909_ _03910_ _03916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09790_ _02432_ _04745_ _04784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08741_ _03856_ _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05953_ _01316_ _01433_ _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_108_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08672_ cpu.pwm_top\[2\] _03801_ _03807_ _03809_ _03810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05884_ _01254_ _01367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09522__A1 _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05605__I _01088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07623_ _02927_ _02966_ _02974_ _00145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_105_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07554_ _02918_ _02932_ _02935_ _00115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06505_ net5 _01982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07485_ cpu.regs\[14\]\[1\] _02889_ _02891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06436_ net95 _01757_ _01914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09224_ _04247_ _04248_ _04249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09155_ cpu.ROM_addr_buff\[5\] _04179_ _04191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06367_ _01753_ _01755_ _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08106_ _03216_ _03367_ _03368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09086_ _04137_ _00832_ _04138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06298_ cpu.regs\[0\]\[6\] cpu.regs\[1\]\[6\] cpu.regs\[2\]\[6\] cpu.regs\[3\]\[6\]
+ _01775_ _00859_ _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_05318_ _00826_ net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_08037_ _03305_ _03306_ _02871_ _00227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_102_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05249_ _00762_ _00763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05075__A1 _00567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09988_ _04936_ _00548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05378__A2 _00866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08939_ _04016_ _00419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_98_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06327__A1 cpu.timer_capture\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06878__A2 _02062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07827__A1 cpu.timer_div\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06346__I _00612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07055__A2 _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10128_ _00027_ clknet_leaf_84_wb_clk_i cpu.base_address\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10059_ _02593_ _04240_ _04242_ _05000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_38_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06318__A1 cpu.uart.divisor\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_29_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_29_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05541__A2 net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07270_ _01082_ _02610_ _02709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06221_ _01692_ _01370_ _01698_ _01699_ _01700_ _01701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_100_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06152_ _00840_ _01633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05103_ _00617_ _00620_ _00621_ _00622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06083_ _01544_ _01565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09911_ _04879_ _00528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_79_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09842_ cpu.pwm_top\[4\] cpu.pwm_counter\[4\] _04824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_13_Left_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08546__A2 cpu.toggle_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09773_ _00688_ _02473_ _04768_ _04769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_06985_ _02426_ _02456_ _02457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08724_ cpu.timer_top\[10\] _03842_ _03846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05936_ _01340_ _01419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08655_ cpu.pwm_counter\[6\] _03795_ _03797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05867_ _01332_ _01342_ _01350_ _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_89_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08586_ _03749_ _03750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07606_ _02964_ _02965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07537_ _01772_ cpu.regs\[12\]\[4\] _02914_ _02924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05798_ _00858_ _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07550__I _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Left_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07468_ _02874_ _02876_ _00088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_64_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07399_ _02812_ _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06419_ _01895_ _01896_ _01897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09207_ _01579_ _01676_ _01767_ _04231_ _04232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_09138_ _03378_ _04173_ _04178_ _00456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_114_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08785__A2 cpu.timer\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09069_ _04125_ _00440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06796__A1 _02271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_31_Left_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06548__A1 _00682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output61_I net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05071__I1 _00590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05429__I3 cpu.regs\[11\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05864__B _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06770_ _02245_ _02244_ _02246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_05721_ _01199_ _01205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10099__A1 _01359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08440_ _03311_ _03633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05652_ _01135_ _01128_ _01107_ _00970_ _01136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_81_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08371_ _03576_ _03563_ _03553_ _03578_ _03579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_105_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05583_ _01040_ _01066_ _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_46_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07322_ cpu.toggle_top\[12\] _02745_ _02748_ _02737_ _02749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05117__I2 cpu.regs\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07253_ _02660_ _02694_ _02695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07184_ _02634_ _02635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06204_ _00982_ _00992_ _01684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_14_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09964__A1 _00904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06135_ _01238_ _01616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06066_ _01453_ _01548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09825_ _04810_ _04811_ _04812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05202__A1 cpu.base_address\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06968_ _02426_ _02439_ _02440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09756_ cpu.startup_cycle\[5\] _04755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09687_ cpu.last_addr\[1\] cpu.ROM_addr_buff\[1\] _04174_ _04697_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08707_ cpu.timer_div_counter\[5\] _03832_ _03834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05919_ _01232_ _01402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08638_ _03784_ _03783_ _03505_ _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06899_ _02373_ _01289_ _02374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08569_ _03725_ cpu.toggle_top\[5\] cpu.toggle_top\[4\] _03730_ _03733_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_10600_ _00494_ clknet_leaf_74_wb_clk_i cpu.startup_cycle\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07258__A2 _02698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10531_ _00425_ clknet_leaf_41_wb_clk_i cpu.uart.divisor\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_40_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10462_ _00357_ clknet_leaf_10_wb_clk_i cpu.pwm_top\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10393_ _00288_ clknet_leaf_37_wb_clk_i cpu.uart.receive_div_counter\[8\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09955__A1 _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07430__A2 cpu.uart.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05992__A2 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07194__A1 _02643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_48_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08694__A1 _02619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10005__A1 cpu.ROM_addr_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10005__B2 cpu.ROM_addr_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_7_0_wb_clk_i clknet_0_wb_clk_i clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08213__A4 _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07566__S _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07940_ cpu.spi.data_out_buff\[3\] _03230_ _03232_ _03233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_44_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_44_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07871_ cpu.timer\[8\] _03170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_92_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09610_ _04600_ _04622_ _00687_ _00484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06822_ _02288_ _02296_ _02298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09580__I _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06753_ _02227_ _02228_ _02229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09541_ _04532_ _04556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05704_ cpu.spi.divisor\[0\] _01188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09472_ _04388_ _04474_ _04489_ _04362_ _04490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_59_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08685__A1 _02755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06684_ _00603_ _00975_ _02160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05499__A1 _00982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05635_ _00644_ _00645_ _01119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07033__C _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08423_ cpu.orig_IO_addr_buff\[4\] _03615_ _03619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09229__A3 _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06160__A2 _00840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08354_ _03552_ _03565_ _00285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_86_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08924__I _02723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05566_ _01049_ _00645_ _01050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07305_ _00903_ _02735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08285_ _03499_ _03511_ _03512_ _00269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_73_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05497_ _00940_ _00983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_116_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07236_ _02658_ _02680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09937__A1 _04851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07167_ _02620_ _02621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06118_ net24 _01113_ _01088_ _01599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06380__S _01681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05423__A1 _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07098_ _02321_ _02562_ _02563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06049_ _01530_ _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07208__C _02610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09808_ cpu.ROM_spi_dat_out\[5\] _04772_ _02715_ _04799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_70_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09739_ _04733_ _04738_ _04742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06923__A1 _02150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_15_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07479__A2 _02885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_25_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10514_ _00409_ clknet_leaf_53_wb_clk_i cpu.spi.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_96_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10445_ _00340_ clknet_leaf_5_wb_clk_i cpu.toggle_ctr\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10376_ _00271_ clknet_leaf_44_wb_clk_i cpu.uart.receiving vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07185__I _02612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05965__A2 _01447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06390__A2 _01211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08744__I _03859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05420_ _00908_ _00909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05351_ net75 cpu.ROM_spi_mode _00842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_16_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08070_ _03333_ _01692_ _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_102_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05282_ _00593_ _00788_ _00792_ _00793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_07021_ _00668_ _00780_ _02492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05653__A1 _01133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08972_ _04041_ _04042_ _04043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05608__I _01091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07923_ _03201_ _03218_ _03219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07854_ _03135_ _03150_ _03152_ _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08919__I _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06805_ _02256_ _02255_ _02281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07785_ _03069_ _03091_ _03092_ _00189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_108_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05343__I cpu.PORTB_DDR\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09524_ _00752_ _04539_ _04540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06736_ _02210_ _02211_ _02212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09455_ _02050_ _04450_ _04473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06667_ _02136_ _02142_ _02143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08406_ _00723_ _03605_ _03606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05618_ _01095_ _01101_ _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05892__A1 cpu.PORTB_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09386_ _04406_ _04407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06598_ _00633_ _00965_ _02074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_22_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08337_ _02872_ _03551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_74_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05549_ _00646_ _01032_ _01033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_61_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08268_ _03477_ _03499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06174__I _01447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07219_ _02665_ _00050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08199_ _03427_ _03442_ _00253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10230_ _00125_ clknet_leaf_126_wb_clk_i cpu.regs\[10\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_72_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07397__A1 _02580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Left_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10161_ _00060_ clknet_leaf_20_wb_clk_i cpu.timer_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05947__A2 _00900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10092_ net69 _05031_ _05032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07149__A1 _02592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05518__I _00878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08897__A1 cpu.spi.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07321__A1 _02746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07872__A2 _03170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07401__C _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05883__A1 _01365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10428_ _00323_ clknet_leaf_57_wb_clk_i cpu.had_int vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10359_ _00254_ clknet_leaf_35_wb_clk_i cpu.uart.div_counter\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_94_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09129__A2 _04169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08888__A1 cpu.timer_capture\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06363__A2 _01840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_69_Left_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07570_ _01158_ _02405_ _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_06521_ cpu.timer_capture\[15\] _01402_ _01616_ _01998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_118_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09240_ _03635_ _04078_ _04235_ _04264_ _04265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_113_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07863__A2 _02697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06452_ net96 _01296_ _01929_ _01930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_103_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09171_ cpu.last_addr\[9\] _04192_ _04203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09065__A1 _02508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06383_ _00982_ _01281_ _01861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05403_ cpu.regs\[8\]\[1\] cpu.regs\[9\]\[1\] cpu.regs\[10\]\[1\] cpu.regs\[11\]\[1\]
+ _00882_ _00884_ _00893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_113_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08122_ _03379_ _03196_ _03375_ _03380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_71_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06418__A3 _01742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05334_ _00841_ net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_08053_ _03317_ _03318_ _03312_ _00231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_78_Left_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07004_ cpu.spi_clkdiv _02475_ _02476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05265_ _00695_ _00773_ _00774_ _00778_ _00008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05196_ _00705_ _00710_ _00711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_3_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08955_ cpu.uart.divisor\[8\] _04026_ _04029_ _04015_ _04030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05338__I cpu.PORTA_DDR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07906_ _03201_ _03203_ _03204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input23_I io_in[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08886_ cpu.timer\[15\] _03946_ _03978_ _03979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07837_ cpu.timer\[12\] _03136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__07551__A1 cpu.regs\[11\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07768_ _03053_ _03076_ _03077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09507_ _04521_ _04522_ _04523_ _00480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06719_ _02194_ _02195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07303__A1 _01004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07699_ _02975_ _03023_ _03025_ _00170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09438_ cpu.PC\[4\] _00745_ _04457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_35_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09369_ _04361_ _04390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06118__B _01088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output91_I net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09359__A2 _04379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06290__B2 _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10213_ _00108_ clknet_leaf_0_wb_clk_i cpu.regs\[12\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10144_ _00043_ clknet_leaf_41_wb_clk_i cpu.uart.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09943__I _04891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07463__I _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10075_ net97 _01863_ _01972_ _05016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_89_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xwrapped_qcpu_110 io_out[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_58_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08294__I _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05050_ _00570_ _00571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06542__I _01109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08740_ _03855_ _03175_ _03856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05952_ _01314_ _01435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08671_ _03808_ _03809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05883_ _01365_ _01165_ _01166_ _01366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__06336__A2 _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07622_ cpu.regs\[8\]\[7\] _02964_ _02974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_105_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05395__I0 cpu.regs\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07553_ cpu.regs\[11\]\[1\] _02933_ _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06504_ cpu.spi.dout\[7\] _01981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_64_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07484_ _01360_ _02888_ _02890_ _00090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07041__C _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06435_ _01326_ _01911_ _01912_ _01913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_32_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09223_ _01162_ _02293_ _04248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_86_Left_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09154_ _04187_ _04188_ _04190_ _00460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_75_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08105_ _03196_ _03213_ _03367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06366_ _01574_ _01827_ _01844_ _01845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09085_ _00697_ _04137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06297_ cpu.regs\[4\]\[6\] cpu.regs\[5\]\[6\] cpu.regs\[6\]\[6\] cpu.regs\[7\]\[6\]
+ _01775_ _00859_ _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_4_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05317_ _00566_ _00820_ _00825_ _00826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_116_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08036_ cpu.uart.dout\[2\] _03301_ _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05248_ _00761_ _00762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07548__I _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09210__A1 _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05179_ _00694_ _00695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_95_Left_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09987_ cpu.PORTA_DDR\[7\] _04926_ _04935_ _04931_ _04936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_99_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08938_ cpu.timer_div\[6\] _03996_ _04014_ _04015_ _04016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_4_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08869_ _03942_ _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_94_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09029__B2 _00978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06015__A1 cpu.PORTB_DDR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10127_ _00026_ clknet_leaf_85_wb_clk_i cpu.base_address\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08510__C _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07193__I _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10058_ _04246_ _04247_ _04245_ _04999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_18_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_69_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_69_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06537__I _02013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05441__I cpu.base_address\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06220_ _01195_ _01700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08491__A2 _03659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06151_ _01173_ _01631_ _01632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05102_ _00583_ _00621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06082_ _01447_ _01562_ _01563_ _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05301__I0 cpu.regs\[8\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09910_ net82 _04869_ _04878_ _04874_ _04879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_111_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09841_ net73 _04823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_111_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09772_ _04733_ _02456_ _04767_ _02487_ _04768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_06984_ _00663_ _00664_ _02456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_95_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08723_ _02624_ _03841_ _03845_ _03844_ _00374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05935_ _01417_ _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08654_ cpu.pwm_counter\[6\] _03795_ _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05866_ _01343_ _01348_ _01349_ _01318_ _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_95_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09259__A1 _00721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08585_ _03200_ _03748_ _03749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07605_ _02963_ _02964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05797_ _01279_ _01280_ _00852_ _01281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_88_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07536_ _02922_ _02915_ _02923_ _00109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05383__I3 cpu.regs\[11\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07467_ _02868_ _02875_ _02876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_9_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09206_ _01354_ _01475_ _04228_ _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_07398_ _00768_ _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06418_ net94 _00613_ _01742_ _01896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_17_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09137_ _04174_ _04177_ _04178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06349_ _01725_ _01736_ _01727_ _01828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_102_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07278__I _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09068_ _04121_ _04115_ _04122_ _04124_ _04125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_60_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06245__A1 _00596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08019_ cpu.spi.data_in_buff\[3\] _03291_ _03294_ cpu.spi.data_in_buff\[4\] _03295_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06796__A2 _00899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06548__A2 _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07745__A1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output54_I net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05071__I2 _00591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05261__I _00682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06293__S _01681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07188__I _02638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06236__A1 cpu.toggle_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06092__I _01321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_116_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_116_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06539__A2 _01681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05436__I _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05211__A2 _00721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05720_ _01203_ _01204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09071__C _04124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05651_ _01134_ _01135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08370_ _03576_ _03577_ _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_105_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05514__A3 _00999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05582_ _01048_ _01055_ _01066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__05171__I _00686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07321_ _02746_ _02747_ _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07252_ _02691_ _02686_ _02693_ _02694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07183_ _00987_ _02634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06203_ _01267_ _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09413__A1 _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06134_ _01591_ _01233_ _01613_ _01614_ _01239_ _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_5_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06065_ _01436_ _01546_ _01547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_47_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05450__A2 _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09824_ cpu.ROM_spi_cycle\[2\] _04811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05346__I cpu.PORTA_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05202__A2 _00712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06967_ _02431_ _02438_ _02439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09755_ _04754_ _00497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09686_ cpu.last_addr\[3\] cpu.ROM_addr_buff\[3\] _04676_ _04696_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08706_ _03826_ _03832_ _03833_ _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_69_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05918_ cpu.timer_capture\[9\] _01401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06898_ _00619_ _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08637_ cpu.pwm_counter\[1\] _03784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05849_ _00799_ _01309_ _01333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_64_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08568_ _03730_ cpu.toggle_top\[4\] cpu.toggle_top\[3\] _03731_ _03732_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08499_ cpu.PC\[13\] _03674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07519_ _01359_ _02910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10530_ _00424_ clknet_leaf_41_wb_clk_i cpu.uart.divisor\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_86_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10461_ _00356_ clknet_leaf_16_wb_clk_i cpu.pwm_counter\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06218__A1 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10392_ _00287_ clknet_leaf_38_wb_clk_i cpu.uart.receive_div_counter\[7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_20_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07718__A1 cpu.regs\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09891__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08446__A2 _03636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10659_ _00553_ clknet_leaf_71_wb_clk_i net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05432__A2 _00920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07870_ _03138_ _03146_ _03141_ _03168_ _03169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_06821_ _02288_ _02296_ _02297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_84_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_84_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09540_ _04554_ _04555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_50_Left_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06752_ _02217_ _02218_ _02228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05703_ _01186_ _01187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09471_ cpu.orig_PC\[6\] _04359_ _04489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_13_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_13_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09882__A1 _04041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08422_ _03609_ _03618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06683_ _02156_ _02158_ _02159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_86_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05634_ _01083_ _01090_ _01118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_clkbuf_leaf_120_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08353_ _02835_ _03563_ _03553_ _03564_ _03565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05565_ _01048_ _01049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09229__A4 _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08284_ cpu.uart.data_buff\[9\] _03471_ _03505_ _03512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07304_ _01256_ _02732_ _02734_ _02724_ _00066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_6_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06448__A1 _01447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07235_ cpu.timer\[3\] _02679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_6_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05496_ _00867_ _00982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_33_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07166_ _02619_ _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_3_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06117_ net62 _01069_ _01596_ _01597_ _01216_ _01598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_100_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07948__A1 _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07097_ _02305_ _02319_ _02320_ _02562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_2_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06460__I _00642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06048_ _00826_ _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05076__I _00596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09807_ cpu.ROM_spi_dat_out\[4\] _04790_ _04792_ _04798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07999_ _03190_ _03253_ _03273_ _03281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09738_ _04738_ _04741_ _00778_ _00493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05726__A3 _01101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08125__A1 _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05804__I _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09669_ _04197_ _04678_ _04679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__05329__I3 cpu.regs\[11\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09625__A1 _00762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06439__B2 _01336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10513_ _00408_ clknet_leaf_53_wb_clk_i cpu.spi.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10444_ _00339_ clknet_leaf_7_wb_clk_i cpu.toggle_ctr\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07667__S _02994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10375_ _00270_ clknet_leaf_47_wb_clk_i cpu.uart.data_buff\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07939__A1 _03231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05725__I0 cpu.PORTA_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05350_ cpu.PORTB_DDR\[2\] net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_71_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_112_Right_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_99_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05281_ _00579_ _00791_ _00792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07020_ _02478_ _02491_ _00739_ _00025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_102_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08971_ _04025_ _04042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07922_ _03217_ _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07853_ _03151_ cpu.timer\[15\] cpu.timer\[14\] _03133_ _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06804_ _02277_ _02279_ _02280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08107__A1 _03366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07784_ _00832_ _03069_ _03092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_108_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09523_ _01002_ _04430_ _04538_ _04434_ _04539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06735_ _02177_ _02178_ _02211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09454_ _04448_ _04472_ _04417_ _00478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06666_ _02140_ _02141_ _02142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08405_ cpu.instr_cycle\[3\] cpu.instr_cycle\[1\] _03605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05617_ _01050_ _01041_ _01101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09385_ _04365_ _04406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08336_ _03514_ _03549_ _03550_ _00282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09607__A1 _00832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06597_ _00618_ _00998_ _02073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_22_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05548_ _00674_ _01031_ _01032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_50_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08267_ _03481_ _03496_ _03498_ _00265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_61_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05479_ _00965_ _00966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_104_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08198_ _03439_ _03405_ _03441_ _03408_ _03442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07218_ cpu.timer_capture\[0\] _02656_ _02663_ _02664_ _02665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08670__I _02638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07149_ _02592_ _02600_ _02605_ _02603_ _00040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_42_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10160_ _00059_ clknet_leaf_19_wb_clk_i cpu.timer_top\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_30_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10091_ _03253_ _03242_ _02517_ _05031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_76_Right_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_58_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_106_Left_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08845__I _01241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_85_Right_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07085__A1 _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10427_ _00322_ clknet_leaf_86_wb_clk_i cpu.orig_PC\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09609__C _04081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08513__C _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_115_Left_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05709__I _00681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08585__A1 _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10358_ _00253_ clknet_leaf_34_wb_clk_i cpu.uart.div_counter\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10289_ _00184_ clknet_leaf_116_wb_clk_i cpu.regs\[3\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_94_Right_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06899__A1 _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06520_ cpu.timer_capture\[7\] _01182_ _01994_ _01996_ _01243_ _01997_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_06451_ _01908_ _01913_ _01928_ _01929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_118_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05402_ _00886_ _00891_ _00892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09170_ cpu.ROM_addr_buff\[9\] _04194_ _04202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06382_ _01146_ _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_8_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08121_ _03098_ _03379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05333_ _00840_ _00841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08052_ cpu.uart.dout\[6\] _03309_ _03318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05264_ _00777_ _00778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_43_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07003_ _02417_ _02418_ _02475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_98_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05195_ _00706_ _00709_ _00710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_3_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08954_ _04027_ _04028_ _04029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07905_ _03202_ _03203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08885_ _03947_ _02651_ _03978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07836_ _03133_ cpu.timer\[14\] cpu.timer\[13\] _03134_ _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_input16_I io_in[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07767_ _02534_ _03072_ _03075_ _03076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_69_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09506_ _00686_ _04523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06718_ _00590_ _00975_ _02194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08500__A1 _03674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07698_ cpu.regs\[4\]\[0\] _03024_ _03025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09437_ _04455_ _04456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06649_ _02121_ _02122_ _02125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_35_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09368_ cpu.orig_PC\[3\] _04388_ _04389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08319_ _03536_ _00279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_62_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09299_ _00759_ _04318_ _04321_ _04284_ _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_50_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10212_ _00107_ clknet_leaf_4_wb_clk_i cpu.regs\[12\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10143_ _00042_ clknet_leaf_41_wb_clk_i cpu.uart.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10074_ _04121_ _01313_ _05014_ _05015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xwrapped_qcpu_100 io_oeb[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_qcpu_111 io_oeb[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_57_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07058__A1 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06281__A2 _00977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input8_I io_in[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07654__I _02994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07781__A2 _03085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05951_ _01316_ _01433_ _01434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08670_ _02638_ _03808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05882_ _01364_ _01365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07621_ _02973_ _00144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05395__I1 cpu.regs\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07552_ _02910_ _02932_ _02934_ _00114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06503_ cpu.timer_top\[7\] _01980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07297__A1 _02727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07483_ cpu.regs\[14\]\[0\] _02889_ _02890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06434_ _01822_ _01910_ _01909_ _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_17_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09222_ _01365_ _02270_ _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09153_ _04189_ _04177_ _04190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_60_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06365_ _01441_ _01829_ _01831_ _01833_ _01843_ _01844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_17_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08104_ _00777_ _03366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08434__B _03600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08797__A1 _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05316_ _00566_ _00822_ _00824_ _00825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09084_ _00697_ _04136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06296_ net124 _01775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_32_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08035_ cpu.uart.receive_buff\[2\] _02881_ _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05247_ _00706_ _00760_ _00709_ _00761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_3_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05349__I cpu.PORTB_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05178_ _00689_ _00693_ _00694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_3_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09986_ _02726_ _04927_ _04935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08937_ _04002_ _04015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08868_ _03964_ _00400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_99_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07819_ cpu.timer_div\[3\] cpu.timer_div_counter\[3\] _03118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08721__A1 _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08799_ _03170_ _03894_ _03904_ _03906_ _03898_ _03907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__05812__I _00654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06263__A2 _01742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05310__I1 _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06015__A2 _01211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10126_ _00025_ clknet_leaf_72_wb_clk_i net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05774__A1 _01256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10057_ _04245_ _04250_ _04998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_18_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08238__C _03474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05541__A4 _00669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07279__A1 _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_38_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_38_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_102_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06150_ cpu.TIE _01171_ _01630_ _01631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_80_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05101_ cpu.regs\[0\]\[6\] _00619_ cpu.regs\[2\]\[6\] cpu.regs\[3\]\[6\] _00615_
+ _00616_ _00620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06081_ _01444_ _01561_ _01560_ _01563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05301__I1 cpu.regs\[9\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_37_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09864__I _04843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09840_ _03207_ _04822_ _00514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_111_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09771_ _00663_ _04766_ _04767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06983_ _02449_ _02454_ _02455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_111_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08722_ cpu.timer_top\[9\] _03842_ _03845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05934_ _00937_ _01416_ _01277_ _01417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_37_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08653_ _03789_ _03794_ _03795_ _00354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05865_ _00849_ _01320_ _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08584_ _03677_ _03747_ _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_05796_ cpu.regs\[8\]\[7\] cpu.regs\[9\]\[7\] cpu.regs\[10\]\[7\] cpu.regs\[11\]\[7\]
+ _00864_ _00865_ _01280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07604_ _01158_ _02912_ _02963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_88_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07535_ cpu.regs\[12\]\[3\] _02914_ _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07466_ cpu.uart.receive_counter\[2\] _02866_ _02875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07987__C _02753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09205_ _01731_ _01819_ _01916_ _01945_ _04230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
X_06417_ _00628_ _01895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05376__S0 _00864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08219__B1 _03453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_76_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07397_ _02580_ _02811_ _02601_ _02763_ _00082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__07559__I _01771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09136_ _04176_ _04177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06348_ _01826_ _01757_ _01827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09067_ _04123_ _04124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_71_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06245__A2 _00985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06279_ net94 _01758_ _01759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08018_ _03286_ _03294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05079__I _00575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07495__S _02886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09707__C _03920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07294__I _02651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09969_ cpu.PORTA_DDR\[2\] _04915_ _04922_ _04920_ _04923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05807__I _01290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07745__A2 _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output47_I net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05071__I3 cpu.regs\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05119__S0 _00630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08933__A1 _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10109_ _05042_ _00563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05650_ cpu.br_rel_dest\[3\] _01134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05581_ _01035_ _01064_ _01065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_clkbuf_leaf_110_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07320_ _02731_ _02747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09661__A2 _04020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07251_ _02692_ _02680_ _02693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07182_ _02633_ _00045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06202_ _01160_ _01680_ _01682_ _00016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06227__A2 _01183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06133_ cpu.timer_capture\[3\] _01235_ _01232_ _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_41_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09808__B _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06064_ _01301_ _01538_ _01545_ _01546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09823_ cpu.ROM_spi_cycle\[3\] _04810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05202__A3 _00716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06966_ cpu.startup_cycle\[2\] _02438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_09754_ _02436_ _04750_ _04753_ _04721_ _04754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08705_ cpu.timer_div_counter\[3\] _03829_ cpu.timer_div_counter\[4\] _03833_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05917_ _01394_ _01398_ _01399_ _01243_ _01400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_09685_ _04189_ cpu.ROM_addr_buff\[4\] _04677_ _04695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_55_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06897_ _02369_ _02371_ _02372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08636_ _03781_ _03783_ _00349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05848_ net90 _00878_ _01331_ _01332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_64_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05362__I _00851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05779_ _01016_ _01263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08567_ cpu.toggle_ctr\[3\] _03731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08498_ _03672_ _03651_ _03673_ _03653_ _00321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_9_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07518_ _02015_ _02901_ _02909_ _00105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07449_ cpu.uart.divisor\[11\] cpu.uart.receive_div_counter\[11\] _02860_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_107_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_40_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07289__I _00776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10460_ _00355_ clknet_leaf_16_wb_clk_i cpu.pwm_counter\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06218__A2 _01114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09119_ _04162_ _00453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09404__A2 _01586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10391_ _00286_ clknet_leaf_35_wb_clk_i cpu.uart.receive_div_counter\[6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_20_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05977__A1 _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09168__A1 _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06368__I _01426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05272__I net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10658_ _00552_ clknet_leaf_71_wb_clk_i net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10589_ _00483_ clknet_leaf_95_wb_clk_i cpu.PC\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08906__A1 _02643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06820_ _02289_ _02295_ _02296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06751_ _02197_ _02198_ _02227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_92_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05702_ _01075_ _01185_ _01186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09470_ _04347_ _04487_ _04488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06682_ _00633_ _02157_ _02158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08421_ _01058_ _03610_ _03617_ _03613_ _00300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_59_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06145__A1 _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05633_ _01081_ _01023_ _01114_ _01116_ _01117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_08352_ _02835_ _03560_ _03564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xclkbuf_leaf_53_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_53_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05564_ cpu.IO_addr_buff\[1\] _01048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__09634__A2 _04296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08283_ cpu.uart.data_buff\[8\] _03465_ _03510_ _03511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05495_ _00981_ net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07303_ _01004_ _02733_ _02734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07234_ _02678_ _00052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07165_ _02516_ _02619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_74_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06116_ net42 _01374_ _01069_ _01597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__08070__A1 _03333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07096_ _02559_ _02560_ _02561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05959__A1 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06047_ _01528_ _01529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_10_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09806_ _04797_ _00505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06389__S _01207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07998_ _03103_ _03242_ _03279_ _03253_ _03280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__09570__A1 _04456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09737_ _04734_ _04740_ _04741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06949_ cpu.startup_cycle\[6\] _02421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__05431__I0 cpu.regs\[12\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09668_ cpu.last_addr\[6\] cpu.last_addr\[5\] cpu.last_addr\[4\] _04677_ _04678_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_09599_ _04610_ _04611_ _04612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08619_ _03753_ _03772_ _00343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_25_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06439__A2 _01784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10512_ _00407_ clknet_leaf_20_wb_clk_i cpu.spi.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10443_ _00338_ clknet_leaf_6_wb_clk_i cpu.toggle_ctr\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10374_ _00269_ clknet_leaf_47_wb_clk_i cpu.uart.data_buff\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06298__S1 _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05178__A2 _00693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06299__S _00851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06375__A1 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07482__I _02886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09313__A1 cpu.PC\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07875__A1 _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06678__A2 _00933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09202__I _04226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05280_ cpu.regs\[0\]\[0\] _00789_ _00790_ cpu.regs\[3\]\[0\] _00785_ _00786_ _00791_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_113_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10016__C _03366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08970_ _00987_ _04041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__05177__I _00692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05810__B1 _01291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_100_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_100_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09805__C _04788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07921_ _03216_ _03195_ _03217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07852_ cpu.timer_top\[15\] _03151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput1 io_in[0] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06803_ _02273_ _02278_ _02279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09522_ _04057_ _04526_ _04537_ _04432_ _04538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07783_ _01678_ _03090_ _02023_ _03091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06118__A1 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06734_ _02205_ _02206_ _02209_ _02210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_66_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09453_ _04381_ _04468_ _04471_ _04472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06665_ _02134_ _02135_ _02141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08404_ _03514_ _00698_ _03604_ _00296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08437__B _03600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09384_ _04391_ _04404_ _04405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05616_ _01010_ _00747_ _01099_ _01100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_08335_ cpu.uart.receive_div_counter\[1\] _03537_ _02824_ _03550_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06596_ _02070_ _02071_ _02068_ _02072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_22_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05547_ _00672_ _01031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_50_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08266_ cpu.uart.data_buff\[5\] _03497_ _03489_ _03498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08951__I _04025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05478_ _00964_ _00965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08197_ _03439_ _03440_ _03441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07217_ _02639_ _02664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05644__A3 _01093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07148_ _01860_ _02598_ _02605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_72_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07079_ _02545_ _00030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09715__C _04721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10090_ _03216_ _03371_ _05030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_58_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06380__I1 cpu.regs\[9\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10124__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08282__A1 _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10426_ _00321_ clknet_leaf_85_wb_clk_i cpu.orig_PC\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08585__A2 _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10357_ _00252_ clknet_leaf_35_wb_clk_i cpu.uart.div_counter\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_94_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10288_ _00183_ clknet_leaf_100_wb_clk_i cpu.regs\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_87_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06450_ _01574_ _01915_ _01923_ _01927_ _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_118_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06520__A1 cpu.timer_capture\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05401_ _00887_ _00890_ _00867_ _00891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_103_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06381_ _01859_ _00018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08273__A1 _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08120_ _00777_ _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05332_ _00593_ _00834_ _00839_ _00840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_22_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08051_ cpu.uart.receive_buff\[6\] _03307_ _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05263_ _00776_ _00777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07002_ _02472_ _02473_ _02474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08025__A1 _03296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06291__I _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09073__I0 _00790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05194_ _00708_ cpu.instr_buff\[14\] _00709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09816__B _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09773__A1 _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08576__A2 _01256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06587__A1 _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08953_ _04025_ _04028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07904_ _03100_ _03195_ _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08884_ _03977_ _00403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06339__A1 _00612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07000__A2 _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07835_ cpu.timer_top\[13\] _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_55_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07766_ _02523_ _03074_ _03075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_69_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07839__B2 cpu.timer_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09505_ _02570_ _04297_ _04522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06717_ _02190_ _02191_ _02192_ _02193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08500__A2 _03611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09436_ _04308_ _04455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07697_ _03021_ _03024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_109_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06648_ _00804_ _01954_ _02124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05370__I _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09367_ _04239_ _04388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06579_ _02052_ _02053_ _02054_ _02055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08318_ net15 _03521_ _03526_ cpu.uart.receive_buff\[7\] _03474_ _03536_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_09298_ _04319_ _04300_ _04320_ _04321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08249_ _03477_ _03484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10211_ _00106_ clknet_leaf_3_wb_clk_i cpu.regs\[12\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output77_I net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10142_ _00041_ clknet_leaf_108_wb_clk_i cpu.br_rel_dest\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10073_ _01941_ _05010_ _01951_ _01940_ _05013_ _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_89_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_qcpu_101 io_oeb[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_97_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_qcpu_112 io_oeb[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_43_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10409_ _00304_ clknet_leaf_56_wb_clk_i cpu.orig_IO_addr_buff\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05950_ _01426_ _01429_ _01432_ _01433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_108_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05881_ _01363_ _01364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07620_ _02942_ cpu.regs\[8\]\[6\] _02963_ _02973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_105_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07551_ cpu.regs\[11\]\[0\] _02933_ _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06502_ _01021_ _01272_ _01979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07482_ _02886_ _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_66_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06433_ _01822_ _01909_ _01910_ _01911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_32_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09221_ _01163_ _02772_ _02778_ _01365_ _04246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_118_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09152_ cpu.last_addr\[4\] _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_60_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06364_ _01438_ _01835_ _01836_ _01453_ _01842_ _01843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_17_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08103_ _03322_ _03360_ _03361_ _00239_ _00233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05315_ _00580_ _00823_ _00824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09083_ _04135_ _00444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06295_ _00743_ _01774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08034_ _03303_ _03304_ _02871_ _00226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05246_ _00705_ _00760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05177_ _00692_ _00693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_110_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08450__B _03633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09985_ _04934_ _00547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05232__A1 _00701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08936_ _02755_ _04009_ _04014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05365__I _00854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08867_ cpu.timer_capture\[11\] _03943_ _03963_ _03951_ _03964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07818_ cpu.timer_div\[4\] cpu.timer_div_counter\[4\] _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08798_ _03170_ _03905_ _03906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_8_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_8_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_67_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07749_ _03059_ _00186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_80_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09419_ _04361_ _04439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_94_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10044__A1 _00693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06099__I0 net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05310__I2 _00818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05476__S _00871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09175__C _04006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10125_ _00024_ clknet_leaf_103_wb_clk_i cpu.regs\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_89_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10056_ _00653_ _01334_ _04226_ _04997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_98_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_100_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08476__A1 _02559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05100_ _00618_ _00619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06080_ _01444_ _01560_ _01561_ _01562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_110_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_78_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_78_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05301__I2 cpu.regs\[10\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09880__I _04843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_107_Right_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09770_ _00664_ _04763_ _04765_ _02434_ _04766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06982_ _02025_ _02442_ _02444_ _02038_ _02454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_111_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08721_ _02708_ _03841_ _03843_ _03844_ _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05933_ _01273_ _01416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09813__C _04788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08652_ cpu.pwm_counter\[5\] _03792_ _03791_ _03795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_07603_ _02015_ _02960_ _00137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05864_ _00971_ _01346_ _01347_ _01348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_37_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08583_ _03746_ _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_05795_ cpu.regs\[12\]\[7\] cpu.regs\[13\]\[7\] cpu.regs\[14\]\[7\] cpu.regs\[15\]\[7\]
+ _00864_ _00865_ _01279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_66_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07534_ _01679_ _02922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07465_ _02873_ _02874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09204_ _01465_ _01444_ _01560_ _01650_ _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__05376__S1 _00865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06416_ _01860_ _01164_ _01892_ _01893_ _01894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_60_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07396_ _02599_ _02811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_8_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09135_ _04175_ _04176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06347_ _01825_ _01826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09066_ _02501_ _04123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_102_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06278_ _01672_ _01745_ _01758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08017_ _03289_ _03293_ _00220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05229_ _00704_ _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05205__A1 cpu.uart.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09968_ _04851_ _04916_ _04922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05095__I _00567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08919_ _02501_ _04002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09899_ _04027_ _04870_ _04871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08458__A1 _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07130__A1 _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10017__A1 _04147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07681__A2 _03011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09958__A1 _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05119__S1 _00631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10108_ _02365_ cpu.regs\[15\]\[5\] _05033_ _05042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09633__C _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10039_ _02474_ _04981_ _04982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_125_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_125_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_105_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05580_ _01037_ _01063_ _01064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_86_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07121__A1 _00692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07250_ _01688_ _02692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_61_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07181_ _02630_ _02613_ _02632_ _02518_ _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_6_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06201_ cpu.regs\[9\]\[3\] _01681_ _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05683__A1 _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06132_ cpu.timer_div\[3\] _01396_ _01609_ _01611_ _01612_ _01613_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_5_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_113_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07395__I _02810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06063_ _01301_ _01544_ _01545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07328__C _02753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09822_ _02416_ _04809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09753_ _02422_ _04740_ _04751_ _04752_ _04753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__06935__A1 _02150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06965_ _02430_ _02437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08704_ cpu.timer_div_counter\[3\] cpu.timer_div_counter\[4\] _03829_ _03832_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_09684_ cpu.last_addr\[6\] _04693_ _04694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05916_ cpu.timer_capture\[1\] _01235_ _01399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06896_ _02370_ _01290_ _02342_ _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08635_ _03782_ _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05847_ _01330_ _01331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_89_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08566_ cpu.toggle_ctr\[4\] _03730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07517_ cpu.regs\[13\]\[7\] _02899_ _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05778_ _01168_ _01262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_92_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08497_ cpu.orig_PC\[12\] _03609_ _03673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07448_ _02845_ _02859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_91_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07379_ _02253_ _02796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09118_ _04161_ cpu.ROM_addr_buff\[11\] _04159_ _04162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07415__A2 cpu.uart.receive_div_counter\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10390_ _00285_ clknet_leaf_35_wb_clk_i cpu.uart.receive_div_counter\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09049_ _04102_ _04109_ _00436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05285__S0 _00785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08679__A1 _02746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_86_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06154__A2 _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07351__A1 _02768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10657_ _00551_ clknet_leaf_70_wb_clk_i net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05665__A1 _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09628__C _04313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10588_ _00482_ clknet_leaf_98_wb_clk_i cpu.PC\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09644__B _04455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05276__S0 _00785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05463__I _00950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06750_ _02220_ _02225_ _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05701_ _01119_ _01185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06681_ _00906_ _02157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08420_ cpu.orig_IO_addr_buff\[3\] _03615_ _03617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05632_ _01064_ _01100_ _01115_ _01116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__07342__A1 _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08351_ _03517_ _03563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_86_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05563_ _01039_ _01042_ _01046_ _01047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08282_ _02726_ _03468_ _03510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08842__A1 _01055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05494_ _00968_ _00980_ _00981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_46_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07302_ _02731_ _02733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07233_ cpu.timer_capture\[2\] _02656_ _02677_ _02664_ _02678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xclkbuf_leaf_93_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_93_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_46_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07164_ _02618_ _00042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_22_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_22_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_42_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06115_ net53 _01593_ _01594_ _01595_ _01596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_07095_ _02057_ _02560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05959__A2 _01340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05638__I _01121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06046_ _01341_ _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09805_ cpu.ROM_spi_dat_out\[4\] _04778_ _04796_ _04788_ _04797_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07997_ _03278_ _03279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06948_ _02419_ _02420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09736_ _04739_ _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09667_ _04184_ _04676_ _04677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_06879_ net1 _02041_ _02355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08618_ _03741_ _03771_ _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09598_ _04578_ _04581_ _04611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08549_ _03707_ _03710_ _03712_ _03713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_25_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10511_ _00406_ clknet_leaf_21_wb_clk_i cpu.spi.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10442_ _00337_ clknet_leaf_7_wb_clk_i cpu.toggle_ctr\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10373_ _00268_ clknet_leaf_48_wb_clk_i cpu.uart.data_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09010__B2 _01004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06379__I _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08824__A1 cpu.timer_capture\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_99_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07938__I _00951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07920_ cpu.spi.counter\[0\] _03216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07851_ _03138_ _03147_ _03149_ _03150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput2 io_in[10] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06802_ _00805_ _00974_ _02278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07782_ net20 _03053_ _03089_ _03090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09521_ _04524_ _04351_ _04537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06733_ _02207_ _02208_ _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_108_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06118__A2 _01113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07315__A1 _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07866__A2 _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09452_ _04443_ _04452_ _04470_ _04413_ _04414_ _04471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06664_ _02137_ _02139_ _02140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08403_ cpu.had_int _03603_ cpu.needs_interrupt _03604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09068__A1 _04121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09383_ _04398_ _04403_ _00751_ _04404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05615_ cpu.br_rel_dest\[7\] _01019_ _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_06595_ _00589_ _01955_ _02071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08334_ _02824_ _03542_ _03544_ _03548_ _03549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_86_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05546_ _01029_ _01030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_52_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08815__A1 _01486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08265_ _03477_ _03497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05477_ _00963_ _00964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_116_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08196_ _03435_ _03440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07216_ _02657_ _02659_ _02660_ _02662_ _02663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07147_ _02590_ _02600_ _02604_ _02603_ _00039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08579__B1 cpu.toggle_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07078_ _02334_ _02533_ _02544_ _02545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06029_ _01510_ _01368_ _01397_ _01511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_100_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06199__I _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09719_ _02462_ _04724_ _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07306__A1 _02735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_6_0_wb_clk_i clknet_0_wb_clk_i clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_2_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09059__A1 _01002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05868__A1 _01326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10425_ _00320_ clknet_leaf_86_wb_clk_i cpu.orig_PC\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_17_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09082__I1 cpu.ROM_addr_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05278__I cpu.regs\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10356_ _00251_ clknet_leaf_34_wb_clk_i cpu.uart.div_counter\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_94_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10287_ _00182_ clknet_leaf_114_wb_clk_i cpu.regs\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_20_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_29_Left_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06348__A2 _01757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09298__A1 _04319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_1_Left_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_56_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05400_ cpu.regs\[4\]\[1\] cpu.regs\[5\]\[1\] cpu.regs\[6\]\[1\] cpu.regs\[7\]\[1\]
+ _00888_ _00889_ _00890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XPHY_EDGE_ROW_38_Left_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_113_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06380_ _01858_ cpu.regs\[9\]\[5\] _01681_ _01859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05331_ _00836_ _00838_ _00593_ _00839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__07076__A3 _02541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08050_ _03315_ _03316_ _03312_ _00230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05262_ _00775_ _00776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07001_ cpu.spi_clkdiv _02418_ _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_52_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09073__I1 _02768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05193_ _00707_ _00708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__09222__A1 _01365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_47_Left_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06587__A2 _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07784__A1 _00832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08952_ _02614_ _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07903_ _03200_ _03201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09525__A2 _04359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08883_ cpu.timer_capture\[14\] _03965_ _03976_ _03968_ _03977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07834_ cpu.timer_top\[14\] _03133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06339__A2 _01685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_95_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09289__A1 _04309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07765_ _03073_ _02329_ _03074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_69_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09504_ _04328_ _04517_ _04520_ _04521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06716_ _00900_ _02190_ _02192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07696_ _03022_ _03023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_56_Left_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09435_ _04387_ _04452_ _04453_ _04390_ _04454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06647_ _02121_ _02122_ _02123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_93_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08962__I _04002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09366_ _04061_ _04387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06578_ cpu.PC\[1\] _02054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_117_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08317_ _03532_ _03535_ _00278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09297_ _02778_ _04319_ _04320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05529_ _00654_ _01011_ _01012_ _01013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_117_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08248_ cpu.uart.data_buff\[1\] _03469_ _03482_ _03483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06275__A1 _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08179_ _03336_ _03424_ _03426_ _03097_ _00249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_EDGE_ROW_65_Left_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09213__A1 _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10210_ _00105_ clknet_leaf_119_wb_clk_i cpu.regs\[13\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09726__C _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10141_ _00040_ clknet_leaf_108_wb_clk_i cpu.br_rel_dest\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10072_ _01941_ _05012_ _05013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_7_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08358__B _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_74_Left_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_qcpu_113 io_oeb[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_57_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_qcpu_102 io_oeb[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_97_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06018__A1 _01492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06018__B2 _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10408_ _00303_ clknet_leaf_56_wb_clk_i cpu.orig_IO_addr_buff\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10339_ _00234_ clknet_leaf_61_wb_clk_i cpu.spi.counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05736__I _01195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07369__I1 _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05880_ cpu.br_rel_dest\[1\] _01363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_108_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07550_ _02930_ _02933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05395__I3 cpu.regs\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06501_ _01717_ _01978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08494__A2 _03626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09220_ _04241_ _04242_ _04243_ _04244_ _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_07481_ _02887_ _02888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06432_ _01901_ _01910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09151_ cpu.ROM_addr_buff\[4\] _04179_ _04188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_60_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09443__A1 _04456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06363_ _01838_ _01840_ _01841_ _01842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_17_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08102_ _03365_ _00239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_83_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07398__I _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09082_ _04133_ cpu.ROM_addr_buff\[2\] _04134_ _04135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05314_ cpu.regs\[8\]\[2\] cpu.regs\[9\]\[2\] cpu.regs\[10\]\[2\] cpu.regs\[11\]\[2\]
+ _00801_ _00574_ _00823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08033_ cpu.uart.dout\[1\] _03301_ _03304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06294_ _01773_ _00017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05245_ _00753_ _00758_ _00759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05176_ _00691_ _00692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07757__A1 _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09984_ cpu.PORTA_DDR\[6\] _04926_ _04933_ _04931_ _04934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05232__A2 _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08935_ _04013_ _00418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_4_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input21_I io_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08957__I _00903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08866_ _03137_ _03953_ _03954_ _03962_ _03963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_98_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07817_ _02517_ _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08797_ _02703_ _03895_ _03905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07748_ _00790_ _03057_ _03058_ _03059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07679_ _02975_ _03011_ _03013_ _00162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09418_ cpu.orig_PC\[4\] _04437_ _04438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10690_ net49 net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09349_ _04370_ _04332_ _04371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05310__I3 cpu.regs\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06420__A1 _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10124_ _00023_ clknet_4_8_0_wb_clk_i cpu.regs\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_101_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10055_ _04987_ _04994_ _04996_ _03366_ _00555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_82_Left_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06487__A1 _01862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_91_Left_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09425__A1 _02334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05301__I3 cpu.regs\[11\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06981_ _02447_ _02449_ _02452_ _02453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_111_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_47_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_47_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08777__I _03275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08720_ _02723_ _03844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05932_ _01412_ _01413_ _01414_ _01415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08164__A1 _03335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08651_ _03792_ _03791_ cpu.pwm_counter\[5\] _03794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05863_ _01141_ _01143_ _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07602_ _02556_ _02960_ _00136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_37_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08582_ _03719_ _03720_ _03738_ _03745_ _03746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05794_ _01277_ _01278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_88_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08467__A2 _03636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07533_ _02920_ _02915_ _02921_ _00108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07464_ _02872_ _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06415_ _01688_ _01278_ _01721_ _01893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09203_ _00846_ _01344_ _01939_ _04228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_97_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09134_ _00689_ _00690_ _04168_ _04175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09416__A1 _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07395_ _02810_ _00081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_115_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06346_ _00612_ _01825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_17_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09065_ _02508_ _04116_ _04122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06277_ _01724_ _01672_ _01745_ _01757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_08016_ cpu.spi.data_in_buff\[2\] _03291_ _03287_ cpu.spi.data_in_buff\[3\] _03293_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05228_ cpu.uart.busy cpu.spi.busy _00719_ _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_8_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05205__A2 cpu.spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05159_ cpu.IO_addr_buff\[7\] cpu.IO_addr_buff\[6\] cpu.IO_addr_buff\[5\] _00676_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_40_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09967_ _04921_ _00542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08918_ _02735_ _03997_ _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09292__B _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09898_ _04868_ _04870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08849_ _03170_ _03946_ _03948_ _03949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09655__A1 _00604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09311__I _04309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10107_ _05041_ _00562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10038_ _04973_ _04980_ _02420_ _04981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08146__A1 _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09894__A1 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09646__A1 _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07121__A2 _02583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06200_ _01159_ _01681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07180_ _02631_ _02616_ _02632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06131_ _01181_ _01612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_14_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06062_ _01541_ _01543_ _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_113_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09821_ _04807_ _04808_ _00509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09752_ _04739_ _04737_ _04752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06964_ cpu.startup_cycle\[4\] _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08703_ _03827_ _03831_ _00368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09885__A1 _04045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09683_ cpu.last_addr\[5\] _04189_ _04677_ _04693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05915_ cpu.timer_div\[1\] _01397_ _01182_ _01398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_55_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06895_ _00603_ _02370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07344__C _02763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08634_ cpu.pwm_counter\[0\] _03782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05846_ _01329_ _01330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08565_ _03726_ _03727_ _03728_ _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05777_ _01260_ _01261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07516_ _02908_ _00104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08496_ _02046_ _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07447_ _02842_ _02854_ _02855_ _02815_ _02857_ _02858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_64_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08970__I _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07378_ _01582_ _02764_ _02794_ _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09117_ cpu.regs\[3\]\[3\] _03082_ _04150_ _04161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06329_ cpu.timer_top\[13\] _01404_ _01621_ _01807_ _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_44_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09048_ cpu.IO_addr_buff\[6\] _04097_ _04108_ _04100_ _04109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06623__A1 _00829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09306__I _04327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output52_I net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07726__I1 cpu.regs\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10656_ _00550_ clknet_leaf_77_wb_clk_i net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_36_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05665__A2 _01071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10587_ _00481_ clknet_leaf_98_wb_clk_i cpu.PC\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_10_Left_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08119__A1 _02621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05276__S1 _00786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09867__A1 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_2_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05700_ _01183_ _01184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_78_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06680_ _02152_ _02155_ _02156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05631_ _00702_ _00717_ _00744_ _01071_ _01115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_116_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08350_ _03561_ _03562_ _00284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08276__B _03505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05562_ _01045_ _01046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07301_ _02731_ _02732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08281_ _03499_ _03508_ _03509_ _00268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06508__C _01122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05493_ _00928_ _00951_ _00979_ _00980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10097__I _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09886__I _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07232_ _02673_ _02659_ _02674_ _02676_ _02677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_27_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07163_ _02608_ _02613_ _02617_ _02518_ _02618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_26_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06114_ _01091_ _01595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07094_ _02558_ _02559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_14_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_62_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_62_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06045_ _01173_ _01526_ _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_74_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09804_ _04780_ _04795_ _04796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07996_ _03190_ _03272_ _03268_ _03278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_5_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06947_ _02418_ _02419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09735_ _02487_ _02481_ _04739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09666_ cpu.last_addr\[2\] cpu.last_addr\[1\] cpu.last_addr\[0\] _04676_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__08965__I _00952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08530__A1 _02755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06878_ _02045_ _02062_ _02350_ _02353_ _02354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08617_ _03756_ _03770_ _03771_ _00342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09597_ _02047_ _00930_ _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05829_ _01299_ _01313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09086__A2 _00832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08548_ _03711_ cpu.toggle_top\[13\] cpu.toggle_top\[12\] _03708_ _03712_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_08479_ _03658_ _03660_ _03650_ _00315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_65_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10510_ _00405_ clknet_leaf_53_wb_clk_i cpu.spi.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10441_ _00336_ clknet_leaf_6_wb_clk_i cpu.toggle_ctr\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_45_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10372_ _00267_ clknet_leaf_63_wb_clk_i cpu.uart.data_buff\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07021__A1 _00668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09480__B _04417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_46_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10639_ _00533_ clknet_leaf_68_wb_clk_i cpu.PORTB_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07850_ cpu.timer_top\[12\] _03136_ _03148_ _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_85_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06801_ _02276_ _02246_ _02277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07781_ _02557_ _03085_ _03088_ _03052_ _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xinput3 io_in[11] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09520_ _04334_ _04526_ _04535_ _04345_ _04536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06732_ _02193_ _02194_ _02208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_36_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_108_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08512__A1 _02735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09451_ _02370_ _04409_ _04469_ _04470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06663_ _00619_ _00975_ _02138_ _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08402_ net17 _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_05614_ _01093_ _01097_ _01098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09382_ _01135_ _04399_ _04402_ _00767_ _04403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_47_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06594_ _02068_ _02069_ _02070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08333_ cpu.uart.receive_div_counter\[2\] cpu.uart.receive_div_counter\[1\] cpu.uart.receive_div_counter\[0\]
+ _03548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_86_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05545_ _01028_ _01029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08264_ cpu.uart.data_buff\[4\] _03491_ _03495_ _03496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_50_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06826__A1 _00907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05476_ _00959_ _00962_ _00871_ _00963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08195_ cpu.uart.div_counter\[13\] _03439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07215_ _01004_ _02661_ _02662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07146_ _01774_ _02599_ _02604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07251__A1 _02692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07077_ _02543_ _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_112_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06028_ cpu.spi.dout\[2\] _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05101__I1 _00619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09718_ _04718_ _04717_ _04724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07979_ _03184_ _03181_ _03261_ _03264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_58_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07813__B _03112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08503__A1 _02621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09649_ _00734_ _00764_ _04432_ _04659_ _04660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_2_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07104__I _02568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10424_ _00319_ clknet_leaf_87_wb_clk_i cpu.orig_PC\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09231__A2 _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10355_ _00250_ clknet_leaf_34_wb_clk_i cpu.uart.div_counter\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_94_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10286_ _00181_ clknet_leaf_112_wb_clk_i cpu.regs\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05294__I cpu.regs\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_2_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05330_ _00581_ _00837_ _00838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05261_ _00682_ _00775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_113_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07000_ _02471_ _00729_ _02472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_72_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05192_ cpu.instr_buff\[15\] _00707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_52_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09222__A2 _02270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_102_Left_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08951_ _04025_ _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07902_ _00775_ _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_08882_ _03944_ _03975_ _03976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07833_ cpu.TIE _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XPHY_EDGE_ROW_81_Right_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_55_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07764_ _02328_ _02216_ net117 _03073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_79_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09503_ _04368_ _04502_ _04519_ _04374_ _04375_ _04520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_06715_ _00618_ _00907_ _02191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07695_ _03021_ _03022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_69_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09434_ cpu.orig_PC\[5\] _04437_ _04453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06646_ cpu.regs\[1\]\[2\] _00996_ _02122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_111_Left_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09365_ _04385_ _04386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06577_ cpu.PC\[2\] _02053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08316_ cpu.uart.receive_buff\[6\] _03522_ _03530_ cpu.uart.receive_buff\[7\] _03535_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05528_ _00708_ _00651_ _01010_ _01012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_47_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09296_ _04287_ _04319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08247_ _02707_ _03465_ _03482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_90_Right_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05459_ _00880_ _00946_ _00947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08178_ cpu.uart.div_counter\[9\] _03388_ _03425_ _03398_ _03426_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_70_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07594__I _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07129_ _01015_ _02586_ _02591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08972__A1 _04041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10140_ _00039_ clknet_leaf_108_wb_clk_i cpu.br_rel_dest\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10071_ _01942_ _05011_ _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08724__A1 cpu.timer_top\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05842__I _01325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_qcpu_114 io_oeb[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xwrapped_qcpu_103 io_oeb[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_93_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10536__CLK clknet_leaf_18_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05289__I _00799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06018__A2 _01035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07215__A1 _01004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10407_ _00302_ clknet_leaf_55_wb_clk_i cpu.orig_IO_addr_buff\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10338_ _00233_ clknet_leaf_64_wb_clk_i net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_119_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_119_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10269_ _00164_ clknet_leaf_110_wb_clk_i cpu.regs\[5\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05529__A1 _00654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_105_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09140__A1 cpu.ROM_addr_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07480_ _02886_ _02887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06500_ net33 _01976_ _01580_ _01977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09691__A2 cpu.ROM_addr_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08284__B _03505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06431_ _01826_ _00999_ _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09150_ _00777_ _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_60_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06362_ _01450_ _01818_ _01841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08101_ _03200_ _03364_ _03365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09081_ _04022_ _04134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06293_ _01772_ cpu.regs\[9\]\[4\] _01681_ _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05313_ _00586_ _00821_ _00822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08032_ cpu.uart.receive_buff\[1\] _02881_ _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05244_ _00757_ _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05199__I cpu.base_address\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05175_ _00690_ _00667_ _00691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08954__A1 _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09983_ _02646_ _04927_ _04933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10054__B net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08934_ cpu.timer_div\[5\] _03996_ _04012_ _04003_ _04013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_110_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_4_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08865_ _00978_ _03955_ _03962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07816_ _01981_ _03104_ _03115_ _00197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_74_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08796_ _03857_ _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input14_I io_in[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07747_ _02523_ _02535_ _02022_ _03052_ _03058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_67_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07678_ cpu.regs\[5\]\[0\] _03012_ _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05379__S0 _00864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09417_ _04239_ _04437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06629_ _02103_ _02104_ _02105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09348_ _04319_ _04370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09279_ _02512_ _04301_ _04302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09198__A1 _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06420__A2 _01784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10123_ _00022_ clknet_leaf_102_wb_clk_i cpu.regs\[2\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10054_ _04987_ _04995_ net77 _04996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_4_7_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08936__A1 _02755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06980_ _02028_ _02033_ _02451_ _02452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA_input6_I io_in[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09382__C _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05931_ _01269_ _01414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08650_ _03781_ _03793_ _00353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05862_ _01345_ _01346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06578__I cpu.PC\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07911__A2 cpu.spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07601_ _02962_ _00135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_37_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_87_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_87_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05793_ _01276_ _01277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08581_ _03712_ _03716_ _03740_ _03744_ _03745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_88_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_16_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_16_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_9_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07532_ cpu.regs\[12\]\[2\] _02916_ _02921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07463_ _00768_ _02872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09202_ _04226_ _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06414_ _01416_ _01863_ _01891_ _01589_ _01892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09133_ cpu.last_addr\[0\] _04174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07394_ _02809_ _02093_ _02775_ _02810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06345_ _01326_ _01823_ _01824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09064_ _00932_ _04121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06276_ _01753_ _01755_ _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_32_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08015_ _03289_ _03292_ _00219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05227_ _00740_ _00718_ _00658_ _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_4_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08927__A1 cpu.timer_div\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05158_ cpu.IO_addr_buff\[4\] _00675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_8_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09966_ cpu.PORTA_DDR\[1\] _04915_ _04919_ _04920_ _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05089_ cpu.regs\[8\]\[5\] cpu.regs\[9\]\[5\] cpu.regs\[10\]\[5\] cpu.regs\[11\]\[5\]
+ _00572_ _00599_ _00609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_0_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09897_ _04868_ _04869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_85_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08917_ _03995_ _04000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08848_ _02707_ _03947_ _03948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06166__A1 _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08779_ _03887_ _03890_ _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08918__A1 _02735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10106_ _01771_ cpu.regs\[15\]\[4\] _05034_ _05041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10037_ _04736_ _04976_ _04979_ _04980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_98_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08562__B _01176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06880__A2 _02354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08082__B2 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06130_ _01610_ _01368_ _01396_ _01611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_53_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06061_ _01364_ _01454_ _01542_ _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_113_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09820_ _02417_ _04769_ _03474_ _04808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08788__I _03864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09751_ _02436_ _04750_ _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06963_ cpu.startup_cycle\[4\] _02430_ _02434_ _02435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__06302__S _00851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05914_ _01396_ _01397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08702_ cpu.timer_div_counter\[3\] _03829_ _03831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09334__A1 _02593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09682_ _04197_ cpu.ROM_addr_buff\[7\] _04678_ _04692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__06148__A1 _00966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06894_ _02338_ _02341_ _02369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08633_ _03551_ _03781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05845_ _01313_ _01328_ _01329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__06101__I _01582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08564_ cpu.toggle_ctr\[3\] _01590_ _01485_ cpu.toggle_ctr\[2\] _03728_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05776_ _00703_ _01021_ _01259_ _01260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__09412__I _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07515_ _01935_ cpu.regs\[13\]\[6\] _02898_ _02908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08495_ _03670_ _03671_ _03667_ _00320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_71_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07446_ cpu.uart.receive_div_counter\[7\] _02856_ _02622_ _02836_ _02857_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_91_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07377_ _02524_ _02790_ _02793_ _02531_ _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09116_ _04160_ _00452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_79_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06328_ _01786_ _01245_ _01805_ _01806_ _01247_ _01807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_45_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09047_ _04079_ _04106_ _04107_ _04108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_20_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06259_ _01730_ _01738_ _01739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09573__A1 _04121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09949_ _02502_ _04908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06139__A1 cpu.timer_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_36_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09322__I _04313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06311__A1 net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10655_ _00549_ clknet_leaf_77_wb_clk_i cpu.ROM_spi_mode vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_24_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09100__I1 _04147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06681__I _00906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10586_ _00480_ clknet_leaf_93_wb_clk_i cpu.PC\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_75_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07878__A1 _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05630_ _01113_ _01114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_59_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09619__A2 _01155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05561_ _01044_ _01040_ _01045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07300_ _01202_ _02730_ _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08280_ cpu.uart.data_buff\[8\] _03497_ _03505_ _03509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05492_ _00971_ _00978_ _00939_ _00979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07231_ _02675_ _02661_ _02676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07162_ _02615_ _02616_ _02617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06113_ net82 _01208_ _01594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07093_ _02050_ _02558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06044_ _00779_ _01171_ _01524_ _01525_ _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_74_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08311__I _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09803_ cpu.ROM_spi_dat_out\[3\] _04779_ _04785_ _04795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07995_ _03274_ _03277_ _00214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06946_ _02415_ _02416_ _02417_ _00660_ _02418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_09734_ _04731_ _04737_ _02481_ _02488_ _04738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xclkbuf_leaf_31_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_31_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_66_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09665_ _02030_ _04674_ _04675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07869__B2 cpu.timer_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07869__A1 cpu.timer_top\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06877_ _02351_ _02352_ _02353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05828_ _01305_ _01311_ _01262_ _01312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08616_ _03704_ _03739_ _03767_ _03771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_09596_ _00971_ _04399_ _04608_ _04396_ _04609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05759_ _01242_ _01243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_25_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08547_ cpu.toggle_ctr\[13\] _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08981__I _04002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08478_ cpu.orig_PC\[6\] _03659_ _03660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_53_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07429_ _02820_ _02827_ _02834_ _02839_ _02840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_80_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10440_ _00335_ clknet_leaf_7_wb_clk_i cpu.toggle_ctr\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09094__I0 _00604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10371_ _00266_ clknet_leaf_63_wb_clk_i cpu.uart.data_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_88_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06532__A1 _01419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10092__A1 net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10638_ _00532_ clknet_leaf_68_wb_clk_i net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_106_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10569_ _00463_ clknet_leaf_83_wb_clk_i cpu.last_addr\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05271__A1 _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09537__A1 _03045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06800_ _02243_ _00965_ _02276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07780_ _03086_ _03087_ _03088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput4 io_in[12] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06731_ _02205_ _02206_ _02207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_108_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09450_ _04410_ _04452_ _04469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08401_ _03601_ _03602_ _03600_ _00295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06662_ _02130_ _02131_ _02138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05490__I _00976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05613_ _01033_ _01096_ _01097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09381_ _04399_ _04401_ _04402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06593_ _02066_ _02067_ _02069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08332_ _03547_ _00281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09897__I _04868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05544_ _00675_ _00676_ _01028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08263_ _03231_ _03486_ _03495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_50_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07214_ _02658_ _02661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05475_ _00960_ _00961_ _00850_ _00962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08194_ _03436_ _03438_ _00252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07145_ _02580_ _02600_ _02601_ _02603_ _00038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_42_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07076_ _02534_ _02535_ _02541_ _02542_ _02543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_100_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06027_ _01507_ _01508_ _01187_ _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__05101__I2 cpu.regs\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07978_ _03181_ _03261_ _03263_ _03097_ _00211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09717_ cpu.mem_cycle\[4\] _04718_ _04717_ _04723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_58_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06929_ net19 _02042_ _02403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08503__A2 _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09648_ _00763_ _04649_ _04658_ _04659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_2_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09579_ _01297_ _01313_ _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10074__A1 _04121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10423_ _00318_ clknet_leaf_87_wb_clk_i cpu.orig_PC\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10354_ _00249_ clknet_leaf_32_wb_clk_i cpu.uart.div_counter\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09519__A1 _04530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10285_ _00180_ clknet_leaf_109_wb_clk_i cpu.regs\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07790__I _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08819__C _03920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10065__A1 _01419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05260_ net18 _00695_ _00728_ _00774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05492__A1 _00971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05191_ cpu.base_address\[5\] _00706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08950_ _01052_ _01185_ _02611_ _04025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_71_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07901_ _03198_ _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08881_ _03933_ _03946_ _03974_ _03975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09930__A1 _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07832_ _03130_ _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06744__A1 _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09502_ _02375_ _04369_ _04518_ _04519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07763_ _03070_ _03071_ _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_55_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06714_ _02188_ _02189_ _02190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07694_ _02911_ _02977_ _03021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_69_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09433_ _04451_ _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06645_ cpu.regs\[1\]\[3\] _00963_ _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09364_ _02052_ _04384_ _04385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08315_ _03532_ _03534_ _00277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10056__A1 _00653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06576_ cpu.PC\[3\] _02052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_117_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09997__A1 _03822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09295_ _04315_ _04317_ _04318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05527_ _00711_ _01010_ _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_28_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08246_ _03471_ _03481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05458_ cpu.regs\[0\]\[3\] _00829_ cpu.regs\[2\]\[3\] cpu.regs\[3\]\[3\] _00882_
+ _00884_ _00946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08177_ cpu.uart.div_counter\[9\] _03421_ _03417_ _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_7_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07128_ _02505_ _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09213__A3 _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05389_ _00849_ _00878_ _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_30_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07059_ _02391_ _02526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_7_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10070_ _01943_ _01946_ _05011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09921__A1 _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_102_Right_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07783__I0 _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_qcpu_104 io_oeb[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_85_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08660__A1 _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10406_ _00301_ clknet_leaf_56_wb_clk_i cpu.orig_IO_addr_buff\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10337_ _00232_ clknet_leaf_44_wb_clk_i cpu.uart.dout\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10268_ _00163_ clknet_leaf_13_wb_clk_i cpu.regs\[5\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10199_ _00094_ clknet_leaf_120_wb_clk_i cpu.regs\[14\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05529__A2 _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07151__A1 _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06430_ _01435_ _01907_ _01908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09979__A1 _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06361_ _01687_ _01337_ _01839_ _01335_ _00716_ _01840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_32_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08100_ _03362_ _03363_ _03364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09080_ _00818_ _02789_ _04130_ _04133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_60_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06292_ _01771_ _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05312_ cpu.regs\[12\]\[2\] cpu.regs\[13\]\[2\] cpu.regs\[14\]\[2\] cpu.regs\[15\]\[2\]
+ _00801_ _00802_ _00821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08031_ _01223_ _03301_ _03302_ _00225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05465__A1 _00928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05243_ _00756_ _00757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07695__I _03021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05174_ _00666_ _00690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05217__A1 _00668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09982_ _04932_ _00546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_110_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08933_ _02750_ _04009_ _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08864_ _03961_ _00399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07815_ cpu.spi.data_in_buff\[7\] _03101_ _03112_ _03115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08795_ _03903_ _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07746_ _01358_ _02407_ _03054_ _03056_ _03057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_79_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09416_ _00752_ _04435_ _04436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07142__A1 _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07677_ _03009_ _03012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05379__S1 _00865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08890__A1 _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06628_ _02088_ _02089_ _02104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07693__A2 _03012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06559_ cpu.mem_cycle\[3\] _02035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_81_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09347_ _04288_ _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09278_ _00742_ _00757_ _04301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_62_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08229_ _03360_ _03463_ _03466_ _03456_ _03467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_90_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08945__A2 _04020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output75_I net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10122_ _00021_ clknet_leaf_102_wb_clk_i cpu.regs\[2\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10053_ _02456_ _04988_ _04993_ _04773_ _04995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09325__I _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07133__A1 _02593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05930_ _00878_ _01261_ _01413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05861_ _00843_ _01344_ _01345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08580_ _03706_ _03702_ _03743_ _03710_ _03744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_07600_ _02365_ _02959_ _02912_ _02962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__06175__A2 _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09649__B1 _04432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05792_ _01263_ _01072_ _01276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07531_ _01583_ _02920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_66_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07462_ _02868_ _02869_ _02871_ _00087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10110__S _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09201_ _00723_ _03624_ _04226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_63_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06413_ _01269_ _01890_ _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_45_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07393_ _01678_ _02764_ _02808_ _02809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09132_ cpu.ROM_addr_buff\[0\] _04172_ _04173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_56_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_56_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_56_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06344_ _01819_ _01821_ _01823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05438__A1 _00715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09063_ _04120_ _00439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06275_ _01640_ _01737_ _01754_ _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08014_ cpu.spi.data_in_buff\[1\] _03291_ _03287_ cpu.spi.data_in_buff\[2\] _03292_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05226_ _00650_ _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_8_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05157_ cpu.IO_addr_buff\[3\] _00674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06938__A1 _02410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09965_ _02502_ _04920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05088_ _00587_ _00607_ _00608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08916_ _03822_ _03999_ _00413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09896_ _01046_ _04842_ _04868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08847_ _03945_ _03947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08984__I _02651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08778_ cpu.timer_capture\[4\] _03888_ _03889_ _03890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05913__A2 _01395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_26_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07729_ _03042_ _00183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07115__A1 _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10671_ _00565_ clknet_leaf_1_wb_clk_i cpu.regs\[15\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06477__I0 _01781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06929__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_65_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10105_ _01679_ _05035_ _05040_ _00561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10036_ _04952_ _04978_ _04979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09343__A2 _00757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07657__A2 _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06060_ _01427_ _01428_ _01542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_113_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09031__A1 _01587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_103_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_103_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09750_ _04749_ _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06962_ _02432_ _02433_ _00662_ _02434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08701_ _03826_ _03829_ _03830_ _00367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09681_ cpu.last_addr\[8\] cpu.ROM_addr_buff\[8\] _04679_ _04691_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_05913_ _00673_ _01395_ _01094_ _01059_ _01396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__09334__A2 _04349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08632_ _03753_ _03780_ _00348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06893_ _02345_ _02348_ _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08542__B1 _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05844_ _00928_ cpu.base_address\[2\] _01328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08563_ cpu.toggle_ctr\[2\] _01485_ _01410_ cpu.toggle_ctr\[1\] _03727_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_05775_ _01018_ _01020_ _01259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_76_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08494_ cpu.orig_PC\[11\] _03626_ _03671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07514_ _02907_ _00103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07445_ _02650_ _02856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_92_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07213__I _02655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08753__B _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07376_ _02526_ _02313_ _02792_ _02564_ _02793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_09115_ _04158_ cpu.ROM_addr_buff\[10\] _04159_ _04160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09270__A1 _00724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06327_ cpu.timer_capture\[13\] _01233_ _01239_ _01806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_45_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09046_ _01860_ _04058_ _04107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06258_ _01633_ _00977_ _01658_ _01738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06084__A1 _01144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05209_ _00723_ _00724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08979__I _02698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06189_ _01575_ _01661_ _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09573__A2 _04349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09948_ _04045_ _04904_ _04907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09879_ _04855_ _00520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_output38_I net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07123__I _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10654_ _00548_ clknet_leaf_58_wb_clk_i cpu.PORTA_DDR\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09261__A1 _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10585_ _00479_ clknet_leaf_93_wb_clk_i cpu.PC\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06075__A1 _01296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_1_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_1_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09013__A1 _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09564__A2 _00929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10019_ _04961_ _04962_ _04953_ _04963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07878__A2 _03176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05560_ _00644_ _01043_ _01044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_59_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05491_ _00977_ _00978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07230_ _00937_ _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07161_ _02612_ _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09252__A1 _00734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06112_ _01207_ _01593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_41_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07092_ _02522_ _02557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_112_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06043_ _00902_ _01292_ _01293_ _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09802_ _04771_ _04793_ _04794_ _00504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07994_ _03272_ _03268_ _03276_ _03277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06945_ cpu.ROM_spi_cycle\[0\] _02417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06112__I _01207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09733_ _04732_ _02427_ _02424_ _04736_ _04737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_09664_ _02461_ _02582_ _04674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06876_ _02149_ _02331_ _02349_ _02352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_96_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09595_ _04399_ _04607_ _04608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08615_ _03739_ _03767_ _03704_ _03770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05827_ _01306_ _01310_ _01311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_71_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_71_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_82_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05758_ _01094_ _01241_ _01242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08546_ _03708_ cpu.toggle_top\[12\] cpu.toggle_top\[11\] _03709_ _03710_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_92_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08477_ _03625_ _03659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09491__A1 _04456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05689_ _01172_ _01173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07428_ _02835_ _02818_ _02825_ _02824_ _02838_ _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_64_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07359_ _02299_ _02309_ _02777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09094__I1 _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10370_ _00265_ clknet_leaf_66_wb_clk_i cpu.uart.data_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09029_ cpu.orig_IO_addr_buff\[3\] _04091_ _04092_ _00978_ _04093_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07557__A1 cpu.regs\[11\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07281__C _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09333__I _04313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09489__B _04455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10637_ _00531_ clknet_leaf_66_wb_clk_i net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_3_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_116_Right_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10568_ _00462_ clknet_leaf_82_wb_clk_i cpu.last_addr\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08840__C _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10499_ _00394_ clknet_leaf_8_wb_clk_i cpu.timer\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09537__A2 _04500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput5 io_in[13] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06730_ _02172_ _02173_ _02206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06771__A2 _00966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06661_ _00949_ _02130_ _02131_ _02137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_36_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08400_ _02846_ _02850_ _03558_ _03593_ _03602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_78_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05612_ _01095_ _01096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06088__B _01326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07720__A1 cpu.regs\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09380_ _02052_ _04068_ _04400_ _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06592_ _02066_ _02067_ _02068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08331_ _03116_ _03546_ _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05543_ _01026_ _01027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08262_ _03481_ _03493_ _03494_ _00264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_52_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05474_ cpu.regs\[0\]\[4\] cpu.regs\[1\]\[4\] cpu.regs\[2\]\[4\] cpu.regs\[3\]\[4\]
+ _00956_ _00957_ _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_22_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07213_ _02655_ _02660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08193_ _03323_ _03434_ _03437_ _03438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06039__A1 _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07144_ _02602_ _02603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07075_ _02520_ _02542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06026_ cpu.spi.divisor\[2\] _01189_ _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07977_ cpu.spi.div_counter\[2\] _03252_ _03262_ _03259_ _03263_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09716_ _04722_ _00490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_58_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06928_ _02392_ _02401_ _02359_ _02402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06777__I _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09647_ _03674_ _00763_ _04658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06859_ _02334_ _01289_ _02081_ _02335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_2_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09578_ _04382_ _04577_ _04591_ _04406_ _04592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_93_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08925__C _04006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08529_ _03695_ _00330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_37_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05325__I0 cpu.regs\[0\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09216__A1 _02593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10422_ _00317_ clknet_leaf_86_wb_clk_i cpu.orig_PC\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07078__I0 _02334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10353_ _00248_ clknet_leaf_32_wb_clk_i cpu.uart.div_counter\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_33_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05856__I _01309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10284_ _00179_ clknet_leaf_109_wb_clk_i cpu.regs\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05800__I1 cpu.regs\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05492__A2 _00978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05190_ cpu.base_address\[4\] _00705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07769__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06441__A1 _01331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_71_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06441__B2 _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07900_ _03197_ _03198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08880_ _03947_ _02698_ _03974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07831_ _03117_ _03118_ _03126_ _03129_ _03130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XPHY_EDGE_ROW_16_Left_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09501_ _04370_ _04502_ _04518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07762_ _02060_ _03071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08497__A2 _03609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06713_ _00589_ _00934_ _02189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07693_ _02992_ _03012_ _03020_ _00169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09432_ _02549_ _04449_ _04450_ _04451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06644_ _02065_ _02119_ _02120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_82_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06575_ cpu.PC\[4\] _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_19_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09363_ _02053_ _02054_ cpu.PC\[0\] _04384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08314_ cpu.uart.receive_buff\[5\] _03522_ _03530_ cpu.uart.receive_buff\[6\] _03534_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05526_ _01009_ _01010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__05450__B _00912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09446__A1 _01774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09294_ cpu.orig_PC\[1\] _04267_ _04316_ _00749_ _04317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_25_Left_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08245_ _03480_ _00261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05457_ _00887_ _00944_ _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08176_ _03421_ _03417_ _03424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05388_ _00877_ _00878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_42_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07127_ _02580_ _02587_ _02588_ _02589_ _00034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_112_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05676__I _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07058_ _02051_ _02055_ _02525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06009_ cpu.uart.divisor\[2\] _01383_ _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_7_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_34_Left_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07932__A1 _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07783__I1 _03090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_qcpu_105 io_oeb[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_97_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_43_Left_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07131__I _02508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10405_ _00300_ clknet_leaf_17_wb_clk_i cpu.orig_IO_addr_buff\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08412__A2 _03611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10336_ _00231_ clknet_leaf_43_wb_clk_i cpu.uart.dout\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_52_Left_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10267_ _00162_ clknet_leaf_13_wb_clk_i cpu.regs\[5\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07923__A1 _03201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10198_ _00093_ clknet_leaf_1_wb_clk_i cpu.regs\[14\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05085__S1 _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_61_Left_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07151__A2 _02598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06360_ _01826_ _01686_ _01839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_17_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06291_ _01770_ _01771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05311_ _00815_ _00819_ _00580_ _00820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput30 sram_out[4] net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08030_ cpu.uart.receive_buff\[0\] _03300_ _03245_ _03302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05242_ _00754_ _00755_ _00746_ _00756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_25_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_116_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_5_0_wb_clk_i clknet_0_wb_clk_i clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_05173_ _00688_ _00689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08403__A2 _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10108__S _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09981_ cpu.PORTA_DDR\[5\] _04926_ _04930_ _04931_ _04932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_12_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08932_ _04011_ _00417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08863_ cpu.timer_capture\[10\] _03943_ _03960_ _03951_ _03961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07814_ _01865_ _03104_ _03114_ _00196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08794_ cpu.timer_capture\[7\] _03870_ _03902_ _03820_ _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_clkbuf_leaf_16_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07745_ net1 _03055_ _02406_ _03056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09415_ _01683_ _04430_ _04433_ _04434_ _04435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07676_ _03010_ _03011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_94_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06627_ _02100_ _02101_ _02102_ _02103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06558_ _02033_ _02034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09346_ _02512_ _04368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_75_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09277_ _04299_ _04300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05509_ _00993_ _00994_ _00850_ _00995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06489_ net97 _01965_ _01966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_35_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08228_ _03454_ _03465_ _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_35_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08159_ _03337_ _03407_ _03411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_101_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06405__A1 cpu.timer_capture\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_55_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10121_ _00020_ clknet_leaf_120_wb_clk_i cpu.regs\[9\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output68_I net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10052_ _04953_ _02459_ _04993_ _04994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07126__I _00686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09658__A1 _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07133__A2 _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_94_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10319_ _00214_ clknet_leaf_50_wb_clk_i cpu.spi.div_counter\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08149__A1 _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05860_ _00712_ _01344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__09649__A1 _00734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05791_ _01266_ _01271_ _01274_ _00902_ _01275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_37_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07530_ _02918_ _02915_ _02919_ _00107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_66_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07461_ _02870_ _02871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09200_ _04222_ _04225_ _00471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10478__CLK clknet_leaf_18_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06412_ _01687_ _01717_ _01889_ _01175_ _01890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_45_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06883__A1 _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07392_ _02798_ _02801_ _02807_ _02531_ _02808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09131_ _04171_ _04172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06343_ _01819_ _01821_ _01822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_72_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05438__A2 _00912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09062_ _00847_ _04115_ _04119_ _04050_ _04120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_44_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_96_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_96_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06274_ _01640_ _01743_ _01754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08013_ _03198_ _03291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05225_ _00726_ _00738_ _00739_ _00010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_25_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_25_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_8_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05156_ _00672_ _00673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_69_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06938__A2 _02359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09964_ _00904_ _04916_ _04919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05087_ cpu.regs\[12\]\[5\] cpu.regs\[13\]\[5\] cpu.regs\[14\]\[5\] cpu.regs\[15\]\[5\]
+ _00572_ _00576_ _00607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_09895_ _04867_ _00524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09888__A1 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08915_ cpu.timer_div\[0\] _03996_ _03998_ _03999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08846_ _03945_ _03946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_99_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08777_ _03275_ _03889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05913__A3 _01094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05989_ _01455_ _01471_ _01472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_95_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07728_ _03004_ cpu.regs\[3\]\[5\] _03033_ _03042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07659_ cpu.regs\[6\]\[2\] _02997_ _03000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10670_ _00564_ clknet_leaf_121_wb_clk_i cpu.regs\[15\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09329_ _04055_ _04351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_11_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07051__A1 _02513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09336__I _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10104_ cpu.regs\[15\]\[3\] _05034_ _05040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10035_ _04974_ _04977_ _02426_ _04978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09103__I0 cpu.regs\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05840__A2 _01322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07475__B _02882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06961_ cpu.startup_cycle\[2\] _02433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08790__A1 cpu.timer_capture\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08700_ cpu.timer_div_counter\[0\] cpu.timer_div_counter\[1\] cpu.timer_div_counter\[2\]
+ _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09680_ cpu.last_addr\[9\] cpu.ROM_addr_buff\[9\] _04689_ _04690_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_05912_ _00647_ _01395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06892_ cpu.PC\[13\] _02366_ _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_08631_ cpu.toggle_ctr\[14\] _03778_ cpu.toggle_ctr\[15\] _03780_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05843_ _01168_ _01310_ _01327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08562_ cpu.toggle_ctr\[1\] _01410_ _01176_ cpu.toggle_ctr\[0\] _03726_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05774_ _01256_ _01257_ _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08493_ _03082_ _03611_ _03670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07513_ _01858_ cpu.regs\[13\]\[5\] _02898_ _02907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10101__A1 _01481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07444_ cpu.uart.receive_div_counter\[6\] _02855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07375_ _02777_ _02791_ _02792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09114_ _04022_ _04159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_79_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06326_ cpu.timer_capture\[5\] _01690_ _01802_ _01804_ _01243_ _01805_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_60_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07281__A1 _02627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09045_ cpu.orig_IO_addr_buff\[6\] _04075_ _04076_ _01957_ _04106_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06257_ _01729_ _01736_ _01737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05208_ _00722_ _00723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06188_ _01637_ _01667_ _01669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_111_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05139_ _00654_ _00655_ _00656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XPHY_EDGE_ROW_8_Left_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09947_ _04906_ _00537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09878_ net62 _04844_ _04854_ _04849_ _04855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08829_ cpu.timer_capture\[13\] _03913_ _03914_ _03932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05898__A2 _01035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10653_ _00547_ clknet_leaf_59_wb_clk_i cpu.PORTA_DDR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_36_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07279__C _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10584_ _00478_ clknet_4_9_0_wb_clk_i cpu.PC\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09066__I _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08524__A1 _02746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07515__S _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10018_ cpu.ROM_addr_buff\[2\] _04950_ _02484_ cpu.ROM_addr_buff\[10\] _04962_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_47_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07314__I _00952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05490_ _00976_ _00977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_116_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07160_ _02614_ _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_54_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06111_ cpu.uart.divisor\[3\] _01592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_81_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07091_ _01933_ _02556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06042_ _01414_ _01522_ _01523_ _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_74_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09801_ cpu.ROM_spi_dat_out\[3\] _04772_ _02715_ _04794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09732_ _04735_ _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07993_ _03275_ _03276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__05121__S0 _00630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06944_ cpu.ROM_spi_cycle\[1\] _02416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08515__A1 _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09663_ _04672_ _04673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06875_ _02043_ _02351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09594_ _03081_ _04484_ _04606_ _04607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08614_ _03751_ _03769_ _00341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05826_ _00800_ _01309_ _01310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_08545_ cpu.toggle_ctr\[11\] _03709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_85_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05757_ _01061_ _01185_ _01241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08476_ _02559_ _03657_ _03658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05688_ _01139_ _01172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07427_ _02836_ cpu.uart.divisor\[1\] _02837_ cpu.uart.receive_div_counter\[0\] _02838_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_64_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_40_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_40_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07358_ _02776_ _00078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05679__I _01162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06309_ cpu.uart.divisor\[5\] _01788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__07254__A1 cpu.timer_capture\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07289_ _00776_ _02723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_33_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09028_ _04063_ _04092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07006__A1 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output50_I net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10636_ _00530_ clknet_leaf_66_wb_clk_i net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_3_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10567_ _00461_ clknet_leaf_82_wb_clk_i cpu.last_addr\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_3_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06922__B _02150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10498_ _00393_ clknet_leaf_25_wb_clk_i cpu.timer\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08993__A1 _01133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput6 io_in[14] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_108_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06660_ _02134_ _02135_ _02136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_108_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05611_ cpu.IO_addr_buff\[4\] _01094_ _01038_ _01095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05731__A1 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06591_ _00602_ _00998_ _02067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08330_ _02836_ _03543_ _03545_ _03546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05542_ _01025_ _01026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_74_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08261_ cpu.uart.data_buff\[4\] _03484_ _03489_ _03494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05473_ cpu.regs\[4\]\[4\] cpu.regs\[5\]\[4\] cpu.regs\[6\]\[4\] cpu.regs\[7\]\[4\]
+ _00956_ _00957_ _00960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_22_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07212_ _02658_ _02659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08192_ _03275_ _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_89_Left_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07143_ _00685_ _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_70_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07074_ _00775_ _02537_ _00689_ _02540_ _02541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_06025_ _01075_ _01057_ _01487_ _01506_ _01507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_77_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08736__A1 _02647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07976_ cpu.spi.div_counter\[2\] _03256_ _03250_ _03262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09715_ _04718_ _04673_ _04720_ _04721_ _04722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_98_Left_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_87_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06927_ _02399_ _02400_ _02401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09646_ _04333_ _04648_ _04344_ _04657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_97_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06858_ _00590_ _02334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09577_ _04588_ _04590_ _04591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05809_ _01024_ _01293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06789_ _02242_ _02264_ _02265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08528_ cpu.toggle_top\[5\] _03690_ _03694_ _03686_ _03695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_92_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08459_ cpu.orig_PC\[1\] _03643_ _03646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10074__A3 _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05325__I1 _00831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10421_ _00316_ clknet_leaf_89_wb_clk_i cpu.orig_PC\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10352_ _00247_ clknet_leaf_32_wb_clk_i cpu.uart.div_counter\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05789__A1 _01110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08727__A1 _02631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10283_ _00178_ clknet_leaf_109_wb_clk_i cpu.regs\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05800__I2 cpu.regs\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07799__I _02619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_113_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06208__I _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10619_ _00513_ clknet_leaf_72_wb_clk_i cpu.ROM_spi_cycle\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08966__A1 _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07830_ cpu.timer_div\[6\] _03127_ cpu.timer_div_counter\[7\] _01995_ _03128_ _03129_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__09391__A1 _02093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07761_ _02047_ _03070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09143__A1 cpu.ROM_addr_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09500_ _04329_ _04502_ _04516_ _04366_ _04517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06712_ cpu.regs\[1\]\[6\] _00876_ _02188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07692_ cpu.regs\[5\]\[7\] _03010_ _03020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_69_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09431_ _02766_ _02560_ _04450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06643_ _02097_ _02118_ _02119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05731__B _01113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09362_ _04382_ _04383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06574_ cpu.PC\[6\] _02050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08313_ _03532_ _03533_ _00276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_87_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05525_ _00649_ _01008_ _01009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07502__I _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09293_ _04267_ _04300_ _04316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08244_ _03116_ _03479_ _03480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_105_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05456_ cpu.regs\[4\]\[3\] cpu.regs\[5\]\[3\] cpu.regs\[6\]\[3\] cpu.regs\[7\]\[3\]
+ _00882_ _00884_ _00944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_105_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08175_ _03402_ _03423_ _00248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05387_ _00876_ _00877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_15_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07126_ _00686_ _02589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_45_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07057_ _02523_ _02524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06008_ cpu.uart.divisor\[10\] _01489_ _01490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_7_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09382__A1 _01135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07959_ cpu.spi.data_out_buff\[7\] _03214_ _03247_ _03248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09685__A2 cpu.ROM_addr_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_qcpu_106 io_oeb[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09629_ _00750_ _04636_ _04640_ _04641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06499__A2 _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08508__I _03678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07412__I _02816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_84_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10404_ _00299_ clknet_leaf_17_wb_clk_i cpu.orig_IO_addr_buff\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07287__C _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05306__S0 _00569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10335_ _00230_ clknet_leaf_43_wb_clk_i cpu.uart.dout\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10266_ _00161_ clknet_leaf_118_wb_clk_i cpu.regs\[6\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10197_ _00092_ clknet_leaf_1_wb_clk_i cpu.regs\[14\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05934__A1 _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09676__A2 cpu.ROM_addr_buff\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05310_ cpu.regs\[0\]\[2\] _00817_ _00818_ cpu.regs\[3\]\[2\] _00569_ _00574_ _00819_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06290_ _01357_ _01723_ _01768_ _01769_ _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
Xinput20 io_in[3] net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_116_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput31 sram_out[5] net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__05465__A3 _00952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05241_ _00744_ _00755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_4_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05172_ _00661_ _00665_ _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_40_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07992__I _02516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09980_ _02502_ _04931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06414__A2 _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08931_ cpu.timer_div\[4\] _04000_ _04010_ _04003_ _04011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_0_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08862_ _03166_ _03953_ _03954_ _03959_ _03960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_4_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09364__A1 _02052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07813_ cpu.spi.data_in_buff\[6\] _03101_ _03112_ _03114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08793_ _02703_ _03861_ _03856_ _03901_ _03869_ _03902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_07744_ _02024_ _03051_ _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_79_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07675_ _03009_ _03010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09414_ _04344_ _04434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06626_ _02098_ _02099_ _02102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_109_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06557_ _02032_ cpu.mem_cycle\[4\] _02033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09345_ _04329_ _04332_ _04364_ _04366_ _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_118_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09276_ _02781_ _02765_ _04299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05508_ cpu.regs\[0\]\[5\] cpu.regs\[1\]\[5\] cpu.regs\[2\]\[5\] cpu.regs\[3\]\[5\]
+ net126 _00857_ _00994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06488_ _00613_ _00629_ _01746_ _01965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_7_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08227_ _03464_ _03465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05439_ _00927_ net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_1_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08158_ _03409_ _03410_ _00244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_101_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08089_ _03339_ _03343_ _03347_ _03352_ _03353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__07602__A1 _02556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07109_ _02285_ _02321_ _02573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10120_ _00019_ clknet_leaf_122_wb_clk_i cpu.regs\[9\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10051_ _04952_ _04991_ _04992_ _04993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_101_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07407__I _01788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09107__A1 _03045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09069__I _04125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10318_ _00213_ clknet_leaf_54_wb_clk_i cpu.spi.div_counter\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10249_ _00144_ clknet_leaf_117_wb_clk_i cpu.regs\[8\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05265__C _00778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05790_ _01273_ _01274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_37_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06580__A1 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06377__B _01478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08148__I _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07460_ _00685_ _02870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_17_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06411_ cpu.toggle_top\[14\] _01625_ _01888_ _01889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07391_ _02552_ _02806_ _02807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09130_ _04170_ _04171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06342_ _01764_ _01820_ _01821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09061_ _02505_ _04116_ _04119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08012_ _03289_ _03290_ _00218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_72_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05438__A3 _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06273_ _01634_ _01648_ _01753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05224_ _00686_ _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_71_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05155_ cpu.IO_addr_buff\[2\] _00672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09585__A1 _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09963_ _04918_ _00541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_77_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05086_ _00600_ _00605_ _00583_ _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_65_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_65_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_90_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08914_ _02615_ _03997_ _03998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09894_ net67 _04856_ _04866_ _04862_ _04867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_85_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08845_ _01241_ _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08776_ _03869_ _03888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08560__A2 cpu.toggle_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input12_I io_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05970__I _01452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07727_ _03041_ _00182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05988_ _01302_ _01323_ _01471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08058__I net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07658_ _02983_ _02996_ _02999_ _00155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06609_ _00588_ _00998_ _02085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07589_ _02927_ _02948_ _02956_ _00129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09328_ _04056_ _04350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_80_Left_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09259_ _00721_ _04282_ _04283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_35_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05210__I _00724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06306__I _01784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10103_ _01583_ _05035_ _05039_ _00560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10034_ cpu.startup_cycle\[6\] _02427_ _02423_ _02437_ _04977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__08551__A2 cpu.toggle_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09103__I1 _02570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07114__I0 _02013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07756__B _03065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06960_ _02431_ _02432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input4_I io_in[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05911_ _01368_ _01391_ _01393_ _01184_ _01394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_06891_ _02046_ _02061_ _02366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08542__A2 _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05842_ _01325_ _01326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08630_ _03753_ _03779_ _00347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_55_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08561_ cpu.toggle_ctr\[5\] _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05773_ _01123_ _01257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08492_ _03668_ _03669_ _03667_ _00319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07512_ _02906_ _00102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07443_ cpu.uart.receive_div_counter\[12\] _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_112_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_112_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_91_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09113_ cpu.regs\[3\]\[2\] _03083_ _04150_ _04158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07374_ _02312_ _02309_ _02791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06325_ _01612_ _01803_ _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_79_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09044_ _04102_ _04105_ _00435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06256_ _01636_ _01638_ _01735_ _01736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_103_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05207_ _00648_ _00722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09437__I _04455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06187_ _01650_ _01667_ _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05138_ cpu.base_address\[1\] cpu.base_address\[0\] _00655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_09946_ cpu.PORTB_DDR\[4\] _04903_ _04905_ _04897_ _04906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05069_ _00589_ _00590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09877_ _04037_ _04845_ _04854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_79_Right_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08828_ _03929_ _03894_ _03904_ _03930_ _03898_ _03931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08759_ _03873_ _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_95_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_109_Left_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10652_ _00546_ clknet_leaf_59_wb_clk_i cpu.PORTA_DDR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09097__I0 cpu.regs\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10583_ _00477_ clknet_leaf_94_wb_clk_i cpu.PC\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_88_Right_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09549__A1 _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05875__I _01358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_118_Left_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_97_Right_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10017_ _04147_ _02483_ _04948_ _04961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_47_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05115__I cpu.regs\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07330__I _02698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06110_ cpu.timer_capture\[11\] _01591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_42_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07090_ _02555_ _00031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06041_ _00977_ _01273_ _01277_ _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_74_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09800_ cpu.ROM_spi_dat_out\[2\] _04790_ _04792_ _04793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07992_ _02516_ _03275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06943_ cpu.ROM_spi_cycle\[4\] _02415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09731_ _04733_ _04734_ _04735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_66_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05121__S1 _00631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06774__A1 _00589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09662_ _04671_ _04672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06874_ _02149_ _02331_ _02349_ _02350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09593_ _04056_ _04602_ _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08613_ _03739_ _03767_ _03769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05825_ _01307_ _01308_ _01309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_89_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05756_ _01239_ _01240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_49_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08544_ cpu.toggle_ctr\[12\] _03708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_85_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08475_ _03621_ _03657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05687_ _01024_ _01171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07426_ _02608_ _02837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07357_ _02771_ _02772_ _02775_ _02776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06308_ cpu.spi.dout\[5\] _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_45_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_80_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_80_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07288_ cpu.timer_top\[5\] _02720_ _02722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09027_ _04074_ _04091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06239_ _01414_ _01718_ _01719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09929_ _04891_ _04893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output43_I net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07190__A1 cpu.uart.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08690__A1 _02727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10635_ _00529_ clknet_leaf_67_wb_clk_i net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_36_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10566_ _00460_ clknet_leaf_82_wb_clk_i cpu.last_addr\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05256__A1 _00763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10497_ _00392_ clknet_leaf_24_wb_clk_i cpu.timer\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput7 io_in[15] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06508__A1 cpu.PORTB_DDR\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07181__A1 _02630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05610_ _01074_ _01094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__05731__A2 _01122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10068__A1 _01262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06590_ cpu.regs\[1\]\[6\] _00965_ _02066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05541_ cpu.instr_cycle\[2\] net25 _00659_ _00669_ _01025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_08260_ cpu.uart.data_buff\[3\] _03491_ _03492_ _03493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05472_ _00954_ _00958_ _00851_ _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_116_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08191_ _03323_ _03388_ _03435_ _03398_ _03436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07211_ _01062_ _02658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07142_ _01683_ _02599_ _02601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07073_ _02036_ _02034_ _02539_ _02540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_42_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_35_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06024_ _01488_ _01505_ _01192_ _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09933__A1 _04031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06747__A1 _00900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07975_ _03256_ cpu.spi.div_counter\[0\] _03261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09714_ _04123_ _04721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_87_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06926_ _02384_ _02393_ _02398_ _02400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_97_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09645_ _04121_ _04654_ _04655_ _04656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06857_ _02072_ _02080_ _02333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05808_ _01263_ _01115_ _01292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_2_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09576_ _04387_ _04577_ _04589_ _04439_ _04590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10059__A1 _02593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06788_ _02260_ _02263_ _02264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05739_ cpu.uart.dout\[0\] _01223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08527_ _02750_ _03691_ _03694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08458_ _02783_ _03641_ _03645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_74_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07409_ _02814_ cpu.uart.receive_div_counter\[13\] cpu.uart.receive_div_counter\[6\]
+ _02815_ _02819_ _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_80_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05325__I2 _00832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08389_ _02851_ _03588_ _03593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_98_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10420_ _00315_ clknet_leaf_89_wb_clk_i cpu.orig_PC\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10351_ _00246_ clknet_leaf_33_wb_clk_i cpu.uart.div_counter\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05089__I1 cpu.regs\[9\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10282_ _00177_ clknet_leaf_111_wb_clk_i cpu.regs\[4\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09924__A1 _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07163__A1 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09360__I _04327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08663__A1 _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07710__I0 _03006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10618_ _00512_ clknet_leaf_72_wb_clk_i cpu.ROM_spi_cycle\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10549_ _00443_ clknet_leaf_88_wb_clk_i cpu.ROM_addr_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_11_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09915__A1 net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09535__I _04296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_119_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07760_ _03058_ _03069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06711_ _02185_ _02186_ _02187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09430_ _04421_ _04449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07691_ _03019_ _00168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06642_ _02112_ _02117_ _02118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06901__A1 _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09361_ _04301_ _04382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06573_ cpu.PC\[7\] _02049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08312_ cpu.uart.receive_buff\[4\] _03522_ _03530_ cpu.uart.receive_buff\[5\] _03533_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_86_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05524_ _01006_ _01007_ _01008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xclkbuf_leaf_19_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_19_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09292_ _04307_ _04314_ _00750_ _04315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08243_ _03476_ _03471_ _03478_ _03479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05455_ _00941_ _00942_ _00880_ _00943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_105_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08174_ _03421_ _03418_ _03422_ _03417_ _03423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05386_ _00875_ _00876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_15_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07125_ _01111_ _02586_ _02588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_30_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07056_ _02522_ _02523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09906__A1 _04851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06007_ _01220_ _01489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_100_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07393__A1 _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07958_ _02726_ _03242_ _03247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07889_ cpu.spi.divisor\[1\] _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07145__A1 _02580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06909_ _02368_ _02350_ _02382_ _02384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xwrapped_qcpu_107 io_out[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09628_ _00760_ _04348_ _04639_ _04313_ _04640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_54_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09559_ _04551_ _04573_ _04523_ _00482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_93_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05459__A1 _00880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10403_ _00298_ clknet_leaf_55_wb_clk_i cpu.orig_IO_addr_buff\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09070__A1 _02514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10334_ _00229_ clknet_leaf_43_wb_clk_i cpu.uart.dout\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05306__S1 _00574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10265_ _00160_ clknet_leaf_117_wb_clk_i cpu.regs\[6\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10196_ _00091_ clknet_leaf_2_wb_clk_i cpu.regs\[14\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06928__B _02359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07136__A1 _01135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput10 io_in[18] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput21 io_in[6] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05240_ _00653_ _00656_ _00754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput32 sram_out[6] net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05171_ _00686_ _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09061__A1 _02505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08930_ _02746_ _04009_ _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08861_ _02675_ _03955_ _03959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07812_ _01787_ _03104_ _03113_ _00195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07914__A3 _00756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08792_ cpu.timer\[7\] _03895_ _03901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07743_ _02557_ _03046_ _03049_ _03053_ _03054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__07127__A1 _02580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08875__A1 _02692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07678__A2 _03012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07674_ _01132_ _02977_ _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_48_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09413_ _04057_ _04422_ _04431_ _04432_ _04433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06625_ _00816_ _01955_ _02101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08890__A4 _02729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06556_ _02031_ _02032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09344_ _04365_ _04366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09275_ _04295_ _04298_ _03868_ _00473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05507_ cpu.regs\[4\]\[5\] cpu.regs\[5\]\[5\] cpu.regs\[6\]\[5\] cpu.regs\[7\]\[5\]
+ net126 _00857_ _00993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06487_ _01862_ _01338_ _01942_ _01330_ _01147_ _01964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__08344__I _03517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08226_ _03386_ _03464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05438_ _00715_ _00912_ _00926_ _00927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__05968__I _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08157_ _03333_ _03406_ _03276_ _03410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07108_ _02570_ _02571_ _02572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05369_ _00858_ _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08088_ _03337_ _02818_ _02825_ _03341_ _03351_ _03352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_3_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07602__A2 _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07039_ net19 _02498_ _02508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_10050_ _02432_ _02433_ _04736_ _04974_ _04992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08563__B1 _01410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07366__A1 _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05652__B _01107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06341__A2 _00966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09291__A1 _04309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09594__A2 _04484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10317_ _00212_ clknet_leaf_54_wb_clk_i cpu.spi.div_counter\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10248_ _00143_ clknet_leaf_115_wb_clk_i cpu.regs\[8\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10179_ _00074_ clknet_leaf_116_wb_clk_i _00004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_89_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08857__A1 _02668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06410_ _01885_ _01886_ _01887_ _01123_ _01888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_17_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07380__I1 _02796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07390_ _02055_ _02805_ _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06341_ _01724_ _00966_ _01820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09060_ _04118_ _00438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06272_ _01733_ _01751_ _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__06096__A1 _01315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08011_ cpu.spi.data_in_buff\[0\] _03199_ _03287_ cpu.spi.data_in_buff\[1\] _03290_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05223_ _00728_ _00733_ _00737_ _00738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_72_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05154_ _00648_ _00649_ _00659_ _00670_ _00671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_69_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09962_ cpu.PORTA_DDR\[0\] _04915_ _04917_ _04908_ _04918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_77_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05085_ cpu.regs\[0\]\[5\] _00603_ _00604_ cpu.regs\[3\]\[5\] _00598_ _00599_ _00605_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_90_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08913_ _03995_ _03997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09893_ _04052_ _04857_ _04866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08844_ _03942_ _03944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08775_ cpu.timer\[4\] _03836_ _03858_ _03886_ _03881_ _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05987_ _01468_ _01469_ _01470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_34_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_34_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07726_ _03002_ cpu.regs\[3\]\[4\] _03034_ _03041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08848__A1 _02707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07520__A1 _01109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07657_ cpu.regs\[6\]\[1\] _02997_ _02999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06608_ _00601_ _00964_ _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07588_ cpu.regs\[10\]\[7\] _02946_ _02956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09327_ _04348_ _04349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06539_ cpu.regs\[9\]\[7\] _01681_ _02016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09258_ _00748_ _04269_ _04281_ _04282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08209_ cpu.uart.clr_hb _03450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09189_ _04212_ _04215_ _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output73_I net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10102_ cpu.regs\[15\]\[2\] _05036_ _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06322__I _01183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10033_ _04732_ _02423_ _02437_ _04975_ _04976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07354__A4 _02583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05382__B _00871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08839__A1 _03176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07578__A1 cpu.regs\[10\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05910_ _01392_ _01368_ _01393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06890_ _01857_ _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05841_ _00970_ _00930_ _00655_ _01325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__06002__A1 _01153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08560_ _03723_ cpu.toggle_top\[6\] _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05772_ cpu.toggle_top\[8\] _01256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_08491_ cpu.orig_PC\[10\] _03659_ _03669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07511_ _01772_ cpu.regs\[13\]\[4\] _02899_ _02906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07442_ _02841_ _02849_ _02852_ _02853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_71_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07373_ _02789_ _02782_ _02790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06324_ cpu.timer_div\[5\] _01801_ _01803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09112_ _04157_ _00451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09043_ cpu.IO_addr_buff\[5\] _04097_ _04104_ _04100_ _04105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_60_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06255_ _01635_ _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_115_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_111_Right_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05206_ _00719_ _00720_ _00721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_13_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06186_ _01569_ _01666_ _01667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05137_ cpu.base_address\[3\] cpu.base_address\[2\] _00654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_111_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09945_ _04041_ _04904_ _04905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05068_ _00588_ _00589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09876_ _04853_ _00519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08827_ _03929_ _03924_ _03930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07741__A1 _02024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08758_ cpu.timer_capture\[1\] _03870_ _03872_ _03820_ _03873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08689_ _02620_ _03822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07709_ _03030_ _00175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10651_ _00545_ clknet_leaf_59_wb_clk_i cpu.PORTA_DDR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09097__I1 _02559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10582_ _00476_ clknet_leaf_94_wb_clk_i cpu.PC\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10016_ _04956_ _04945_ _04960_ _03366_ _00552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05891__I _01210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09088__I1 cpu.ROM_addr_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09237__A1 cpu.Z vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_25_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06040_ _01175_ _01519_ _01521_ _01261_ _00909_ _01522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_TAPCELL_ROW_74_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07991_ _03272_ _03252_ _03273_ _03259_ _03274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09730_ cpu.startup_cycle\[0\] _04734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06774__A2 _00906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06942_ _02414_ _00024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09273__I _04296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05734__C _01088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09661_ _02492_ _04020_ _00732_ _04671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06873_ _02345_ _02348_ _02349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07723__A1 _01583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09592_ _04387_ _04603_ _04604_ _04390_ _04605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08612_ _03756_ _03767_ _03768_ _00340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05824_ _00874_ net121 _01308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05755_ _01238_ _01239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09476__A1 _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08543_ _03702_ _03705_ _03706_ _03707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_85_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10086__A2 _05024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08474_ _03655_ _03656_ _03650_ _00314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05686_ _01169_ _01170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_9_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_64_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07425_ cpu.uart.receive_div_counter\[1\] _02836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_64_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07356_ _02774_ _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_73_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07287_ _02635_ _02719_ _02721_ _02716_ _00062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06307_ cpu.timer_top\[5\] _01786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_32_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08451__A2 _03636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09026_ _04084_ _04090_ _00432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06238_ _01174_ _01715_ _01716_ _01717_ _00950_ _01718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_33_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06169_ _01637_ _01650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06214__A1 net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09928_ _04891_ _04892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09859_ _00733_ _00737_ net89 _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_96_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output36_I net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09219__A1 _01135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10634_ _00528_ clknet_leaf_67_wb_clk_i net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_102_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06047__I _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10565_ _00459_ clknet_leaf_82_wb_clk_i cpu.last_addr\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09358__I _04296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05256__A2 _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10496_ _00391_ clknet_leaf_24_wb_clk_i cpu.timer\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_109_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07953__A1 _02646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06300__S1 _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08211__B _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput8 io_in[16] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06508__A2 _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_108_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05540_ _01023_ _01024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08130__A1 _03364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05471_ cpu.regs\[8\]\[4\] cpu.regs\[9\]\[4\] cpu.regs\[10\]\[4\] cpu.regs\[11\]\[4\]
+ _00956_ _00957_ _00958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_08190_ _03323_ _03434_ _03435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07210_ cpu.timer\[0\] _02657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_55_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07141_ _02599_ _02600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07072_ _02463_ _02538_ _02539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_70_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06444__B2 _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06023_ _01490_ _01504_ _01194_ _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07974_ _03257_ _03260_ _02871_ _00210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09713_ _04672_ _04710_ _04719_ _04720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_87_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06925_ net118 _02393_ _02398_ _02399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07960__B _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09644_ _00932_ _04654_ _04455_ _04655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06856_ _02083_ _02096_ _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05807_ _01290_ _01291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__05183__A1 cpu.TIE vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09575_ cpu.orig_PC\[10\] _04437_ _04589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06787_ _02261_ _02262_ _02263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05738_ _01196_ _01219_ _01221_ _01222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08526_ _03693_ _00329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08457_ _03642_ _03644_ _03633_ _00309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05669_ _01152_ _01153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07408_ _02816_ _02817_ cpu.uart.receive_div_counter\[5\] _02818_ _02819_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_65_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05325__I3 cpu.regs\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08388_ _02851_ _03588_ _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_98_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07339_ _02761_ _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_45_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10350_ _00245_ clknet_leaf_33_wb_clk_i cpu.uart.div_counter\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06435__A1 _01326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09009_ _04063_ _04076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10281_ _00176_ clknet_leaf_116_wb_clk_i cpu.regs\[4\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07426__I _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_57_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08112__A1 _03366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07161__I _02612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09860__A1 _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06674__A1 cpu.regs\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10617_ _00511_ clknet_leaf_72_wb_clk_i cpu.ROM_spi_cycle\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08415__A2 _03611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09612__A1 _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10548_ _00442_ clknet_leaf_88_wb_clk_i cpu.ROM_addr_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_51_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10479_ _00374_ clknet_leaf_19_wb_clk_i cpu.timer_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07926__A1 _00904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08720__I _02723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06710_ _02137_ _02146_ _02186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_63_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07690_ _03006_ cpu.regs\[5\]\[6\] _03009_ _03019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_69_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06641_ _02115_ _02116_ _02117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09360_ _04327_ _04381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06572_ cpu.PC\[8\] _02048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08311_ _03401_ _03532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_82_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05523_ _00648_ cpu.instr_cycle\[3\] cpu.instr_cycle\[1\] _00670_ _01007_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_09291_ _04309_ _04300_ _04312_ _04313_ _04314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_47_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08242_ cpu.uart.data_buff\[0\] _03453_ _03477_ _03478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_74_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05454_ cpu.regs\[8\]\[3\] cpu.regs\[9\]\[3\] cpu.regs\[10\]\[3\] cpu.regs\[11\]\[3\]
+ _00888_ _00889_ _00942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xclkbuf_leaf_59_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_59_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_74_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07862__B1 cpu.timer\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08173_ _03421_ _03392_ _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05385_ _00862_ _00868_ _00872_ _00874_ _00875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__07020__B _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07124_ _02586_ _02587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07055_ _01528_ _01011_ _01143_ _02522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_112_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06006_ cpu.uart.dout\[2\] _00012_ _01488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05640__A2 _01122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_93_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07957_ _03235_ _03244_ _03246_ _00207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07246__I _02639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08786__B _02697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06908_ _02368_ _02350_ _02382_ _02383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07888_ _03181_ cpu.spi.divisor\[2\] _03182_ cpu.spi.div_counter\[7\] _03185_ _03186_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_69_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09627_ _04303_ _04638_ _04639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_54_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06839_ _02306_ _02311_ _02315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xwrapped_qcpu_108 io_out[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09558_ _04328_ _04569_ _04572_ _04573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08509_ _02615_ _03680_ _03681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09489_ _04504_ _04505_ _04455_ _04506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_38_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Left_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10402_ _00297_ clknet_leaf_55_wb_clk_i cpu.orig_IO_addr_buff\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10333_ _00228_ clknet_leaf_44_wb_clk_i cpu.uart.dout\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05631__A2 _00717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10264_ _00159_ clknet_leaf_114_wb_clk_i cpu.regs\[6\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10195_ _00090_ clknet_leaf_3_wb_clk_i cpu.regs\[14\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07156__I _02610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_21_Left_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09371__I _04273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07136__A2 _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09833__A1 _03207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput11 io_in[19] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput22 io_in[7] net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput33 sram_out[7] net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05170_ _00685_ _00686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_12_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05870__A2 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05622__A2 _01065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08860_ _03958_ _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07811_ cpu.spi.data_in_buff\[5\] _03107_ _03112_ _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_4_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08791_ _03899_ _03900_ _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07742_ _03052_ _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05138__A1 cpu.base_address\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07673_ _02992_ _02997_ _03008_ _00161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09412_ _04303_ _04432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06624_ _02098_ _02099_ _02100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06886__A1 _02359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09124__I0 cpu.regs\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09343_ _02511_ _00757_ _04365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07730__S _03033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06555_ cpu.mem_cycle\[5\] _02031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09274_ _02768_ _04297_ _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05506_ _00990_ _00991_ _00850_ _00992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06486_ net97 _01962_ _01963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08225_ _03456_ _03362_ _03463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05437_ _00925_ _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_15_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_95_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08156_ _03333_ _03405_ _03407_ _03408_ _03409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05368_ _00857_ _00858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_16_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07107_ _02558_ _02560_ _02571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08087_ _03349_ _02622_ _02837_ _03350_ _03351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_05299_ cpu.regs\[12\]\[1\] cpu.regs\[13\]\[1\] cpu.regs\[14\]\[1\] cpu.regs\[15\]\[1\]
+ _00568_ _00573_ _00809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07038_ _02507_ _00027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08989_ _04055_ _04056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09191__I _04213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06326__B1 _01802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05652__C _00970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05224__I _00686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08079__B1 _02630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09366__I _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_4_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_4_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10316_ _00211_ clknet_leaf_57_wb_clk_i cpu.spi.div_counter\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10247_ _00142_ clknet_leaf_125_wb_clk_i cpu.regs\[8\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10178_ _00011_ clknet_leaf_89_wb_clk_i cpu.instr_cycle\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10113__A1 _02014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09282__A2 _00762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06340_ _01818_ _01819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07293__A1 _02647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06271_ _01734_ _01737_ _01740_ _01750_ _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08010_ _02873_ _03289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05222_ _00734_ _00735_ _00736_ _00730_ _00699_ _00737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_60_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05153_ _00669_ _00670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08180__I _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09961_ _02707_ _04916_ _04917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_77_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08793__A1 _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05084_ cpu.regs\[2\]\[5\] _00604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_90_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08912_ _03995_ _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09892_ _04865_ _00523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08843_ _03942_ _03943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08774_ _03884_ _03885_ _03886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05986_ _01465_ _01466_ _01430_ _01469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07725_ _01679_ _03035_ _03040_ _00181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06859__A1 _02334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07656_ _02975_ _02996_ _02998_ _00154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_74_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_74_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_48_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06607_ _02081_ _02082_ _02083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07587_ _02955_ _00128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09326_ _04277_ _04348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06538_ _02014_ _02015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09257_ _04270_ _04275_ _04280_ _00747_ _04281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_7_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08208_ _03427_ _03449_ _00255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06469_ _01899_ _01903_ _01898_ _01946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09188_ _04078_ _04214_ _00723_ _04215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08139_ _03348_ _03345_ _03395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10101_ _01481_ _05035_ _05038_ _00559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output66_I net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10032_ _04748_ _04974_ _04975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_4_4_0_wb_clk_i clknet_0_wb_clk_i clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05889__I _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07275__A1 _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_15_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_113_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05589__A1 _01070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08527__A1 _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06389__I0 cpu.PORTA_DDR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05840_ _01319_ _01322_ _01323_ _01324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05771_ _01176_ _01178_ _01250_ _01253_ _01254_ _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_07510_ _01680_ _02900_ _02905_ _00101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08490_ _03083_ _03657_ _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07441_ _02847_ _02850_ _02851_ cpu.uart.divisor\[13\] _02852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_clkbuf_leaf_54_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07372_ _02788_ _02789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06323_ _01787_ _01187_ _01799_ _01800_ _01801_ _01802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__07266__A1 cpu.timer_capture\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09111_ _04156_ cpu.ROM_addr_buff\[9\] _04148_ _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09042_ _00740_ _04069_ _04071_ _04103_ _04094_ _04104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_5_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06254_ _01441_ _01734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05205_ cpu.uart.busy cpu.spi.busy _00720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06185_ _01531_ _00936_ _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05136_ cpu.instr_buff\[15\] _00651_ cpu.base_address\[5\] _00652_ _00653_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xclkbuf_leaf_121_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_121_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_13_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07519__I _01359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09944_ _04891_ _04904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05067_ cpu.regs\[1\]\[4\] _00588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09875_ net61 _04844_ _04852_ _04849_ _04853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08826_ cpu.timer\[13\] _03929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_93_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07741__A2 _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08757_ _03176_ _03871_ _03860_ _03872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05969_ _01298_ _00848_ _01320_ _01452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_95_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08688_ _03821_ _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07708_ _03004_ cpu.regs\[4\]\[5\] _03021_ _03030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07639_ _01678_ _02987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10650_ _00544_ clknet_leaf_60_wb_clk_i cpu.PORTA_DDR\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09309_ _02788_ _04330_ _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_36_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10581_ _00475_ clknet_leaf_105_wb_clk_i cpu.PC\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08034__B _02871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08757__A1 _03176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08509__A1 _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10015_ _02435_ _04959_ _04945_ _04960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05743__A1 cpu.uart.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_4_Left_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05412__I _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08748__A1 _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05106__S0 _00615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07990_ _03272_ _03268_ _03273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06941_ cpu.regs\[2\]\[7\] _02413_ _02363_ _02414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09660_ _02442_ _04670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08611_ cpu.toggle_ctr\[7\] _03766_ _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06872_ _02346_ _02118_ _02347_ _02348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__05734__A1 _01214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09591_ cpu.orig_PC\[11\] _04437_ _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05823_ net122 _00868_ _01307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05754_ _01046_ _01096_ _01238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08542_ cpu.toggle_ctr\[11\] _01624_ _01520_ _03703_ _03706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_85_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08473_ cpu.orig_PC\[5\] _03643_ _03656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07424_ cpu.uart.receive_div_counter\[5\] _02835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_77_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_59_Left_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05685_ _01168_ _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_92_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05322__I _00829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07239__A1 cpu.timer_capture\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07355_ _02523_ _02535_ _02520_ _02773_ _02774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_116_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07286_ cpu.timer_top\[4\] _02720_ _02721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08633__I _03551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06306_ _01784_ _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_33_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09025_ _00673_ _04067_ _04089_ _04082_ _04090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06237_ _01260_ _01717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07249__I cpu.timer\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06168_ _01634_ _01648_ _01649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_40_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06214__A2 _01210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Left_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05119_ cpu.regs\[12\]\[7\] cpu.regs\[13\]\[7\] cpu.regs\[14\]\[7\] cpu.regs\[15\]\[7\]
+ _00630_ _00631_ _00637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06099_ net28 _01579_ _01580_ _01581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09927_ _01101_ _04842_ _04891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08911__A1 _01054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09858_ _04823_ _04837_ _04838_ _04839_ _03288_ _00515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_09789_ _04783_ _00502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08809_ _03912_ _03915_ _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_68_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_77_Left_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09467__A2 _04484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06150__A1 cpu.TIE vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09219__A2 _02271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10633_ _00527_ clknet_leaf_65_wb_clk_i net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_52_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10564_ _00458_ clknet_leaf_77_wb_clk_i cpu.last_addr\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10495_ _00390_ clknet_leaf_25_wb_clk_i cpu.timer\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07159__I _01419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07402__A1 _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09155__A1 cpu.ROM_addr_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput9 io_in[17] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08718__I _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09458__A2 _00701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08130__A2 _03386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05470_ _00005_ _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_55_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07140_ _02598_ _02599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05327__S0 _00570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07071_ _02027_ _02030_ _02538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06022_ _01491_ _01503_ _01196_ _01504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09394__A1 _02513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09712_ _04718_ _02539_ _04719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07973_ _03258_ _03250_ _03259_ _03260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05955__A1 _00844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06924_ _02395_ _02397_ _02398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_87_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09643_ cpu.PC\[13\] _04653_ _04654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06855_ _02187_ _02329_ _02330_ _02331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09574_ _00751_ _04584_ _04587_ _04588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05806_ _01289_ _01290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08525_ cpu.toggle_top\[4\] _03690_ _03692_ _03686_ _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06786_ _02258_ _02259_ _02262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05737_ cpu.uart.divisor\[8\] _01220_ _01221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06132__A1 cpu.timer_div\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08456_ cpu.orig_PC\[0\] _03643_ _03644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05668_ _01151_ _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_37_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08387_ _03580_ _03591_ _00292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07407_ _01788_ _02818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_80_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05599_ _01037_ _01082_ _01083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07338_ _00768_ _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_98_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07269_ _02707_ _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_60_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09008_ _04074_ _04075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10280_ _00175_ clknet_leaf_100_wb_clk_i cpu.regs\[4\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09688__A2 cpu.ROM_addr_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_85_Left_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_57_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06674__A2 _01286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10616_ _00510_ clknet_leaf_71_wb_clk_i cpu.ROM_spi_cycle\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_94_Left_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09612__A2 _04499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10547_ _00441_ clknet_leaf_96_wb_clk_i cpu.base_address\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_118_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10478_ _00373_ clknet_leaf_18_wb_clk_i cpu.timer_top\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_71_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05937__A1 _01419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06640_ _02109_ _02111_ _02116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06362__A1 _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05796__S0 _00864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06571_ cpu.PC\[10\] _02047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08310_ _03519_ _03531_ _00275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05522_ _00648_ _01006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09290_ _04270_ _04313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08241_ _03470_ _03477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05801__S _00852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05453_ cpu.regs\[12\]\[3\] cpu.regs\[13\]\[3\] cpu.regs\[14\]\[3\] cpu.regs\[15\]\[3\]
+ _00888_ _00889_ _00941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_103_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08172_ cpu.uart.div_counter\[8\] _03421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05384_ _00873_ _00853_ _00874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_70_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07614__A1 cpu.regs\[8\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07123_ _02585_ _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05476__I0 _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07728__S _03033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07054_ _02520_ _02521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_88_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_28_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_28_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06005_ cpu.spi.busy _01079_ _01487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_2_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05640__A3 _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05928__A1 _01410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07956_ cpu.spi.data_out_buff\[5\] _03218_ _03245_ _03246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input28_I sram_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06907_ _02378_ _02381_ _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_106_Right_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07887_ _03184_ cpu.spi.divisor\[3\] _03182_ cpu.spi.div_counter\[7\] _03185_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09626_ _04623_ _00763_ _04637_ _04638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_54_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06838_ _02307_ _02313_ _02314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xwrapped_qcpu_109 io_out[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09557_ _04443_ _04555_ _04571_ _04547_ _04375_ _04572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_06769_ _00588_ _00876_ _02245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08508_ _03678_ _03680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09488_ _02569_ _02606_ _04505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_38_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08439_ cpu.orig_IO_addr_buff\[7\] _03627_ _03632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10401_ _00296_ clknet_leaf_57_wb_clk_i cpu.needs_interrupt vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10332_ _00227_ clknet_leaf_47_wb_clk_i cpu.uart.dout\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output96_I net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05092__A1 _00567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10263_ _00158_ clknet_leaf_118_wb_clk_i cpu.regs\[6\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10194_ _00089_ clknet_leaf_45_wb_clk_i cpu.uart.receive_counter\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09530__A1 _00790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_32_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09099__I _04022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput12 io_in[1] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_83_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05420__I _00908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput23 io_in[8] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08731__I _02723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05458__I0 cpu.regs\[0\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07810_ _03111_ _03112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08790_ cpu.timer_capture\[6\] _03888_ _03889_ _03900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08572__A2 cpu.toggle_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07741_ _02024_ _03051_ _03052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08324__A2 _03518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05138__A2 cpu.base_address\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07672_ cpu.regs\[6\]\[7\] _02995_ _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09411_ _04418_ _04068_ _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06623_ _00829_ _00997_ _02099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06886__A2 _02361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08088__A1 _03337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06554_ _02029_ _02030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09124__I1 _03674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09342_ _04346_ _04357_ _04363_ _04364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05505_ cpu.regs\[8\]\[5\] cpu.regs\[9\]\[5\] cpu.regs\[10\]\[5\] cpu.regs\[11\]\[5\]
+ net125 _00857_ _00991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_118_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09273_ _04296_ _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06638__A2 _02064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06485_ net95 net96 _01757_ _01962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_16_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08224_ _03462_ _00258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_117_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05436_ _00924_ _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_117_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08155_ _03383_ _03408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_95_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05367_ _00005_ _00857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_16_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07106_ _02569_ _02570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08086_ cpu.uart.div_counter\[0\] _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05298_ _00803_ _00807_ _00579_ _00808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_100_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07257__I _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07037_ _00764_ _02496_ _02506_ _02503_ _02507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08988_ _01140_ _04055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07939_ _03231_ _03225_ _03232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06326__A1 cpu.timer_capture\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09609_ _04575_ _04618_ _04619_ _04621_ _04081_ _04622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_97_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08079__B2 _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08037__B _02871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10315_ _00210_ clknet_leaf_57_wb_clk_i cpu.spi.div_counter\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07167__I _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10246_ _00141_ clknet_leaf_126_wb_clk_i cpu.regs\[8\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10177_ _00010_ clknet_leaf_58_wb_clk_i cpu.instr_cycle\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06565__A1 _02024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06317__A1 _01788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_44_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07630__I _02978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08490__A1 _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06270_ _01440_ _01743_ _01749_ _01548_ _01750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05221_ _00696_ _00722_ _00736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05152_ net71 _00661_ _00665_ _00668_ _00669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__09990__A1 _03822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09960_ _04914_ _04916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_77_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05083_ _00602_ _00603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08911_ _01054_ _01077_ _01234_ _02611_ _03995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_40_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09891_ net66 _04856_ _04864_ _04862_ _04865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_85_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08842_ _01055_ _01234_ _02611_ _03942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA_clkbuf_leaf_83_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08773_ cpu.timer\[3\] _03875_ cpu.timer\[4\] _03885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05985_ _00845_ _01001_ _01141_ _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_07724_ cpu.regs\[3\]\[3\] _03034_ _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07655_ cpu.regs\[6\]\[0\] _02997_ _02998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06606_ _00590_ _01288_ _02082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_40_Left_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_75_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07586_ _02942_ cpu.regs\[10\]\[6\] _02945_ _02955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09325_ _00750_ _04347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06537_ _02013_ _02014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_62_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09256_ _01163_ _04277_ _04279_ _04270_ _04280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_8_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06468_ _01944_ _01945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_43_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_43_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08207_ cpu.uart.div_counter\[15\] _03445_ _03448_ _03449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05419_ _00907_ _00908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06399_ cpu.uart.dout\[6\] _01369_ _01874_ _01876_ _01080_ _01877_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_09187_ _04073_ _04213_ _04214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08233__A1 _03364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08138_ _03350_ _03392_ _03393_ _03394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07036__A2 _02505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08069_ cpu.uart.div_counter\[4\] _03333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_101_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10100_ cpu.regs\[15\]\[1\] _05036_ _05038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10031_ _02421_ _04755_ _02436_ _04974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__07715__I _03033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output59_I net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06011__A3 _01046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05770__A2 _01202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08472__A1 _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06066__I _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09724__A1 _04169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06389__I1 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10229_ _00124_ clknet_leaf_0_wb_clk_i cpu.regs\[10\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05770_ _01096_ _01202_ _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_55_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_0_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07440_ cpu.uart.receive_div_counter\[13\] _02851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_9_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07360__I _02270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07371_ _02053_ _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06322_ _01183_ _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09110_ cpu.regs\[3\]\[1\] _03664_ _04150_ _04156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09041_ cpu.orig_IO_addr_buff\[5\] _04091_ _04092_ _00999_ _04103_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_115_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06253_ _01726_ _01732_ _01733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05204_ _00704_ _00718_ _00658_ _00719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_4_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06184_ _01654_ _01659_ _01664_ _01665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05135_ cpu.base_address\[4\] _00652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_96_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09943_ _04891_ _04903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05066_ _00586_ _00587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09874_ _04851_ _04845_ _04852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08825_ _03927_ _03928_ _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input10_I io_in[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08756_ cpu.timer\[1\] _03862_ _03871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08794__C _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05055__I _00575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05968_ _01450_ _01451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05899_ net7 _01372_ _01379_ _01381_ _01382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_95_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08687_ cpu.pwm_top\[6\] _03814_ _03819_ _03820_ _03821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07707_ _03029_ _00174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07638_ _02985_ _02980_ _02986_ _00148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07569_ _02927_ _02933_ _02944_ _00121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09308_ _02781_ _02766_ _04330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05268__A1 _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08454__A1 _02768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10580_ _00474_ clknet_leaf_90_wb_clk_i cpu.PC\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09239_ _04059_ _04238_ _04257_ _04263_ _04264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_8_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07646__S _02978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10014_ _04957_ _04958_ _04953_ _04959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_116_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05743__A2 _01079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06940__A1 _02013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_63_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09945__A1 _04041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_75_Right_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_105_Left_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06940_ _02013_ _02407_ _02411_ _02412_ _02413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input2_I io_in[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06871_ _02065_ _02119_ _02347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05982__A2 _01340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08610_ _03721_ _03722_ _03762_ _03767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_05822_ _01299_ _01300_ _01306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_89_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_84_Right_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09590_ _04602_ _04603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05753_ _01182_ _01231_ _01233_ _01236_ _01237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_08541_ _03703_ _01520_ _03701_ _03704_ _03705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_106_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08472_ _02550_ _03641_ _03655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05684_ cpu.C _01168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07423_ _02828_ _02829_ _02830_ _02831_ _02833_ _02834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XPHY_EDGE_ROW_114_Left_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07354_ _00775_ _02537_ _00689_ _02583_ _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_72_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07285_ _02710_ _02720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06305_ _01783_ _01784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08135__B _03364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_93_Right_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09024_ _01153_ _04070_ _04072_ _04088_ _04079_ _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_06236_ cpu.toggle_top\[12\] _01625_ _01716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_103_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05670__A1 _01153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07974__B _02871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06167_ _01426_ _01639_ _01647_ _01648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05118_ _00632_ _00635_ _00621_ _00636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06098_ _01424_ _01580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09926_ _04890_ _00532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05049_ _00569_ _00570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07175__A1 _02627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09857_ _03784_ _03782_ cpu.pwm_counter\[3\] _03786_ _04839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_09788_ cpu.ROM_spi_dat_out\[1\] _04778_ _04782_ _04721_ _04783_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08808_ cpu.timer_capture\[9\] _03913_ _03914_ _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08739_ _03130_ _03855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09413__C _04432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08675__A1 _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10632_ _00526_ clknet_leaf_65_wb_clk_i net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10563_ _00457_ clknet_leaf_77_wb_clk_i cpu.last_addr\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09927__A1 _01101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10494_ _00389_ clknet_leaf_25_wb_clk_i cpu.timer\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07650__A2 _02981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05661__A1 _01010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06213__I0 cpu.PORTA_DDR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10481__CLK clknet_leaf_18_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07903__I _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08666__A1 _02735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06677__B1 _01286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09091__A1 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07070_ _02536_ _02537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_42_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06254__I _01441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05327__S1 _00827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06021_ _01500_ _01501_ _01502_ _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05652__A1 _01135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07641__A2 _02980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05404__A1 _00880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09711_ _02035_ _04718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07972_ _03202_ _03259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06923_ _02150_ _02340_ _02396_ _02397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_87_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09642_ _04651_ _04633_ _04652_ _04653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06854_ _02120_ _02148_ _02330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09573_ _04121_ _04349_ _04586_ _04344_ _04587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05805_ _01288_ _01289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06785_ _02252_ _02254_ _02249_ _02261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05736_ _01195_ _01220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_77_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08524_ _02746_ _03691_ _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05333__I _00840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08455_ _03626_ _03643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05667_ cpu.br_rel_dest\[2\] _01151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08386_ cpu.uart.receive_div_counter\[12\] _03557_ _03588_ _03590_ _03591_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07406_ cpu.uart.receive_div_counter\[9\] _02817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05598_ _01039_ _01038_ _01082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07337_ _02586_ _02760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_98_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07268_ _02614_ _02707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_5_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07632__A2 _02980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09909__A1 _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06219_ net10 _01204_ _01200_ _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07199_ _02647_ _02636_ _02648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09007_ _04073_ _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09909_ _04037_ _04870_ _04878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07148__A1 _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08896__A1 _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output41_I net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05243__I _00756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08982__C _04050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10615_ _00509_ clknet_leaf_71_wb_clk_i cpu.ROM_spi_cycle\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_3_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10546_ _00440_ clknet_leaf_96_wb_clk_i cpu.base_address\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_3_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10477_ _00372_ clknet_leaf_29_wb_clk_i cpu.timer_div_counter\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_118_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05418__I _00906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08729__I _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07633__I _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05796__S1 _00865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05153__I _00669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06570_ cpu.PC\[12\] _02046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05521_ _01005_ net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07311__A1 _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08240_ cpu.uart.data_buff\[1\] _03476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05452_ _00896_ _00940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08171_ _03402_ _03420_ _00247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07862__A2 cpu.timer\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07122_ _02536_ _02583_ _02584_ _02493_ _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_70_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05383_ cpu.regs\[8\]\[0\] cpu.regs\[9\]\[0\] cpu.regs\[10\]\[0\] cpu.regs\[11\]\[0\]
+ _00856_ _00860_ _00873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_70_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07053_ _01132_ _02020_ _02520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05625__A1 _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06004_ cpu.timer_capture\[10\] _01486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_11_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07378__A1 _01582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_68_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_68_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07955_ _03111_ _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08878__A1 cpu.timer_capture\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06906_ _02379_ _02380_ _02381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07886_ _03183_ _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09625_ _00762_ _04625_ _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07543__I _02014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06837_ _02299_ _02312_ _02309_ _02313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_09556_ _00806_ _04369_ _04570_ _04571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06768_ _00816_ _00933_ _02244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05719_ _01027_ _01030_ _01202_ _01203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_09487_ _04477_ _04478_ _04503_ _04504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08507_ _03678_ _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06699_ _02170_ _02174_ _02175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08438_ cpu.IO_addr_buff\[7\] _03622_ _03631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05998__I _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05864__A1 _00971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08369_ _02830_ _03571_ _03577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_46_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10400_ _00295_ clknet_leaf_38_wb_clk_i cpu.uart.receive_div_counter\[15\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10331_ _00226_ clknet_leaf_45_wb_clk_i cpu.uart.dout\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05616__A1 _01010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output89_I net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10262_ _00157_ clknet_leaf_111_wb_clk_i cpu.regs\[6\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05631__A4 _01071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10193_ _00088_ clknet_leaf_47_wb_clk_i cpu.uart.receive_counter\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06041__A1 _00977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_34_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput13 io_in[20] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09046__A1 _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput24 io_in[9] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09597__A2 _00930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10529_ _00423_ clknet_leaf_40_wb_clk_i cpu.uart.divisor\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_12_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05458__I1 _00829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07628__I _02978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06280__A1 _01757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_73_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07791__C _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06032__A1 _01486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07740_ _02536_ _03050_ _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06583__A2 _02058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07671_ _03007_ _00160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07532__A1 cpu.regs\[12\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09410_ _04348_ _04430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06622_ _00588_ _00964_ _02098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06553_ _02028_ _02029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09341_ _04358_ _04332_ _04360_ _04362_ _04363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_59_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09285__A1 _00970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05504_ cpu.regs\[12\]\[5\] cpu.regs\[13\]\[5\] cpu.regs\[14\]\[5\] cpu.regs\[15\]\[5\]
+ _00956_ _00957_ _00990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_09272_ _01007_ _04296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_115_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_115_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06484_ _01655_ _01960_ _01961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08223_ cpu.uart.counter\[1\] _03458_ _03460_ _03461_ _03462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_90_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05435_ _00923_ _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_08154_ _03333_ _03406_ _03407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05366_ _00855_ _00856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_113_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08085_ _03348_ _03349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_70_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07105_ _02049_ _02569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07036_ _02497_ _02505_ _02506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06271__A1 _01734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05297_ cpu.regs\[0\]\[1\] _00805_ _00806_ cpu.regs\[3\]\[1\] _00801_ _00802_ _00807_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_101_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08548__B1 cpu.toggle_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08987_ _04054_ _00429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07771__A1 _00818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07938_ _00951_ _03231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07869_ cpu.timer_top\[10\] _03166_ _03167_ cpu.timer_top\[9\] _03168_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09608_ _04291_ _04603_ _04620_ _04547_ _04621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_104_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09539_ _03060_ _04552_ _04553_ _04554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_39_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06617__I _00831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_118_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09928__I _04891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10314_ _00209_ clknet_leaf_62_wb_clk_i cpu.spi.div_counter\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09200__A1 _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10245_ _00140_ clknet_leaf_127_wb_clk_i cpu.regs\[8\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10176_ _00009_ clknet_leaf_89_wb_clk_i cpu.instr_cycle\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07183__I _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09019__B2 _02668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05220_ cpu.instr_buff\[14\] _00735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05151_ _00666_ _00667_ _00668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_52_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08242__A2 _03453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05082_ _00601_ _00602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09890_ _04048_ _04857_ _04864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_90_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08910_ _02727_ _03989_ _03994_ _00412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06005__A1 cpu.spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08841_ _03941_ _00396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_85_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08772_ _02685_ _02679_ _03879_ _03884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_05984_ _01465_ _01466_ _01443_ _01467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07723_ _01583_ _03035_ _03039_ _00180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08917__I _03995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07654_ _02994_ _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06605_ _02072_ _02080_ _02081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_94_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09241__C _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07585_ _02954_ _00127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09324_ _04334_ _04331_ _04343_ _04345_ _04346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_8_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06536_ _01479_ _01977_ _02012_ _02013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_106_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09255_ _04276_ _04278_ _04279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06467_ _01942_ _01943_ _01944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05819__A1 _01111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08206_ cpu.uart.div_counter\[15\] _03391_ _03443_ _03448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08481__A2 _03659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06492__B2 _01321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05418_ _00906_ _00907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06398_ _01224_ _01875_ _01876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09186_ _04019_ _04062_ _04213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08233__A2 _03358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05349_ cpu.PORTB_DDR\[1\] net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_08137_ _03387_ _03393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07268__I _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08068_ cpu.uart.divisor\[11\] cpu.uart.div_counter\[11\] _03332_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_101_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_83_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_83_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_31_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07019_ _02477_ _02480_ _02490_ _02491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_12_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_12_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_12_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10030_ _04709_ _04972_ _04939_ _04973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09483__I _04499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06900__I _00634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07744__A1 _02024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09249__A1 _00928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07178__I cpu.uart.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06235__A1 cpu.toggle_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09393__I _04226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10228_ _00123_ clknet_leaf_0_wb_clk_i cpu.regs\[10\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07735__A1 _03045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10159_ _00058_ clknet_leaf_18_wb_clk_i cpu.timer_top\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08160__A1 _03337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06458__S _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07370_ _02787_ _00079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06321_ cpu.spi.divisor\[5\] _01606_ _01190_ _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_17_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09040_ _02870_ _04102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06252_ _01331_ _01727_ _01731_ _01451_ _01732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_72_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05203_ _00711_ _00717_ _00718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__08215__A2 _03453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06183_ _01144_ _01639_ _01663_ _01548_ _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07423__B1 _02830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05134_ cpu.instr_buff\[14\] _00651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_111_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09942_ _04902_ _00536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_96_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05065_ _00002_ _00586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09873_ _00925_ _04851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08824_ cpu.timer_capture\[12\] _03913_ _03914_ _03928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08755_ _03869_ _03870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05201__A2 _00715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09479__A1 _02559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07706_ _03002_ cpu.regs\[4\]\[4\] _03022_ _03029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05967_ _01328_ _01345_ _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_05898_ _01380_ _01035_ _01371_ _01381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08686_ _03808_ _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07637_ cpu.regs\[7\]\[2\] _02981_ _02986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07568_ cpu.regs\[11\]\[7\] _02931_ _02944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06519_ _01995_ _01397_ _01690_ _01996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_76_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09307_ _04301_ _04329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07499_ _01132_ _02885_ _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09238_ _01268_ _04258_ _04262_ _04263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_90_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09169_ _03201_ _04201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_8_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06768__A2 _00933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output71_I net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10013_ cpu.ROM_addr_buff\[9\] _02484_ _02452_ _04958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_99_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09890__A1 _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08292__I _03517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07636__I _01582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06870_ _02097_ _02346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05821_ _01301_ _01302_ _01304_ _01305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_77_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05752_ cpu.timer_capture\[0\] _01235_ _01236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08540_ cpu.toggle_ctr\[9\] _03704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_106_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08471_ _02051_ _03651_ _03654_ _03653_ _00313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__07304__C _02724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05683_ _01163_ _01165_ _01166_ _01167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07422_ cpu.uart.divisor\[10\] _02829_ _02832_ _02608_ _02833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_106_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05498__A2 _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09633__A1 _02513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07353_ _02293_ _02772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_115_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07284_ _02710_ _02719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06298__I1 cpu.regs\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06304_ _00983_ _01778_ _01782_ _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_33_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09023_ cpu.orig_IO_addr_buff\[2\] _04075_ _04076_ _02675_ _04088_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06235_ cpu.toggle_top\[4\] _01252_ _01714_ _01254_ _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_32_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06166_ _01640_ _01646_ _01647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05117_ cpu.regs\[0\]\[7\] _00634_ cpu.regs\[2\]\[7\] cpu.regs\[3\]\[7\] _00630_
+ _00631_ _00635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06097_ _01529_ _01531_ _01578_ _01579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09925_ net58 _04880_ _04889_ _04885_ _04890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05422__A2 _00908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05048_ _00568_ _00569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09856_ cpu.pwm_counter\[5\] _03792_ cpu.pwm_counter\[7\] cpu.pwm_counter\[6\] _04838_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_08807_ _03275_ _03914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09787_ _04779_ _04736_ _04780_ _04781_ _04782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06999_ _02419_ _02470_ _02471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08124__A1 _03195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08738_ _02727_ _03848_ _03854_ _03851_ _00380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08669_ _02739_ _03802_ _03807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10631_ _00525_ clknet_leaf_65_wb_clk_i net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09624__A1 _04455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10562_ _00456_ clknet_leaf_77_wb_clk_i cpu.last_addr\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10493_ _00388_ clknet_leaf_25_wb_clk_i cpu.timer\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05661__A2 _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06213__I1 net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08115__A1 _02621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09863__A1 _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06677__A1 cpu.regs\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06677__B2 _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09615__A1 _00591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06020_ _01074_ _01051_ _01197_ _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_70_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05652__A2 _01128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07971_ _03256_ _03258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09710_ _03789_ _04716_ _04717_ _00489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06922_ _02339_ _02340_ _02150_ _02396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09641_ _04623_ _00931_ _04652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06853_ _02216_ _02327_ _02328_ _02329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_93_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09572_ _04068_ _04576_ _04585_ _04348_ _04586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05804_ _01287_ _01288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06784_ _02258_ _02259_ _02260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05735_ cpu.uart.divisor\[0\] _01200_ _01206_ _01218_ _01219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08523_ _03678_ _03691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08454_ _02768_ _03641_ _03642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05666_ _01149_ _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_37_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08385_ _02854_ _03589_ _03570_ _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07405_ cpu.uart.divisor\[9\] _02816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05597_ _01080_ _01081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_45_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07336_ _02759_ _00073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_21_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07267_ _02706_ _00057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09006_ _04060_ _04073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06218_ net2 _01114_ _01089_ _01697_ _01698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_07198_ _02646_ _02647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06149_ _00924_ _01589_ _01629_ _01293_ _01630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_14_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09908_ _04877_ _00527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07148__A2 _02598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09839_ net74 _03748_ _04822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_29_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_24_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_1_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10614_ _00508_ clknet_leaf_74_wb_clk_i cpu.ROM_spi_dat_out\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10545_ _00439_ clknet_leaf_96_wb_clk_i cpu.base_address\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_118_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10476_ _00371_ clknet_leaf_29_wb_clk_i cpu.timer_div_counter\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05634__A2 _01090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_63_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08336__A1 _03514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_69_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05520_ _01002_ _01004_ _01005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_47_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05451_ _00715_ _00924_ _00938_ _00939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08170_ cpu.uart.div_counter\[7\] _03418_ _03419_ _03420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07121_ _00692_ _02583_ _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05382_ _00863_ _00869_ _00871_ _00872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_88_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07052_ _02519_ _00029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_88_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06003_ cpu.toggle_top\[2\] _01485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_23_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07954_ cpu.spi.data_out_buff\[6\] _03230_ _03243_ _03244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06050__A2 _00923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07885_ cpu.spi.div_counter\[3\] _03183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06905_ _02083_ _02096_ _02344_ _02380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09624_ _04455_ _04634_ _04635_ _00766_ _04636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06836_ _02300_ _02308_ _02312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_54_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_37_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_37_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09555_ _04370_ _04555_ _04570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06767_ _00789_ _02243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_93_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05718_ _01044_ _01032_ _01202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08506_ _01033_ _02730_ _03678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_clkbuf_leaf_108_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09486_ _04479_ _04503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06698_ _02172_ _02173_ _02174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08437_ _03629_ _03630_ _03600_ _00303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05649_ _00657_ _01133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_34_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06510__B1 _01985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_102_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08368_ cpu.uart.receive_div_counter\[9\] _03576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08299_ _02863_ _03520_ _03524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07319_ _00987_ _02746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10330_ _00225_ clknet_leaf_47_wb_clk_i cpu.uart.dout\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10261_ _00156_ clknet_leaf_110_wb_clk_i cpu.regs\[6\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10192_ _00087_ clknet_leaf_46_wb_clk_i cpu.uart.receive_counter\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_6_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05455__S _00880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07670__S _02994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07402__C _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput14 io_in[21] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06018__C _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput25 rst_n net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_10528_ _00422_ clknet_leaf_41_wb_clk_i cpu.uart.divisor\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05607__A2 _01090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10459_ _00354_ clknet_leaf_108_wb_clk_i cpu.pwm_counter\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05791__B2 _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07670_ _03006_ cpu.regs\[6\]\[6\] _02994_ _03007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_59_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06621_ _02083_ _02096_ _02097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06552_ cpu.mem_cycle\[0\] _02028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09340_ _04361_ _04362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05503_ _00652_ _00987_ _00988_ _00989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09271_ _00725_ _00772_ _04292_ _04294_ _03624_ _04295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_47_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08222_ _02752_ _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_47_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06483_ _01953_ _01958_ _01960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05434_ _00917_ _00922_ _00923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_31_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08153_ _03325_ _03397_ _03406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05365_ _00854_ _00855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08084_ cpu.uart.div_counter\[1\] _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07104_ _02568_ _00032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07599__A2 _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07035_ net12 _02498_ _02505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05296_ cpu.regs\[2\]\[1\] _00806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_101_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05339__I cpu.PORTB_DDR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08986_ _02845_ _04040_ _04053_ _04050_ _04054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_input33_I sram_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07937_ _03213_ _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_97_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07868_ cpu.timer\[9\] _03167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_39_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09702__C _04124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07799_ _02619_ _03105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09607_ _00832_ _04596_ _04620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06819_ _02292_ _02294_ _02295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09538_ _03071_ _04420_ _04553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08318__C _03474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07287__A1 _02635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09469_ _01860_ _04349_ _04486_ _04355_ _04487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_47_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07039__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10313_ _00208_ clknet_leaf_61_wb_clk_i cpu.spi.data_out_buff\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09149__C _04006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09944__I _04891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05249__I _00762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10244_ _00139_ clknet_leaf_127_wb_clk_i cpu.regs\[8\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10175_ _00008_ clknet_leaf_89_wb_clk_i net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07464__I _02872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05712__I _01195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05150_ cpu.mem_cycle\[1\] cpu.mem_cycle\[0\] _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08778__A1 cpu.timer_capture\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07639__I _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09059__C _04050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07450__B2 _02630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05081_ cpu.regs\[1\]\[5\] _00601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_90_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06005__A2 _01079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08840_ cpu.timer_capture\[15\] _03870_ _03940_ _03820_ _03941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_109_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08771_ _03882_ _03883_ _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05983_ cpu.C _01310_ _01466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07722_ cpu.regs\[3\]\[2\] _03036_ _03039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09522__C _04432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07653_ _02995_ _02996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06604_ _02079_ _02080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09323_ _04344_ _04345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07584_ _02940_ cpu.regs\[10\]\[5\] _02945_ _02954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06535_ _01014_ _02011_ _02012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_90_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09254_ cpu.PC\[0\] _00761_ _04278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_8_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06466_ _00643_ _01289_ _01943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05819__A2 _00799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08205_ _03446_ _03447_ _03321_ _00254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09185_ _01007_ _04212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05417_ _00886_ _00891_ _00897_ _00894_ _00906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_06397_ cpu.uart.divisor\[14\] _01700_ _01875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08136_ _03391_ _03392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05348_ cpu.PORTB_DDR\[0\] net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__07441__B2 cpu.uart.divisor\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08067_ _03324_ _03326_ _03328_ _03330_ _03331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__05069__I _00589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05279_ cpu.regs\[2\]\[0\] _00790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07018_ _02481_ _02486_ _02435_ _02489_ _02490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_101_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09194__A1 cpu.TIE vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07744__A2 _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08969_ _04025_ _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_52_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_52_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09497__A2 _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09004__I _01734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05532__I _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08843__I _03942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10227_ _00122_ clknet_leaf_0_wb_clk_i cpu.regs\[10\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07735__A2 _02058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10158_ _00057_ clknet_leaf_30_wb_clk_i cpu.timer_capture\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_89_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10089_ _05029_ _00556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_89_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09488__A2 _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05442__I _00929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06171__A1 _00950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06538__I _02014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06320_ cpu.uart.dout\[5\] _01369_ _01796_ _01798_ _01081_ _01799_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_85_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06251_ _01730_ _01731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05202_ cpu.base_address\[1\] _00712_ _00716_ _00717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_13_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06182_ _01660_ _01662_ _01663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05133_ cpu.br_rel_dest\[5\] _00650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09941_ cpu.PORTB_DDR\[3\] _04892_ _04901_ _04897_ _04902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05064_ _00583_ _00584_ _00585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05285__I0 cpu.regs\[8\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09176__A1 cpu.ROM_addr_buff\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09872_ _04850_ _00518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08923__A1 _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08823_ cpu.timer\[12\] _03836_ _03881_ _03926_ _03927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__07037__C _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08754_ _03859_ _03869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05966_ _01441_ _01431_ _01444_ _01448_ _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_07705_ _02987_ _03023_ _03028_ _00173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05897_ net22 _01380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08685_ _02755_ _03811_ _03819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07636_ _01582_ _02985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07567_ _02943_ _00120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06518_ cpu.timer_div\[7\] _01995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_76_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09306_ _04327_ _04328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09651__A2 _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09237_ cpu.Z _01099_ _04237_ _04261_ _04262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07498_ _02015_ _02889_ _02897_ _00097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_106_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06449_ _01347_ _01904_ _01924_ _01926_ _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__06465__A2 _01862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09168_ _04187_ _04199_ _04200_ _00464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_50_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08119_ _02621_ _03377_ _00237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09099_ _04022_ _04148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_31_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output64_I net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05728__A1 cpu.PORTB_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10012_ cpu.ROM_addr_buff\[1\] _04950_ _02483_ cpu.ROM_addr_buff\[5\] cpu.ROM_addr_buff\[13\]
+ _02465_ _04957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__08914__A1 _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07189__I _02639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09158__A1 _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05437__I _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05820_ _01303_ _01304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06392__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07652__I _02994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_19_Left_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05751_ _01037_ _01057_ _01234_ _01235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_08470_ cpu.orig_PC\[4\] _03636_ _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05682_ _01150_ _01166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07421_ cpu.uart.receive_div_counter\[0\] _02832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07352_ _01358_ _02764_ _02770_ _02771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06303_ _00982_ _01781_ _01782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_17_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07283_ _02631_ _02711_ _02718_ _02716_ _00061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06298__I2 cpu.regs\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Left_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09022_ _04084_ _04087_ _00431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06234_ _01712_ _01713_ _01714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06165_ _01643_ _01645_ _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_4_3_0_wb_clk_i clknet_0_wb_clk_i clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_41_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05116_ _00633_ _00634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06096_ _01315_ _01547_ _01567_ _01577_ _01578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_09924_ _04052_ _04881_ _04889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05047_ _00000_ _00568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05347__I cpu.PORTA_DDR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09855_ _04830_ _04833_ _04836_ _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_99_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08806_ _03869_ _03913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_37_Left_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09786_ cpu.ROM_spi_dat_out\[0\] _04779_ _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06998_ _02457_ _02470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_14_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07562__I _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06383__A1 _00982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08737_ cpu.timer_top\[15\] _03849_ _03854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05949_ _01426_ _01431_ _01432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08668_ _03806_ _00358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07619_ _02972_ _00143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10630_ _00524_ clknet_leaf_68_wb_clk_i net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_95_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08599_ _03751_ _03759_ _00336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_24_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_46_Left_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10561_ _00455_ clknet_leaf_79_wb_clk_i cpu.ROM_addr_buff\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10492_ _00387_ clknet_leaf_26_wb_clk_i cpu.timer\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05661__A3 _01144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06297__S1 _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05949__A1 _01426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_53_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_55_Left_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09560__A1 _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_101_Right_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_64_Left_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05720__I _01203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_92_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07970_ _03252_ _03254_ _03256_ _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_73_Left_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05167__I _00682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06921_ _02379_ _02378_ _02394_ _02395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_87_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09640_ _04623_ _00931_ _04651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06852_ _02185_ _02186_ _02328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06365__A1 _01441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_109_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_109_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09571_ _03070_ _04484_ _04585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05803_ _01286_ _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06783_ _02231_ _02232_ _02259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06117__A1 net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05734_ _01214_ _01215_ _01217_ _01088_ _01218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_89_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09303__A1 _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08522_ _03678_ _03690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08453_ _03621_ _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07404_ _01866_ _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_93_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05665_ _01147_ _01071_ _01148_ _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08384_ _03585_ _03581_ _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05630__I _01113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05596_ _01076_ _01079_ _01080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_58_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07335_ cpu.toggle_top\[15\] _02745_ _02758_ _02753_ _02759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_21_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07266_ cpu.timer_capture\[7\] _02684_ _02705_ _02689_ _02706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_33_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06217_ _01378_ _01695_ _01696_ _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09005_ _04071_ _04072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07197_ _01785_ _02646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06148_ _00966_ _01273_ _01277_ _01628_ _01629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06079_ _01454_ _00908_ _01561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09907_ net81 _04869_ _04876_ _04874_ _04877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07493__S _02886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09542__A1 _04530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09838_ _03288_ _04818_ _04821_ _00513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__05403__I0 cpu.regs\[8\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09769_ _02439_ _04735_ _04749_ _04764_ _04765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_57_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10613_ _00507_ clknet_leaf_75_wb_clk_i cpu.ROM_spi_dat_out\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07608__A1 cpu.regs\[8\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10544_ _00438_ clknet_leaf_84_wb_clk_i cpu.base_address\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10475_ _00370_ clknet_leaf_28_wb_clk_i cpu.timer_div_counter\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_118_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05890__I0 cpu.PORTA_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_7_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_7_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_9_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06595__A1 _00589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05450_ _00932_ _00937_ _00912_ _00938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05381_ _00870_ _00871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07120_ _02581_ _02582_ _02583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_70_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_81_Left_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_70_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07051_ _02513_ _02496_ _02515_ _02518_ _02519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_42_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06002_ _01153_ _01165_ _01166_ _01484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09221__B1 _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05389__A2 _00878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07953_ _02646_ _03242_ _03243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07884_ cpu.spi.divisor\[7\] _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09524__A1 _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06904_ _02336_ _02343_ _02379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06338__A1 _01774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09623_ _04309_ _04625_ _04635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06835_ _02307_ _02310_ _02311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_54_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07840__I cpu.timer_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09554_ _04329_ _04555_ _04568_ _04366_ _04569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06766_ _02226_ _02236_ _02242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05717_ net6 _01201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08505_ _03677_ _00739_ _00324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09485_ _04501_ _04502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06697_ _02168_ _02169_ _02173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_38_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_77_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_77_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08157__B _03276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08436_ cpu.orig_IO_addr_buff\[6\] _03627_ _03630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05648_ _01109_ _01131_ _01132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_34_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08367_ _03552_ _03575_ _00288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06510__B2 _01986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05579_ _01038_ _01047_ _01053_ _01062_ _01063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07318_ _02731_ _02745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08298_ _03522_ _03523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08263__A1 _03231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07249_ cpu.timer\[5\] _02691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10260_ _00155_ clknet_leaf_13_wb_clk_i cpu.regs\[6\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10191_ _00086_ clknet_leaf_46_wb_clk_i cpu.uart.receive_counter\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_6_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09118__I1 cpu.ROM_addr_buff\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput15 io_in[23] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput26 sram_out[0] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10527_ _00012_ clknet_leaf_44_wb_clk_i cpu.uart.clr_hb vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_12_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05458__I3 cpu.regs\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07197__I _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10458_ _00353_ clknet_leaf_16_wb_clk_i cpu.pwm_counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10389_ _00284_ clknet_leaf_38_wb_clk_i cpu.uart.receive_div_counter\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05240__A1 _00653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06620_ _02092_ _02095_ _02096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06477__S _00871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06551_ _02026_ _02027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_87_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08493__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05502_ _00968_ _00980_ _00988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09270_ _00724_ _04293_ _04294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06482_ _01953_ _01958_ _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08221_ _03459_ cpu.uart.counter\[1\] _03454_ _03460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05180__I net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05433_ _00919_ _00921_ _00922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08152_ _03387_ _03405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05364_ _00004_ _00854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08083_ _02828_ _03344_ cpu.uart.div_counter\[8\] _02831_ _03346_ _03347_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_70_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05295_ _00804_ _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07103_ _02373_ _02567_ _02543_ _02568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07034_ _02504_ _00026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08548__A2 cpu.toggle_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_124_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_124_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08985_ _04052_ _04042_ _04053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07936_ _03220_ _03227_ _03229_ _00203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input26_I sram_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05355__I _00844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07867_ cpu.timer\[10\] _03166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07798_ _03103_ _03104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09606_ _04594_ _04603_ _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06818_ _02293_ _00974_ _02294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_104_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09537_ _03045_ _04500_ _04552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06749_ _02223_ _02224_ _02225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08484__A1 _03045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09468_ _04350_ _04473_ _04485_ _04353_ _04486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08419_ _01031_ _03610_ _03616_ _03613_ _00299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09399_ _04418_ _04379_ _04419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09984__A1 cpu.PORTA_DDR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output94_I net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10312_ _00207_ clknet_leaf_61_wb_clk_i cpu.spi.data_out_buff\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06798__A1 _02270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10243_ _00138_ clknet_leaf_4_wb_clk_i cpu.regs\[8\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09165__C _04006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10174_ _00073_ clknet_leaf_12_wb_clk_i cpu.toggle_top\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05222__A1 _00734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09960__I _04914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05525__A2 _01008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06722__A1 cpu.regs\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07480__I _02886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07770__I0 _01582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05080_ cpu.regs\[4\]\[5\] cpu.regs\[5\]\[5\] cpu.regs\[6\]\[5\] cpu.regs\[7\]\[5\]
+ _00598_ _00599_ _00600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_0_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08770_ cpu.timer_capture\[3\] _03870_ _03437_ _03883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05982_ _00800_ _01340_ _01465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07721_ _01481_ _03035_ _03038_ _00179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06713__A1 _00589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07652_ _02994_ _02995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06603_ _02077_ _02078_ _02079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07583_ _02953_ _00126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_87_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09322_ _04313_ _04344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06534_ _01133_ _01172_ _02010_ _02011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09253_ _04276_ _04277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06465_ _01937_ _01862_ _01942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06396_ _01866_ _01370_ _01872_ _01873_ _01700_ _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_08204_ _03329_ _03439_ _03398_ _03440_ _03447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_90_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09184_ _04201_ _04210_ _04211_ _00469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05416_ _00905_ net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_62_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08135_ _03331_ _03357_ _03364_ _03391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__09966__A1 cpu.PORTA_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05347_ cpu.PORTA_DDR\[2\] net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_70_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08066_ cpu.uart.divisor\[14\] _03329_ cpu.uart.div_counter\[13\] _02814_ _03330_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_31_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05278_ cpu.regs\[1\]\[0\] _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07017_ _02488_ _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07565__I _01934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08968_ _04039_ _00425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07919_ cpu.spi.data_out_buff\[0\] _03214_ _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08899_ cpu.spi.divisor\[3\] _03984_ _03988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_92_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_92_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05063__S0 _00571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05813__I _01296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_21_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_21_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_66_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06180__A2 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07680__A2 _03012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10226_ _00121_ clknet_leaf_126_wb_clk_i cpu.regs\[11\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06312__C _01121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10157_ _00056_ clknet_leaf_29_wb_clk_i cpu.timer_capture\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_55_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10088_ _01262_ _04997_ _05028_ _04931_ _05029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07499__A2 _02885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08448__A1 _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06250_ _01729_ _01730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09948__A1 _04045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05201_ _00713_ _00715_ _00716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09865__I _04843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07586__S _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06181_ _01554_ _01661_ _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10009__C _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05132_ net25 _00649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_110_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09940_ _04037_ _04893_ _04901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05063_ cpu.regs\[4\]\[4\] cpu.regs\[5\]\[4\] cpu.regs\[6\]\[4\] cpu.regs\[7\]\[4\]
+ _00571_ _00576_ _00584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_115_Right_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05985__A2 _01001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09871_ net60 _04844_ _04848_ _04849_ _04850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_96_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08822_ _03856_ _03924_ _03925_ _03926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08753_ _03863_ _03867_ _03868_ _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05965_ _01445_ _01447_ _01448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07704_ cpu.regs\[4\]\[3\] _03022_ _03028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05896_ _01070_ _01376_ _01377_ _01378_ _01379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_08684_ _03818_ _00362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07635_ _02983_ _02980_ _02984_ _00147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07566_ _02942_ cpu.regs\[11\]\[6\] _02930_ _02943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06517_ _01981_ _01187_ _01992_ _01993_ _01184_ _01994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_09305_ _04284_ _04327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_35_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08165__B _03276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09236_ _01003_ _04259_ _01265_ _01290_ _04260_ _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__06464__I _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07497_ cpu.regs\[14\]\[7\] _02887_ _02897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07111__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06448_ _01447_ _01925_ _01926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09167_ cpu.last_addr\[8\] _04192_ _04200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06379_ _01857_ _01858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08118_ _03098_ _03367_ _03376_ _03371_ _03377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09098_ cpu.ROM_addr_buff\[6\] _04147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_43_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08049_ cpu.uart.dout\[5\] _03309_ _03316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07295__I _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05976__A2 _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10011_ net72 _04956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05728__A2 _01211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output57_I net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09443__C _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09015__I _04081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07102__A1 _02556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_82_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10209_ _00104_ clknet_leaf_121_wb_clk_i cpu.regs\[13\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05750_ _01061_ _01234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_77_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08669__A1 _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05681_ _01164_ _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07420_ cpu.uart.divisor\[8\] _02831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XTAP_TAPCELL_ROW_85_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07351_ _02768_ _02524_ _02542_ _02769_ _02770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_06302_ _01779_ _01780_ _00851_ _01781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07282_ cpu.timer_top\[3\] _02712_ _02718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09021_ _01054_ _04067_ _04086_ _04082_ _04087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06233_ cpu.pwm_top\[4\] _01619_ _01125_ _01713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06164_ _01539_ _01543_ _01644_ _01645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05115_ cpu.regs\[1\]\[7\] _00633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06095_ _01569_ _01570_ _01573_ _01576_ _01577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_40_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09923_ _04888_ _00531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05046_ _00566_ _00567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_clkbuf_4_12_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09854_ cpu.pwm_top\[1\] _04826_ _04834_ cpu.pwm_top\[2\] _04835_ _04836_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA_clkbuf_leaf_127_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07843__I cpu.timer_top\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08805_ _03909_ _03894_ _03904_ _03911_ _03898_ _03912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_09785_ _04770_ _04780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06997_ _02420_ _02468_ _02469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06383__A2 _01281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08736_ _02647_ _03848_ _03853_ _03851_ _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05363__I _00852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05948_ _01333_ _01430_ _01431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08667_ cpu.pwm_top\[1\] _03801_ _03805_ _03697_ _03806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05879_ _01160_ _01360_ _01362_ _00013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_71_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07618_ _02940_ cpu.regs\[8\]\[5\] _02963_ _02972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_83_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08598_ _03731_ _03757_ _03759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_24_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07549_ _02931_ _02932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_101_Left_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10560_ _00454_ clknet_leaf_88_wb_clk_i cpu.ROM_addr_buff\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07635__A2 _02980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10491_ _00386_ clknet_leaf_27_wb_clk_i cpu.timer\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05646__A1 _01110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09219_ _01135_ _02271_ _04244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_80_Right_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09454__B _04417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10689_ net49 net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06920_ _02372_ _02377_ _02394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07663__I _01771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09551__A2 _04359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05799__S1 _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06851_ _02241_ _02325_ _02326_ _02327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_93_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09570_ _04456_ _04582_ _04583_ _04396_ _04584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06782_ _02247_ _02248_ _02257_ _02258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05802_ _01281_ _01285_ _00896_ _01286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05733_ net21 _01216_ _01217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08521_ _03689_ _00328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08452_ _03132_ _03618_ _03640_ _03620_ _00308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_26_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07403_ cpu.uart.divisor\[13\] _02814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_05664_ _00707_ cpu.instr_buff\[14\] _00682_ _01008_ _01148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_08383_ cpu.uart.receive_div_counter\[12\] _03585_ _03581_ _03588_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_92_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05595_ _01075_ _01078_ _01079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_58_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07334_ _02652_ _02747_ _02758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_21_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07265_ _02703_ _02686_ _02674_ _02704_ _02705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06216_ net63 _01213_ _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09004_ _01734_ _04071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07196_ _02645_ _00047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06147_ _01269_ _01627_ _01628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05358__I _00712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06078_ _01559_ _01560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09906_ _04851_ _04870_ _04876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07573__I _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09837_ _02415_ _04806_ _04820_ _04821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__06410__C _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07553__A1 cpu.regs\[11\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09768_ _02431_ _02438_ _04743_ cpu.startup_cycle\[0\] _04764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_57_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05093__I _00612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05403__I1 cpu.regs\[9\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08719_ cpu.timer_top\[8\] _03842_ _03843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09699_ _04684_ _04686_ _04687_ _04708_ _04709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_69_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06917__I _02360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09058__A1 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10612_ _00506_ clknet_leaf_74_wb_clk_i cpu.ROM_spi_dat_out\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10543_ _00437_ clknet_leaf_56_wb_clk_i cpu.IO_addr_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10474_ _00369_ clknet_leaf_28_wb_clk_i cpu.timer_div_counter\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08569__B1 cpu.toggle_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06044__A1 _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06595__A2 _01955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06320__C _01081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05217__B _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09297__A1 _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05858__B2 _01340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05380_ _00007_ _00870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07050_ _02517_ _02518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_70_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06001_ _01160_ _01482_ _01483_ _00014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10084__I _05017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09221__B2 _01365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09221__A1 _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09873__I _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06035__A1 cpu.timer_top\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07952_ _03211_ _03242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07883_ _03180_ _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06903_ _02372_ _02377_ _02378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07535__A1 cpu.regs\[12\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09622_ _03672_ _00931_ _04633_ _04634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06834_ _02300_ _02308_ _02309_ _02310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09553_ _04561_ _04565_ _04567_ _04568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_54_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08504_ cpu.toggle_clkdiv _03677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06765_ _02238_ _02240_ _02241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05716_ _01199_ _01200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_77_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09484_ _02569_ _04498_ _04500_ _04501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06696_ _02171_ _02154_ _02172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08435_ cpu.IO_addr_buff\[6\] _03622_ _03629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05647_ _01130_ _01131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__05849__A1 _00799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08366_ _02830_ _03563_ _03553_ _03574_ _03575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06510__A2 _01035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08952__I _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05578_ _01057_ _01061_ _01062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_46_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07317_ _02744_ _00069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08297_ _03516_ _03521_ _03522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_46_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06274__A1 _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_46_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_46_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07248_ _02690_ _00054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_104_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07179_ _00952_ _02631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09212__A1 _00909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06026__A1 cpu.spi.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10190_ _00085_ clknet_leaf_14_wb_clk_i _00003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_6_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05551__I _01034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06888__I0 _00591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput16 io_in[26] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput27 sram_out[1] net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09451__A1 _02370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10526_ _00421_ clknet_leaf_88_wb_clk_i cpu.rom_data_dist vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06265__A1 _01586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05312__I0 cpu.regs\[12\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06315__C _01793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10457_ _00352_ clknet_leaf_108_wb_clk_i cpu.pwm_counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06017__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10388_ _00283_ clknet_leaf_37_wb_clk_i cpu.uart.receive_div_counter\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05240__A2 _00656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06550_ _02025_ _02026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_114_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05501_ _00986_ _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06481_ _01895_ _01957_ _01925_ _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08220_ _03452_ _03459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08493__A2 _03611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05432_ _00887_ _00920_ _00896_ _00921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_117_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08151_ _03402_ _03404_ _00243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09442__A1 _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05363_ _00852_ _00853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_28_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08082_ _02828_ _03344_ _03345_ _02608_ _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_99_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05294_ cpu.regs\[1\]\[1\] _00804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06292__I _01771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07102_ _02556_ _02521_ _02566_ _02567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07033_ _00760_ _02496_ _02500_ _02503_ _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_30_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07756__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08984_ _02651_ _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07935_ cpu.spi.data_out_buff\[1\] _03223_ _03228_ _03229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08947__I _04022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07866_ cpu.timer_top\[7\] _02703_ _03164_ _03165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09605_ _04382_ _04603_ _04617_ _04406_ _04618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input19_I io_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07797_ _03100_ _03103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06817_ _02243_ _02293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_104_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09536_ _03664_ _04550_ _04551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06748_ _00831_ _00974_ _02224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09467_ _02558_ _04484_ _04485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08418_ cpu.orig_IO_addr_buff\[2\] _03615_ _03616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06679_ _02152_ _02153_ _02154_ _02155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_93_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09398_ cpu.PC\[4\] _04418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08349_ _03556_ _03559_ _03437_ _03562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_104_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06247__A1 _00596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10311_ _00206_ clknet_leaf_60_wb_clk_i cpu.spi.data_out_buff\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06798__A2 _00976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10242_ _00137_ clknet_leaf_119_wb_clk_i cpu.regs\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10173_ _00072_ clknet_leaf_12_wb_clk_i cpu.toggle_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05222__A2 _00735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09018__I _03551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10106__I0 _01771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07770__I1 _03078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06486__A1 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06238__B2 _00950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10509_ _00404_ clknet_leaf_8_wb_clk_i cpu.timer_capture\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05997__B1 _01477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05461__A2 _00943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05981_ _01429_ _01440_ _01449_ _01463_ _01464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_07720_ cpu.regs\[3\]\[1\] _03036_ _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07651_ _02405_ _02977_ _02994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06602_ _00602_ _01956_ _02078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07582_ _02938_ cpu.regs\[10\]\[4\] _02946_ _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_87_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06533_ _01115_ _02007_ _02009_ _02010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09321_ _04337_ _04340_ _04342_ _04343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09252_ _00734_ _00651_ _04276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_44_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06464_ _01640_ _01941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_8_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06395_ net13 _01372_ _01200_ _01873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_106_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08203_ cpu.uart.div_counter\[14\] _03445_ _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09183_ cpu.last_addr\[13\] _04176_ _04211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05415_ _00847_ _00879_ _00904_ _00905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__09415__A1 _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08134_ _03385_ _03390_ _03321_ _00240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06229__A1 cpu.timer_capture\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05346_ cpu.PORTA_DDR\[1\] net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_55_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08065_ cpu.uart.div_counter\[14\] _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_33_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07846__I cpu.timer_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05277_ _00002_ _00787_ _00788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07016_ _02487_ _02488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08967_ cpu.uart.divisor\[11\] _04026_ _04038_ _04035_ _04039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08154__A1 _03333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07918_ _03213_ _03214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08898_ _02627_ _03983_ _03987_ _00407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07849_ _03134_ cpu.timer\[13\] _03148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05063__S1 _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09519_ _04530_ _04533_ _04534_ _04535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_38_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_72_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_61_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_61_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_81_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05979__B1 _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10225_ _00120_ clknet_leaf_121_wb_clk_i cpu.regs\[11\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10156_ _00055_ clknet_leaf_29_wb_clk_i cpu.timer_capture\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10087_ _04575_ _05009_ _05027_ _04997_ _05028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09893__A1 _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05225__B _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09645__A1 _04121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05506__I0 _00990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05200_ _00714_ _00715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_105_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10159__CLK clknet_leaf_18_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06180_ _01152_ net92 _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05131_ cpu.instr_cycle\[2\] _00648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07666__I _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05062_ _00581_ _00583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09870_ _04123_ _04849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09881__I _04843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08821_ _03921_ _03916_ cpu.timer\[12\] _03925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_117_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08752_ _03649_ _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05964_ _01446_ _01447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08683_ cpu.pwm_top\[5\] _03814_ _03817_ _03809_ _03818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07703_ _02985_ _03023_ _03027_ _00172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05895_ _01113_ _01378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07634_ cpu.regs\[7\]\[1\] _02981_ _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09636__A1 _03674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07565_ _01934_ _02942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06516_ cpu.spi.divisor\[7\] _01189_ _01608_ _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09304_ _04326_ _00474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07496_ _02896_ _00096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09235_ _01264_ _01272_ _04260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06447_ _01831_ _01909_ _01910_ _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09166_ cpu.ROM_addr_buff\[8\] _04194_ _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05673__A2 _01145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06378_ _01357_ _01817_ _01856_ _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_08117_ _03098_ _03375_ _03376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09097_ cpu.regs\[2\]\[6\] _02559_ _04130_ _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_71_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05329_ cpu.regs\[8\]\[3\] cpu.regs\[9\]\[3\] cpu.regs\[10\]\[3\] cpu.regs\[11\]\[3\]
+ _00569_ _00827_ _00837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08048_ cpu.uart.receive_buff\[5\] _03307_ _03315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07670__I0 _03006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10010_ _04955_ _00551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09999_ _04944_ _04945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09875__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09627__A1 _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06861__A1 _00603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08366__A1 _02830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10208_ _00103_ clknet_leaf_124_wb_clk_i cpu.regs\[13\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05719__A3 _01202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10139_ _00038_ clknet_leaf_108_wb_clk_i cpu.br_rel_dest\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09866__A1 _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05680_ _01106_ _01164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_85_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09618__A1 _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07350_ _02392_ _02299_ _02529_ _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06301_ cpu.regs\[8\]\[6\] cpu.regs\[9\]\[6\] cpu.regs\[10\]\[6\] cpu.regs\[11\]\[6\]
+ _01775_ _01282_ _01780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_18_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07281_ _02627_ _02711_ _02717_ _02716_ _00060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09020_ _01365_ _04070_ _04072_ _04085_ _04079_ _04086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA_rebuffer9_I _00854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06232_ cpu.timer_top\[12\] _01247_ _01621_ _01711_ _01712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__05655__A2 _01065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06163_ _01152_ _01531_ _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05114_ cpu.regs\[4\]\[7\] cpu.regs\[5\]\[7\] cpu.regs\[6\]\[7\] cpu.regs\[7\]\[7\]
+ _00630_ _00631_ _00632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05407__A2 _00895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06094_ _01574_ _01575_ _01576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09922_ net57 _04880_ _04887_ _04885_ _04888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05045_ _00003_ _00566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09853_ cpu.pwm_top\[3\] cpu.pwm_counter\[3\] _04835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09784_ _02488_ _04779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08804_ _03909_ _03910_ _03911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06996_ _02429_ _02435_ _02441_ _02467_ _02468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_08735_ cpu.timer_top\[14\] _03849_ _03853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05947_ _00814_ _00900_ _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08666_ _02735_ _03802_ _03805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05878_ cpu.regs\[9\]\[0\] _01361_ _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09609__A1 _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08597_ _03756_ _03757_ _03758_ _00335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07617_ _02971_ _00142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05894__A2 _01070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07548_ _02930_ _02931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_52_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07096__A1 _02559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07479_ _02405_ _02885_ _02886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_10490_ _00385_ clknet_leaf_27_wb_clk_i cpu.timer\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09218_ _01153_ _02796_ _04243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09149_ _04184_ _04172_ _04186_ _04006_ _00459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_102_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06385__I _01862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05637__A2 _01120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05729__I _01068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06850_ _02215_ _02214_ _02326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__05464__I _00951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05801_ _01283_ _01284_ _00852_ _01285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06781_ _02255_ _02256_ _02257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05732_ _01034_ _01216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_89_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08520_ cpu.toggle_top\[3\] _03679_ _03688_ _03686_ _03689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08451_ cpu.orig_flags\[3\] _03636_ _03640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05663_ _00716_ _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06509__B _01216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07402_ _02595_ _02811_ _02607_ _02813_ _00085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_08382_ _03580_ _03587_ _00291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05594_ _01049_ _01077_ _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_73_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07333_ _02757_ _00072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_21_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07264_ _02661_ _01291_ _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_118_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_118_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06215_ _01374_ _01693_ _01694_ _01121_ _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_09003_ _04069_ _04070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07195_ cpu.uart.divisor\[5\] _02623_ _02644_ _02640_ _02645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06146_ _01174_ _01623_ _01626_ _01260_ _00936_ _01627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_14_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06077_ _01533_ _01534_ _01559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09905_ _04875_ _00526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09836_ _04809_ _00660_ _04819_ _04820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05374__I _00854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09767_ _04743_ _04734_ _04748_ _04763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06979_ _02026_ _02450_ _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_57_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05403__I2 cpu.regs\[10\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09698_ cpu.last_addr\[13\] _04682_ _04688_ _04707_ _04708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_08718_ _03840_ _03842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_107_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08649_ _03792_ _03791_ _03793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_1_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10611_ _00505_ clknet_leaf_74_wb_clk_i cpu.ROM_spi_dat_out\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10542_ _00436_ clknet_leaf_55_wb_clk_i cpu.IO_addr_buff\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05619__A2 _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05977__C _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10473_ _00368_ clknet_leaf_28_wb_clk_i cpu.timer_div_counter\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07616__I0 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09297__A2 _04319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05858__A2 _01336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06000_ cpu.regs\[9\]\[1\] _01361_ _01483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08980__A1 _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07951_ _03235_ _03240_ _03241_ _00206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06902_ _02374_ _02376_ _02377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07882_ cpu.spi.div_counter\[2\] _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08732__A1 _02635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09621_ _04631_ _04632_ _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06833_ _02270_ _00908_ _02309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09552_ _04358_ _04555_ _04566_ _04439_ _04567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06764_ _02239_ _02240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08503_ _02621_ _03603_ _00323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05715_ _01036_ _01198_ _01199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_54_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09288__A2 _01364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09483_ _04499_ _04500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06695_ _02152_ _02153_ _02171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07342__C _02763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08434_ _03623_ _03628_ _03600_ _00302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_19_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05849__A2 _01309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05646_ _01110_ _01014_ _01129_ _01130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08365_ _02830_ _03571_ _03574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05577_ _01060_ _01061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_18_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08799__A1 _03170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07316_ cpu.toggle_top\[11\] _02732_ _02743_ _02737_ _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08296_ _02863_ _03520_ _03515_ _03521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_6_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07247_ cpu.timer_capture\[4\] _02684_ _02688_ _02689_ _02690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_61_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07178_ cpu.uart.divisor\[3\] _02630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09212__A2 _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06129_ cpu.spi.dout\[3\] _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07223__A1 _02668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_86_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_86_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_15_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_15_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05785__A1 _00656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10662__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09819_ _04806_ _04807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08723__A1 _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput17 io_in[28] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput28 sram_out[2] net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_52_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10525_ _00420_ clknet_leaf_30_wb_clk_i cpu.timer_div\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06265__A2 net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09974__I _04914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10456_ _00351_ clknet_leaf_108_wb_clk_i cpu.pwm_counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10387_ _00282_ clknet_leaf_39_wb_clk_i cpu.uart.receive_div_counter\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05320__S0 _00570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06480_ _01956_ _01957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05500_ _00985_ _00986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05898__B _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05431_ cpu.regs\[12\]\[2\] cpu.regs\[13\]\[2\] cpu.regs\[14\]\[2\] cpu.regs\[15\]\[2\]
+ _00856_ _00860_ _00920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_08150_ cpu.uart.div_counter\[3\] _03389_ _03403_ _03384_ _03404_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_7_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05362_ _00851_ _00852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_16_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07101_ _02557_ _02561_ _02565_ _02531_ _02566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08081_ cpu.uart.div_counter\[0\] _03345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__06500__I0 net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10095__I _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05293_ cpu.regs\[4\]\[1\] cpu.regs\[5\]\[1\] cpu.regs\[6\]\[1\] cpu.regs\[7\]\[1\]
+ _00801_ _00802_ _00803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07032_ _02502_ _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_70_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_23_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07205__A1 _02652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07756__A2 _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08983_ _04051_ _00428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07934_ _03111_ _03228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07865_ _01980_ cpu.timer\[7\] _03163_ _03164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09604_ _04605_ _04616_ _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_39_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07796_ _03101_ _03102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06816_ _02157_ _02290_ _02291_ _02292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_104_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09535_ _04296_ _04550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06747_ _00900_ _02219_ _02222_ _02223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09466_ _04055_ _04484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06678_ _00601_ _00933_ _02154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_19_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_62_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05629_ _01087_ _01112_ _01113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08417_ _03608_ _03615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_80_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09397_ _04380_ _04416_ _04417_ _00476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08348_ _03556_ _03557_ _03558_ _03560_ _03561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08279_ cpu.uart.data_buff\[7\] _03465_ _03507_ _03508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06247__A2 _00985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10310_ _00205_ clknet_leaf_60_wb_clk_i cpu.spi.data_out_buff\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05099__I cpu.regs\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10241_ _00136_ clknet_leaf_114_wb_clk_i cpu.regs\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05758__A1 _01094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10172_ _00071_ clknet_leaf_12_wb_clk_i cpu.toggle_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05222__A3 _00736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06183__A1 _01144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05930__A1 _00878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09121__A1 _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10508_ _00403_ clknet_leaf_8_wb_clk_i cpu.timer_capture\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05297__I0 cpu.regs\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10439_ _00334_ clknet_leaf_7_wb_clk_i cpu.toggle_ctr\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_107_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05980_ _01462_ _01463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_85_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07650_ _02992_ _02981_ _02993_ _00153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06601_ _02075_ _02076_ _02077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07581_ _02922_ _02947_ _02952_ _00125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06532_ _01419_ _01270_ _01721_ _02008_ _02009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09320_ _04337_ _04340_ _04341_ _04342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09251_ _02765_ _04274_ _04275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08202_ _03393_ _03444_ _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06463_ _01851_ _01906_ _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06394_ net4 _01114_ _01089_ _01871_ _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_09182_ cpu.ROM_addr_buff\[13\] _04185_ _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05414_ _00903_ _00904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_62_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08133_ _03350_ _03389_ _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05345_ cpu.PORTA_DDR\[0\] net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_114_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08064_ _02845_ _03327_ cpu.uart.div_counter\[14\] _02847_ _03328_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_71_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07015_ _00661_ _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09179__A1 cpu.ROM_addr_buff\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05276_ cpu.regs\[4\]\[0\] cpu.regs\[5\]\[0\] cpu.regs\[6\]\[0\] cpu.regs\[7\]\[0\]
+ _00785_ _00786_ _00787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08926__A1 _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input31_I sram_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08966_ _04037_ _04028_ _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07917_ _03210_ _03213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08897_ cpu.spi.divisor\[2\] _03984_ _03987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07848_ _03141_ _03144_ _03146_ _03147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07811__B _03112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07779_ _02044_ net115 _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_38_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09518_ _04530_ _04533_ _04341_ _04534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_65_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09449_ _04383_ _04452_ _04467_ _04407_ _04468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_38_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09406__A2 _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09738__B _00778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_30_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_30_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10224_ _00119_ clknet_leaf_116_wb_clk_i cpu.regs\[11\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10155_ _00054_ clknet_leaf_30_wb_clk_i cpu.timer_capture\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10086_ _05015_ _05024_ _05026_ _04327_ _05027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05292__I _00786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07408__A1 _02816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05130_ _00646_ _00647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06631__A2 _02064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05061_ _00577_ _00578_ _00581_ _00582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05285__I3 cpu.regs\[11\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08908__A1 _02647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08820_ cpu.timer\[12\] _03921_ _03916_ _03924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_21_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08751_ cpu.timer_capture\[0\] _03866_ _03867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05963_ _00969_ _00929_ _01346_ _01446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_05894_ net60 _01070_ _01377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08682_ _02750_ _03811_ _03817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_49_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07702_ cpu.regs\[4\]\[2\] _03024_ _03027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07633_ _01480_ _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_88_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07564_ _02941_ _00119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06515_ cpu.uart.dout\[7\] _01369_ _01081_ _01991_ _01992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_09303_ _02783_ _04212_ _04325_ _04124_ _04326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07495_ _01935_ cpu.regs\[14\]\[6\] _02886_ _02896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_90_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09234_ _00743_ _01259_ _04259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06446_ _01831_ _01910_ _01909_ _01924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_17_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09165_ _04197_ _04172_ _04198_ _04006_ _00463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_63_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08116_ cpu.spi.counter\[0\] cpu.spi.counter\[1\] _03099_ _03375_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_44_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06377_ net31 _01425_ _01478_ _01855_ _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_31_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09096_ _04145_ _00447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05328_ _00586_ _00835_ _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08047_ _03313_ _03314_ _03312_ _00229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_101_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05259_ _00725_ _00771_ _00772_ cpu.instr_cycle\[3\] _00773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_112_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05377__I _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09572__A1 _04068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09998_ _02470_ _00692_ _02468_ _02487_ _04944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_08949_ _00728_ _04023_ _04024_ _00421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09312__I _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05664__A3 _00682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06613__A2 _01955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06377__A1 net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10207_ _00102_ clknet_leaf_120_wb_clk_i cpu.regs\[13\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10138_ _00037_ clknet_4_10_0_wb_clk_i cpu.br_rel_dest\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10069_ _01937_ _01948_ _05010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_82_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07280_ cpu.timer_top\[2\] _02712_ _02717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06300_ cpu.regs\[12\]\[6\] cpu.regs\[13\]\[6\] cpu.regs\[14\]\[6\] cpu.regs\[15\]\[6\]
+ _01775_ _01282_ _01779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_73_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06231_ _01689_ _01616_ _01709_ _01710_ _01246_ _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_26_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07677__I _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06162_ _01641_ _01642_ _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05113_ _00599_ _00631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06093_ _01549_ _01572_ _01575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09921_ _04048_ _04881_ _04887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05197__I cpu.base_address\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09852_ _03786_ _04834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09783_ _04770_ _04778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08803_ cpu.timer\[8\] _03905_ _03910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06995_ _02453_ _02455_ _02466_ _02467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08734_ _02643_ _03848_ _03852_ _03851_ _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05946_ _01427_ _01428_ _01429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_96_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08457__B _03633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08665_ _03804_ _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05877_ _01159_ _01361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06915__I0 _00604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08596_ cpu.toggle_ctr\[2\] _03754_ _03758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07616_ _02938_ cpu.regs\[8\]\[4\] _02964_ _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_62_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07547_ _01158_ _02929_ _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_91_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08293__A1 _03514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08971__I _04025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07478_ _01138_ _01156_ _02884_ _02885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_118_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06429_ _01851_ _01906_ _01907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09217_ _01587_ _02093_ _04242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09148_ cpu.ROM_addr_buff\[3\] _04185_ _04186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09079_ _04132_ _00443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_15_Left_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output62_I net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06359__A1 _01329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05582__A2 _01055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_24_Left_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_33_Left_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09536__A1 _03664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_42_Left_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05800_ cpu.regs\[0\]\[7\] cpu.regs\[1\]\[7\] cpu.regs\[2\]\[7\] cpu.regs\[3\]\[7\]
+ _00855_ _01282_ _01284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09839__A2 _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06780_ _02248_ _02247_ _02256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05731_ net59 _01122_ _01113_ _01215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08450_ _03638_ _03639_ _03633_ _00307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05662_ _01020_ _01146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08381_ _03585_ _03563_ _03558_ _03586_ _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07401_ _02592_ _02811_ _02605_ _02813_ _00084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__05480__I _00966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05593_ _00645_ _01077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07332_ cpu.toggle_top\[14\] _02745_ _02756_ _02753_ _02757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_18_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_51_Left_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07263_ cpu.timer\[7\] _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_45_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06214_ net43 _01210_ _01694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08027__A1 _03296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07194_ _02643_ _02636_ _02644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09002_ _04068_ _04069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_54_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06145_ _01624_ _01625_ _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06589__A1 _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06076_ _01336_ _01532_ _01535_ _01451_ _01557_ _01558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_09904_ net80 _04869_ _04873_ _04874_ _04875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_111_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09835_ _04810_ _04811_ _02416_ _04819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09766_ _03207_ _04762_ _00500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06978_ _02035_ _02037_ _02450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_57_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05403__I3 cpu.regs\[11\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09697_ _04690_ _04691_ _04692_ _04706_ _04707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_08717_ _03840_ _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05929_ cpu.toggle_top\[9\] _01367_ _01409_ _01411_ _01175_ _01412_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_107_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08648_ cpu.pwm_counter\[4\] _03792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_1_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05390__I _00852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08579_ _03741_ cpu.toggle_top\[10\] cpu.toggle_top\[9\] _03742_ _03743_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10610_ _00504_ clknet_leaf_74_wb_clk_i cpu.ROM_spi_dat_out\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10541_ _00435_ clknet_leaf_55_wb_clk_i cpu.IO_addr_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09766__A1 _03207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10472_ _00367_ clknet_leaf_28_wb_clk_i cpu.timer_div_counter\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09518__A1 _04530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09037__I _04081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_2_0_wb_clk_i clknet_0_wb_clk_i clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_75_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_13_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07950_ cpu.spi.data_out_buff\[4\] _03218_ _03228_ _03241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06901_ _02375_ _01956_ _02073_ _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07881_ cpu.spi.div_counter\[4\] cpu.spi.divisor\[4\] _03179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09620_ cpu.PC\[11\] _01155_ _04612_ _04632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06832_ _02253_ _00877_ _00935_ _02293_ _02308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09551_ cpu.orig_PC\[9\] _04359_ _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06763_ _02196_ _02212_ _02239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05714_ _01051_ _01197_ _01198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08502_ _03675_ _03676_ _03667_ _00322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_54_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09482_ _02049_ _02050_ _02765_ _02057_ _04499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_06694_ _02168_ _02169_ _02170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_52_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08433_ cpu.orig_IO_addr_buff\[5\] _03627_ _03628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05645_ _01111_ _01128_ _01107_ _01001_ _01129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_08364_ _02821_ _03567_ _03573_ _03097_ _00287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_86_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05576_ _00673_ _01059_ _01060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_62_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09996__A1 net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07315_ _02742_ _02733_ _02743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08295_ cpu.uart.receive_counter\[0\] cpu.uart.receive_counter\[1\] cpu.uart.receive_counter\[3\]
+ cpu.uart.receive_counter\[2\] _03520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_116_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07246_ _02639_ _02689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07177_ _02629_ _00044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06128_ _01605_ _01607_ _01608_ _01609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__05085__I1 _00603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06059_ _01539_ _01540_ _01541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05785__A2 _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09818_ _02417_ _04769_ _04806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_94_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09749_ _04733_ _04731_ _04748_ _04749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xclkbuf_leaf_55_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_55_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_68_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08364__C _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput18 io_in[29] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_64_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput29 sram_out[3] net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10524_ _00419_ clknet_leaf_31_wb_clk_i cpu.timer_div\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10455_ _00350_ clknet_leaf_17_wb_clk_i cpu.pwm_counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09203__A3 _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10386_ _00281_ clknet_leaf_39_wb_clk_i cpu.uart.receive_div_counter\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05320__S1 _00827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05430_ _00853_ _00918_ _00919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_28_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05361_ _00850_ _00851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_16_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07100_ _02526_ _02563_ _02564_ _02565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08080_ cpu.uart.div_counter\[10\] _03344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_70_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06500__I1 _01976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05292_ _00786_ _00802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_113_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07031_ _02501_ _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08982_ cpu.uart.divisor\[14\] _04040_ _04049_ _04050_ _04051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07933_ cpu.spi.data_out_buff\[2\] _03212_ _03226_ _03227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09902__A1 _04031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07864_ _03160_ _03161_ _03162_ _03163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09603_ _04609_ _04615_ _00751_ _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06716__A1 _00900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06815_ _02243_ _00817_ _00877_ _00935_ _02291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_39_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07795_ _03100_ _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_104_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08469__A1 _02803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09534_ _04525_ _04549_ _04523_ _00481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06746_ _02219_ _02221_ _02222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09465_ _04456_ _04473_ _04482_ _04434_ _04483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06677_ cpu.regs\[1\]\[7\] _00876_ _01286_ _00789_ _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_19_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05628_ _00647_ _01032_ _01112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08416_ _01049_ _03610_ _03614_ _03613_ _00298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_59_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09969__A1 cpu.PORTA_DDR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09396_ _03649_ _04417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08347_ _03556_ _03559_ _03560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05559_ cpu.IO_addr_buff\[0\] _01043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08278_ _02646_ _03468_ _03507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_102_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_102_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07229_ _02655_ _02674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10240_ _00135_ clknet_leaf_102_wb_clk_i cpu.regs\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05758__A2 _01241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08944__A2 _00736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10171_ _00070_ clknet_leaf_12_wb_clk_i cpu.toggle_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_110_Right_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07683__A2 _03011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_7_Left_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10507_ _00402_ clknet_leaf_8_wb_clk_i cpu.timer_capture\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05297__I1 _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07199__A1 _02647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10438_ _00333_ clknet_leaf_7_wb_clk_i cpu.toggle_ctr\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10369_ _00264_ clknet_leaf_65_wb_clk_i cpu.uart.data_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_90_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05057__S0 _00572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06600_ _02073_ _02074_ _02076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07580_ cpu.regs\[10\]\[3\] _02946_ _02952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06531_ _01292_ _01957_ _02008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_0_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_0_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_34_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09250_ _01162_ _04273_ _04274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08201_ _03383_ _03443_ _03444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06462_ _01528_ _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06393_ _01378_ _01869_ _01870_ _01871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_90_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09181_ _04201_ _04208_ _04209_ _00468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05413_ _00902_ _00903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08132_ _03388_ _03389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05344_ cpu.PORTA_DDR\[7\] net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_71_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09828__C _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08063_ cpu.uart.div_counter\[15\] _03327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_70_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05275_ _00001_ _00786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07014_ _02447_ _02482_ _02485_ _02486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08965_ _00952_ _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_110_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07916_ _03211_ _03212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input24_I io_in[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08896_ _02624_ _03983_ _03986_ _00406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05663__I _00716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08179__C _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07847_ _03145_ cpu.timer\[11\] cpu.timer\[10\] _03142_ _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07778_ _02187_ _02329_ _02330_ _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_79_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06729_ _02201_ _02203_ _02204_ _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09517_ _04531_ _04532_ _04533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_65_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09448_ _04454_ _04466_ _04467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09379_ _04056_ _04385_ _04400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output92_I net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05838__I _01321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10223_ _00118_ clknet_leaf_125_wb_clk_i cpu.regs\[11\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_70_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_70_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10154_ _00053_ clknet_leaf_21_wb_clk_i cpu.timer_capture\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10085_ _01346_ _05025_ _05009_ _00847_ _01939_ _05026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_89_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08605__A1 _02882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05060_ _00580_ _00581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08750_ _03865_ _03866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05962_ _01442_ _01443_ _01445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05893_ _01092_ _01373_ _01375_ _01376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08681_ _03816_ _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_49_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07344__A1 _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07701_ _02983_ _03023_ _03026_ _00171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07632_ _02975_ _02980_ _02982_ _00146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07895__A2 cpu.spi.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09302_ _00725_ _00772_ _03624_ _04324_ _04325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07563_ _02940_ cpu.regs\[11\]\[5\] _02930_ _02941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06514_ _01196_ _01988_ _01989_ _01990_ _01991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__07203__I _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07494_ _02895_ _00095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09233_ _04214_ _04252_ _04258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06445_ _01919_ _01922_ _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_15_0_wb_clk_i clknet_0_wb_clk_i clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_90_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09164_ cpu.ROM_addr_buff\[7\] _04185_ _04198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08115_ _02621_ _03374_ _00236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06376_ _01424_ _01854_ _01855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09095_ _04144_ cpu.ROM_addr_buff\[5\] _04134_ _04145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05327_ cpu.regs\[12\]\[3\] cpu.regs\[13\]\[3\] cpu.regs\[14\]\[3\] cpu.regs\[15\]\[3\]
+ _00570_ _00827_ _00835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08046_ cpu.uart.dout\[4\] _03309_ _03314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05258_ cpu.instr_cycle\[1\] _00772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08969__I _04025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09021__A1 _01054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05189_ _00703_ _00704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05830__A1 _01155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09997_ _03822_ _04943_ _00550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08948_ _02537_ _04023_ _04024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05393__I _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08879_ _03973_ _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07335__A1 cpu.toggle_top\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_88_Left_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08835__A1 cpu.timer_capture\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07638__A2 _02980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05664__A4 _01008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_97_Left_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06074__B2 _01331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06074__A1 _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09484__B _04500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10206_ _00101_ clknet_leaf_2_wb_clk_i cpu.regs\[13\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05424__I1 cpu.regs\[1\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10137_ _00036_ clknet_leaf_105_wb_clk_i cpu.br_rel_dest\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10068_ _01262_ _04059_ _05008_ _05009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06230_ cpu.timer_capture\[12\] _01232_ _01238_ _01710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09659__B _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06161_ _01134_ _00841_ _01642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05112_ _00598_ _00630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06092_ _01321_ _01574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09920_ _04886_ _00530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09851_ _04827_ _03782_ _03786_ _04831_ _04832_ _04833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09782_ _04777_ _00501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06994_ _00691_ _02460_ _02465_ _02466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08802_ cpu.timer\[9\] _03909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08733_ cpu.timer_top\[13\] _03849_ _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06102__I _01583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05945_ _01161_ _00799_ _01428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05941__I _01148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08664_ cpu.pwm_top\[0\] _03801_ _03803_ _03697_ _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05876_ _01359_ _01360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08595_ cpu.toggle_ctr\[2\] _03754_ _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_07615_ _02922_ _02965_ _02970_ _00141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_62_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07546_ _02018_ _01131_ _02929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_118_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09216_ _02593_ _04240_ _04241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07477_ _01172_ _01145_ _02884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_107_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06428_ _01847_ _01897_ _01905_ _01906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_16_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09147_ _04170_ _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06359_ _01329_ _01837_ _01838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09078_ _04131_ cpu.ROM_addr_buff\[1\] _04023_ _04132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_31_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08029_ _03300_ _03301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_102_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06213__S _01207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output55_I net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07308__A1 cpu.toggle_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08808__A1 cpu.timer_capture\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06531__A2 _01957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07547__A1 _01158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07462__B _02871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05730_ _01092_ _01209_ _01212_ _01213_ _01214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_89_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_42_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07181__C _02518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05661_ _01010_ _01140_ _01144_ _01107_ _01145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_08380_ _03585_ _03581_ _03586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07400_ _02590_ _02811_ _02604_ _02813_ _00083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05592_ _01075_ _01056_ _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07331_ _02755_ _02747_ _02756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07262_ _02702_ _00056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06286__B2 _01322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06286__A1 _01435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10082__A2 _05017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06213_ cpu.PORTA_DDR\[4\] net55 _01207_ _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07193_ _02642_ _02643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09001_ _04055_ _04068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06144_ _01123_ _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06075_ _01296_ _01556_ _01557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05936__I _01340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09903_ _04861_ _04874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09834_ _04810_ _04816_ _02415_ _04818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_127_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_127_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_81_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09765_ cpu.spi_clkdiv _02479_ _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06977_ _02444_ _02038_ _02448_ _02449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_29_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09696_ _04147_ _04694_ _04703_ _04705_ _04706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_69_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08716_ _01090_ _02709_ _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_57_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05671__I _00930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05928_ _01410_ _01178_ _01367_ _01411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__06767__I _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08647_ _03789_ _03790_ _03791_ _00352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_1_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05859_ _01310_ _01343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_95_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08578_ _03704_ _03742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_37_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07529_ cpu.regs\[12\]\[1\] _02916_ _02919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10540_ _00434_ clknet_leaf_55_wb_clk_i cpu.IO_addr_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10471_ _00366_ clknet_leaf_28_wb_clk_i cpu.timer_div_counter\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07777__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05846__I _01329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_126_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10064__A2 _01290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06268__A1 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07301__I _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10669_ _00563_ clknet_leaf_123_wb_clk_i cpu.regs\[15\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07457__B _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_9_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07176__C _02518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09509__A2 _04379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06440__A1 _00654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06900_ _00634_ _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07880_ cpu.spi.div_counter\[0\] cpu.spi.divisor\[0\] _03178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06831_ _02289_ _02295_ _02307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05491__I _00977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09550_ _00752_ _04564_ _04565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06762_ _02226_ _02236_ _02237_ _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05713_ _01029_ _01084_ _01197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08501_ cpu.orig_PC\[13\] _03626_ _03676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_54_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09481_ _02558_ _02767_ _02560_ _04498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__09898__I _04868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08432_ _03626_ _03627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07299__A3 _02729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06693_ _02123_ _02124_ _02169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05644_ _01117_ _01124_ _01093_ _01127_ _01128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_19_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08363_ cpu.uart.receive_div_counter\[7\] _03542_ _03572_ _03573_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05575_ _01058_ _01030_ _01059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_46_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08294_ _03401_ _03519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_102_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07314_ _00952_ _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_62_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07245_ _02685_ _02686_ _02674_ _02687_ _02688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_6_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07176_ cpu.uart.divisor\[2\] _02613_ _02628_ _02518_ _02629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_42_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06127_ _01186_ _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_42_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08042__I _02872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05085__I2 _00604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06058_ _01151_ net92 _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05666__I _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09817_ _04771_ _04804_ _04805_ _00508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09748_ _02431_ _02433_ _04748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09679_ cpu.last_addr\[8\] _04679_ _04689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08487__A2 _03659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_68_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_95_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_95_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06498__A1 _01315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_24_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_24_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_65_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput19 io_in[2] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_91_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10523_ _00418_ clknet_leaf_30_wb_clk_i cpu.timer_div\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10454_ _00349_ clknet_leaf_17_wb_clk_i cpu.pwm_counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10385_ _00280_ clknet_leaf_39_wb_clk_i cpu.uart.receive_div_counter\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_70_Left_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_60_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05528__A3 _01010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06200__I _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08478__A2 _03659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06489__A1 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08127__I _03383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05360_ _00006_ _00850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XTAP_TAPCELL_ROW_31_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07031__I _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05291_ _00568_ _00801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07030_ _00683_ _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_70_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06661__A1 _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08981_ _04002_ _04050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07932_ _00926_ _03225_ _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07863_ _01864_ _02697_ _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09602_ _04392_ _04613_ _04614_ _04615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06814_ _02253_ _02157_ _02290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_39_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07794_ _03098_ _03099_ cpu.spi.counter\[4\] _03094_ _03100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_09533_ _04381_ _04544_ _04548_ _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_104_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06745_ _00602_ _02157_ _02221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09464_ _04477_ _04480_ _04481_ _04482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06676_ _02150_ _02151_ _02152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_19_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05152__A1 net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08415_ cpu.orig_IO_addr_buff\[1\] _03611_ _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09395_ _04381_ _04408_ _04415_ _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05627_ cpu.br_rel_dest\[0\] _01111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08346_ _02822_ _03548_ _03559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05558_ _00647_ _01041_ _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08277_ _03499_ _03504_ _03506_ _00267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_6_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05489_ _00975_ _00976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07228_ _02672_ _02673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_115_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07159_ _01419_ _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_14_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06404__A1 cpu.timer_capture\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10170_ _00069_ clknet_leaf_3_wb_clk_i cpu.toggle_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08157__A1 _03333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09657__A1 _02513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_69_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09331__I _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08880__A2 _02698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10506_ _00401_ clknet_leaf_8_wb_clk_i cpu.timer_capture\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05297__I2 _00806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10437_ _00332_ clknet_leaf_11_wb_clk_i cpu.toggle_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_78_Right_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10368_ _00263_ clknet_leaf_65_wb_clk_i cpu.uart.data_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_90_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10299_ _00194_ clknet_leaf_52_wb_clk_i cpu.spi.dout\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08410__I _03609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09506__I _00686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_108_Left_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09896__A1 _01046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05255__B _00735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05057__S1 _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09648__A1 _00763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_87_Right_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06530_ _01978_ _01784_ _02004_ _02006_ _02007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06461_ _01937_ _01938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_16_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08200_ cpu.uart.div_counter\[14\] _03439_ _03440_ _03443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_56_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05412_ _00901_ _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_8_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_117_Left_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06392_ net66 _01213_ _01870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09180_ cpu.last_addr\[12\] _04176_ _04209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08131_ _03387_ _03388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05343_ cpu.PORTB_DDR\[7\] net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_70_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09397__B _04417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08062_ _02859_ cpu.uart.div_counter\[15\] _03325_ _02630_ _03326_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_71_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06634__A1 _00831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05274_ _00000_ _00785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_96_Right_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07013_ cpu.ROM_addr_buff\[3\] _02483_ _02484_ cpu.ROM_addr_buff\[7\] _02452_ _02485_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_12_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10055__C _03366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08964_ _04036_ _00424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_110_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07915_ _03210_ _03211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08895_ cpu.spi.divisor\[1\] _03984_ _03986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07846_ cpu.timer_top\[11\] _03145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input17_I io_in[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07777_ _03082_ _03084_ _03085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06728_ _02199_ _02200_ _02204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09516_ _04524_ _00848_ _04532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_65_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09447_ _04347_ _04462_ _04465_ _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_109_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06659_ _02106_ _02107_ _02135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09378_ _02511_ _00735_ _04399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08329_ _02836_ _03537_ _03544_ _03545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08075__B1 _03335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09754__C _04721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10222_ _00117_ clknet_leaf_127_wb_clk_i cpu.regs\[11\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10153_ _00052_ clknet_leaf_22_wb_clk_i cpu.timer_capture\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09326__I _04277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09878__A1 net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10084_ _05017_ _05025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07728__I1 cpu.regs\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06864__A1 _00619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08605__A2 _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08369__A1 _02830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07041__A1 _00735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input9_I io_in[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09869__A1 _04031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05961_ _01442_ _01443_ _01444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07700_ cpu.regs\[4\]\[1\] _03024_ _03026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05892_ cpu.PORTB_DDR\[1\] _01374_ _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08680_ cpu.pwm_top\[4\] _03814_ _03815_ _03809_ _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_49_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07631_ cpu.regs\[7\]\[0\] _02981_ _02982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07562_ _01857_ _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06513_ cpu.uart.divisor\[15\] _01489_ _00012_ _01990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_76_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09301_ _00724_ _04323_ _04324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07493_ _01858_ cpu.regs\[14\]\[5\] _02886_ _02895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09232_ _00902_ _04019_ _04062_ _04256_ _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06444_ _01439_ _01897_ _01921_ _01453_ _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_35_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09163_ cpu.last_addr\[7\] _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_16_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06375_ net95 _01297_ _01853_ _01854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_114_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08114_ _03099_ _03367_ _03373_ _03371_ _03374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_90_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05326_ _00828_ _00833_ _00581_ _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09094_ _00604_ _02550_ _04130_ _04144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_9_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08045_ cpu.uart.receive_buff\[4\] _03307_ _03313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05257_ _00741_ _00752_ _00759_ _00770_ _00771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_112_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05188_ _00702_ _00703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09996_ net75 _04938_ _04942_ _04759_ _04943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_86_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08947_ _04022_ _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08878_ cpu.timer_capture\[13\] _03965_ _03972_ _03968_ _03973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_99_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07829_ _03122_ cpu.timer_div_counter\[2\] _03127_ cpu.timer_div\[6\] _03128_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08532__A1 cpu.toggle_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07099__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06454__B _01478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07023__A1 _00693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10205_ _00100_ clknet_leaf_2_wb_clk_i cpu.regs\[13\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10136_ _00035_ clknet_leaf_105_wb_clk_i cpu.br_rel_dest\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_89_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10067_ _05003_ _05007_ _00748_ _05008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_32_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06160_ _01586_ _00840_ _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05111_ _00629_ net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_06091_ _01549_ _01572_ _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_71_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09850_ cpu.pwm_top\[6\] cpu.pwm_counter\[6\] _04832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09781_ cpu.ROM_spi_dat_out\[0\] _04771_ _04776_ _04721_ _04777_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06993_ _02461_ _02464_ _02465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08801_ _03907_ _03908_ _00389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08732_ _02635_ _03848_ _03850_ _03851_ _00377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05944_ _01363_ _00814_ _01427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08663_ _02615_ _03802_ _03803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05875_ _01358_ _01359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_88_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08594_ _03749_ _03756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07614_ cpu.regs\[8\]\[3\] _02964_ _02970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_62_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07545_ _02927_ _02916_ _02928_ _00113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07476_ _02883_ _00089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10085__B1 _05009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08293__A3 _03518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09215_ _02796_ _04240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06427_ _01847_ _01904_ _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09146_ cpu.last_addr\[3\] _04184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__09242__A2 _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06358_ _01825_ _01686_ _01837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09077_ _00806_ _02783_ _04130_ _04131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06289_ net30 _01425_ _01478_ _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05309_ cpu.regs\[2\]\[2\] _00818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_32_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08028_ _02877_ _02878_ _03300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_49_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_49_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_4_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09979_ _02642_ _04927_ _04930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_105_Right_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_95_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_116_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07244__A1 _00967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10119_ _00018_ clknet_leaf_124_wb_clk_i cpu.regs\[9\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05660_ _01141_ _01143_ _01144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05730__A1 _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05591_ _01074_ _00679_ _01075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07330_ _02698_ _02755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10538__CLK clknet_leaf_18_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07261_ cpu.timer_capture\[6\] _02684_ _02701_ _02689_ _02702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09000_ _04066_ _04067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06212_ cpu.uart.divisor\[4\] _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_98_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07192_ _01688_ _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06143_ cpu.toggle_top\[11\] _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06589__A3 _02064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06074_ _00924_ _01339_ _01534_ _01331_ _01556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09902_ _04031_ _04870_ _04873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09833_ _03207_ _04817_ _00512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07209__I _02655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10063__C _04213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09764_ _04761_ _00499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06976_ _02025_ _02030_ _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_29_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08715_ _03827_ _03839_ _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09695_ cpu.last_addr\[5\] cpu.ROM_addr_buff\[5\] _04704_ _04705_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_57_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05927_ cpu.toggle_top\[1\] _01410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_107_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09160__A1 _04147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08646_ cpu.pwm_counter\[3\] _03788_ _03791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_1_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05858_ _01333_ _01336_ _01339_ _01340_ _01341_ _01342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_64_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05789_ _01110_ _01072_ _01272_ _01021_ _01273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_37_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08577_ cpu.toggle_ctr\[10\] _03741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_49_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07528_ _01481_ _02918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07459_ cpu.uart.receive_counter\[1\] _02865_ _02866_ _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_91_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10470_ _00365_ clknet_leaf_33_wb_clk_i cpu.timer_div_counter\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09129_ _02471_ _04169_ _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08726__A1 cpu.timer_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06201__A2 _01681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09151__A1 cpu.ROM_addr_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10668_ _00562_ clknet_leaf_123_wb_clk_i cpu.regs\[15\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10599_ _00493_ clknet_leaf_73_wb_clk_i cpu.startup_cycle\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__08413__I _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06361__C _00716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06830_ _02288_ _02296_ _02302_ _02306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_06761_ _02234_ _02235_ _02237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05712_ _01195_ _01196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09142__A1 _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08500_ _03674_ _03611_ _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09480_ _04496_ _04497_ _04417_ _00479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_54_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06692_ _02165_ _02166_ _02167_ _02168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08431_ _03625_ _03626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05643_ _01125_ _01126_ _01127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08362_ _03570_ _03571_ _03572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05574_ cpu.IO_addr_buff\[3\] _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_58_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08293_ _03514_ _02881_ _03518_ _00271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_102_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07313_ _02741_ _00068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07244_ _00967_ _02680_ _02687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07175_ _02627_ _02616_ _02628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06126_ cpu.spi.divisor\[3\] _01606_ _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05085__I3 cpu.regs\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06431__A2 _00999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06057_ _01152_ _01530_ _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_70_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09816_ cpu.ROM_spi_dat_out\[7\] _04772_ _02715_ _04805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06959_ cpu.startup_cycle\[3\] _02431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09747_ _04222_ _04747_ _00496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09678_ _04204_ cpu.ROM_addr_buff\[10\] _04680_ _04688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_68_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08629_ cpu.toggle_ctr\[14\] _03778_ _03779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_81_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_64_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_64_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10522_ _00417_ clknet_leaf_30_wb_clk_i cpu.timer_div\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05857__I _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10453_ _00348_ clknet_leaf_5_wb_clk_i cpu.toggle_ctr\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10384_ _00279_ clknet_leaf_43_wb_clk_i cpu.uart.receive_buff\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07513__S _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05290_ _00800_ net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08143__I _03383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07610__A1 cpu.regs\[8\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08980_ _04048_ _04042_ _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07931_ _03213_ _03225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07862_ _01864_ cpu.timer\[6\] cpu.timer\[5\] _01786_ _03161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_09601_ _04392_ _04602_ _04396_ _04614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06813_ _02267_ _02268_ _02289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_39_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07793_ cpu.spi.counter\[2\] _03099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09532_ _04443_ _04527_ _04546_ _04547_ _04414_ _04548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_104_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06744_ _00901_ _02219_ _02220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09463_ _04477_ _04480_ _04273_ _04481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_19_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06675_ _00789_ _00875_ _02151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08414_ _01055_ _03610_ _03612_ _03613_ _00297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_59_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05626_ _01017_ _01110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09394_ _02513_ _04386_ _04412_ _04413_ _04414_ _04415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08345_ _03544_ _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_80_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05557_ _01040_ _01041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07222__I _00909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08276_ cpu.uart.data_buff\[7\] _03497_ _03505_ _03506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05488_ _00974_ _00975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07227_ cpu.timer\[2\] _02672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07158_ _02612_ _02613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05677__I _01111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06109_ cpu.toggle_top\[3\] _01590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__10235__D _00130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08988__I _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07089_ _02370_ _02554_ _02544_ _02555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_100_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_4_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_111_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_111_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07904__A2 _03195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05915__A1 cpu.timer_div\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10505_ _00400_ clknet_leaf_9_wb_clk_i cpu.timer_capture\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05297__I3 cpu.regs\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10436_ _00331_ clknet_leaf_10_wb_clk_i cpu.toggle_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10367_ _00262_ clknet_leaf_63_wb_clk_i cpu.uart.data_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05454__I0 cpu.regs\[8\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10298_ _00193_ clknet_leaf_42_wb_clk_i cpu.spi.dout\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07307__I _02639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05382__A2 _00869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06460_ _00642_ _01937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05411_ _00900_ _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_16_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08130_ _03364_ _03386_ _03387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06391_ _01374_ _01867_ _01868_ _01121_ _01869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_71_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05342_ cpu.PORTA_DDR\[6\] net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_16_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08061_ cpu.uart.div_counter\[3\] _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_70_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06634__A2 _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05273_ _00784_ cpu.ROM_spi_mode net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_113_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07012_ _02454_ _02484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08963_ _02828_ _04026_ _04034_ _04035_ _04036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07914_ _00722_ _03209_ _00756_ _01066_ _03210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_110_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08894_ _02708_ _03983_ _03985_ _00405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07217__I _02639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07845_ _03142_ _03143_ cpu.timer\[9\] _03139_ _03144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_79_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07776_ _03083_ _03071_ _03084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09515_ _02048_ _01344_ _04531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06727_ _02190_ _02202_ _02203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_65_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09446_ _01774_ _04430_ _04464_ _04355_ _04465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06658_ _02128_ _02133_ _02134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05609_ _01089_ _01092_ _01093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09377_ _04392_ _04395_ _04397_ _04398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06589_ _00949_ _02063_ _02064_ _02065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_117_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08328_ _03538_ _03544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_105_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08259_ _00926_ _03486_ _03492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06625__A2 _01955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10221_ _00116_ clknet_leaf_127_wb_clk_i cpu.regs\[11\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output78_I net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10152_ _00051_ clknet_leaf_22_wb_clk_i cpu.timer_capture\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10083_ _01468_ _05016_ _05023_ _05024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06313__A1 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08066__A1 cpu.uart.divisor\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06206__I _01685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05110__I _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10419_ _00314_ clknet_leaf_90_wb_clk_i cpu.orig_PC\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_61_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05960_ _01430_ _01443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05891_ _01210_ _01374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_49_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07630_ _02978_ _02981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08541__A2 _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07561_ _02939_ _00118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06512_ cpu.uart.divisor\[7\] _01502_ _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09300_ _04300_ _04302_ _04322_ _04291_ _04323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_07492_ _02894_ _00094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09231_ cpu.orig_flags\[1\] _04239_ _04255_ _04256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06443_ _00629_ _01920_ _01921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_90_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09162_ _04187_ _04195_ _04196_ _00462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06374_ _01822_ _01824_ _01845_ _01852_ _01853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_08113_ _03099_ _03370_ _03373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_83_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07500__I _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05325_ cpu.regs\[0\]\[3\] _00831_ _00832_ cpu.regs\[3\]\[3\] _00570_ _00827_ _00833_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09093_ _04143_ _00446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08044_ _03308_ _03310_ _03312_ _00228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05256_ _00763_ _00767_ _00769_ _00770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_31_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05187_ _00701_ _00702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_4_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09995_ _02422_ _02428_ _02437_ _04939_ _04941_ _04942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_08946_ _02638_ _00733_ _04021_ _04022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__06791__A1 _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08877_ _03944_ _03971_ _03972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07828_ cpu.timer_div_counter\[6\] _03127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_79_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05690__I _01100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07759_ _03068_ _00187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07099__A2 _02361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09429_ _02550_ _04379_ _04448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09548__A1 _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10204_ _00099_ clknet_leaf_2_wb_clk_i cpu.regs\[13\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05424__I3 cpu.regs\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10135_ _00034_ clknet_leaf_105_wb_clk_i cpu.br_rel_dest\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_89_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10066_ _01003_ _04213_ _05006_ _05007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_82_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07582__I0 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06534__A1 _01133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10011__I net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10094__A1 _02885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09236__B1 _01290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07320__I _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05110_ _00628_ _00629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_41_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06090_ _01550_ _01571_ _01572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08800_ cpu.timer_capture\[8\] _03888_ _03889_ _03908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09780_ _04772_ _04775_ _04776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06992_ _02032_ _02462_ _02036_ _02463_ _02464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06773__A1 _00899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08731_ _02723_ _03851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05943_ _01306_ _01426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08662_ _03800_ _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06525__A1 cpu.toggle_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07613_ _02920_ _02965_ _02969_ _00140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05874_ _01167_ _01295_ _01356_ _01357_ _01358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_08593_ _03753_ _03754_ _03755_ _00334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_49_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08278__A1 _02646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07544_ cpu.regs\[12\]\[7\] _02914_ _02928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07475_ _02879_ _02881_ _02882_ _02883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10085__B2 _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09214_ _04060_ _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06426_ _01901_ _01903_ _01904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_118_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08326__I _03517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07230__I _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09145_ _03378_ _04182_ _04183_ _00458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08770__B _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06357_ _01826_ _01746_ _01836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09076_ _00727_ _04130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_71_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09585__C _04081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05308_ _00816_ _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06288_ _01012_ _01767_ _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_114_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08027_ _03296_ _03299_ _00224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05239_ _00711_ _00656_ _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_31_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_73_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09950__A1 cpu.PORTB_DDR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09978_ _04929_ _00545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_89_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_89_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_99_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08929_ _03995_ _04009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_18_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_18_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_99_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08505__A2 _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07140__I _02598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05255__A1 _00734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10118_ _00017_ clknet_leaf_123_wb_clk_i cpu.regs\[9\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05802__I0 _01281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10049_ _00663_ _04990_ _04991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06507__A1 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07180__A1 _02631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_11_Left_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05590_ _00671_ _01074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06375__B _01853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07260_ _02660_ _02700_ _02701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06211_ cpu.spi.dout\[4\] _01691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07191_ _02641_ _00046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_54_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06142_ _01590_ _01177_ _01620_ _01622_ _01254_ _01623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_41_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06073_ _01548_ _01553_ _01554_ _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09901_ _04872_ _00525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_111_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09832_ _04810_ _04816_ _04817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_6_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09763_ _04732_ _04757_ _04758_ _04760_ _03474_ _04761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06975_ _02442_ _02445_ _02446_ _02447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08714_ cpu.timer_div_counter\[7\] _03838_ _03839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_4_9_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09694_ _04189_ _04677_ _04704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05926_ _01405_ _01406_ _01407_ _01408_ _01409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xrebuffer10 net123 net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_107_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07171__A1 _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08645_ cpu.pwm_counter\[3\] _03788_ _03790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_1_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05857_ _01147_ _01341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08765__B _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08576_ _03739_ _01256_ _03718_ _03720_ _03740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08484__C _03653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05788_ _00703_ _01099_ _01272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07527_ _02910_ _02915_ _02917_ _00106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_37_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07458_ cpu.uart.receive_counter\[0\] cpu.uart.receive_counter\[1\] _02864_ _02868_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__08056__I _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06409_ cpu.toggle_top\[6\] _01177_ _01887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07389_ _02803_ _02804_ _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09128_ _00666_ _04168_ _04169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_118_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09059_ _01002_ _04115_ _04117_ _04050_ _04118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_9_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07135__I _02514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07162__A1 _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10162__CLK clknet_leaf_18_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10667_ _00561_ clknet_leaf_0_wb_clk_i cpu.regs\[15\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08414__A1 _01055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10598_ _00492_ clknet_leaf_70_wb_clk_i cpu.mem_cycle\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05228__A1 cpu.uart.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09914__A1 _04041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput90 net90 sram_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05087__S0 _00572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06760_ _02234_ _02235_ _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05711_ _01036_ _01052_ _01119_ _01195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_06691_ _02163_ _02164_ _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_77_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08430_ _03624_ _03606_ _03625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05642_ _01083_ _01120_ _01126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08361_ _02821_ _03567_ _03571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_05573_ _01056_ _01057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_34_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08292_ _03517_ _03518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_102_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08653__A1 _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07312_ cpu.toggle_top\[10\] _02732_ _02740_ _02737_ _02741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_6_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07929__B _03112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07243_ _02658_ _02686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_33_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07174_ _00925_ _02627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06125_ _01076_ _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05314__S1 _00574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06056_ _01535_ _01537_ _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09815_ cpu.ROM_spi_dat_out\[6\] _04790_ _04792_ _04804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09746_ _02432_ _04745_ _04747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06958_ _02421_ cpu.startup_cycle\[5\] _02430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09677_ cpu.last_addr\[11\] cpu.ROM_addr_buff\[11\] _04681_ _04687_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_05909_ cpu.spi.dout\[1\] _01392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_96_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06889_ _02364_ _00021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06794__I _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08628_ _03750_ _03777_ _03778_ _00346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_84_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08559_ _03722_ _03723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_92_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10521_ _00416_ clknet_leaf_30_wb_clk_i cpu.timer_div\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_9_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10452_ _00347_ clknet_leaf_5_wb_clk_i cpu.toggle_ctr\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10383_ _00278_ clknet_leaf_43_wb_clk_i cpu.uart.receive_buff\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_33_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_33_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_92_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07758__I0 _00806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07293__C _02724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05697__A1 _01094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08883__A1 cpu.timer_capture\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05113__I _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08424__I _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer1 _02331_ net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07930_ _03220_ _03222_ _03224_ _00202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05621__A1 _01081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07861_ _01786_ cpu.timer\[5\] cpu.timer\[4\] _01689_ _03159_ _03160_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_07792_ cpu.spi.counter\[3\] _03098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09600_ _03081_ _00932_ _04612_ _04613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06812_ _02277_ _02273_ _02278_ _02288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XTAP_TAPCELL_ROW_39_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09531_ _04373_ _04547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06743_ _02217_ _02218_ _02219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_104_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09462_ _04478_ _04479_ _04480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06674_ cpu.regs\[1\]\[7\] _01286_ _02150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_19_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08413_ _02602_ _03613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09393_ _04226_ _04414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05625_ _00740_ _01014_ _01108_ _01109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_08344_ _03517_ _03557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05556_ cpu.IO_addr_buff\[3\] cpu.IO_addr_buff\[2\] _01040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_19_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09858__C _03288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08275_ _00776_ _03505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05958__I _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05487_ _00973_ _00974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07226_ _02671_ _00051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07157_ _01198_ _02611_ _02612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__09051__A1 _01133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_1_0_wb_clk_i clknet_0_wb_clk_i clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_06108_ _01276_ _01589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07088_ _02365_ _02553_ _02542_ _02554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06039_ _01520_ _01257_ _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_12_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09729_ cpu.startup_cycle\[1\] _04733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__09106__A2 cpu.regs\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05471__S0 _00956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08865__A1 _00978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10504_ _00399_ clknet_leaf_9_wb_clk_i cpu.timer_capture\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09042__A1 _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10435_ _00330_ clknet_leaf_11_wb_clk_i cpu.toggle_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10366_ _00261_ clknet_leaf_64_wb_clk_i cpu.uart.data_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_51_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10297_ _00192_ clknet_leaf_42_wb_clk_i cpu.spi.dout\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07108__A1 _02570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07659__A2 _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05410_ _00899_ _00900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06390_ net46 _01211_ _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05341_ cpu.PORTB_DDR\[6\] net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_70_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_90_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09281__A1 _00762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08060_ _02843_ _03323_ cpu.uart.div_counter\[8\] _02831_ _03324_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_05272_ net75 _00784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07011_ _02449_ _02483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_113_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07993__I _03275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08962_ _04002_ _04035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08893_ cpu.spi.divisor\[0\] _03984_ _03985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07913_ _00679_ _03209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_110_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07844_ cpu.timer\[10\] _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07898__A2 _03195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_3_Left_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07775_ _03070_ _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09514_ _04504_ _04528_ _04529_ _04530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06726_ _02188_ _02189_ _02202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09445_ _04350_ _04451_ _04463_ _04353_ _04464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06657_ _02129_ _02132_ _02133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05608_ _01091_ _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_74_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09376_ _04392_ _04385_ _04396_ _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06588_ _00633_ _00935_ _02064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08327_ _03542_ _03540_ _03543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05539_ _00702_ _01017_ _01022_ _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_47_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08258_ _03464_ _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Left_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_105_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07209_ _02655_ _02656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09024__A1 _01153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05833__A1 _01315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08189_ cpu.uart.div_counter\[11\] _03428_ _03434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_42_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10220_ _00115_ clknet_leaf_127_wb_clk_i cpu.regs\[11\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_76_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10151_ _00050_ clknet_leaf_22_wb_clk_i cpu.timer_capture\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10082_ _01655_ _05017_ _05022_ _05023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_58_Left_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_67_Left_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09263__A1 _01298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10418_ _00313_ clknet_leaf_86_wb_clk_i cpu.orig_PC\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10349_ _00244_ clknet_leaf_33_wb_clk_i cpu.uart.div_counter\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_76_Left_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07318__I _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05890_ cpu.PORTA_DDR\[1\] net80 _01208_ _01373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_49_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08829__A1 cpu.timer_capture\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07560_ _02938_ cpu.regs\[11\]\[4\] _02931_ _02939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06378__B _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06511_ net14 _01372_ _01383_ _01987_ _01988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_88_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09230_ _04245_ _04250_ _04253_ _04254_ _04255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_07491_ _01772_ cpu.regs\[14\]\[4\] _02887_ _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06442_ _00613_ _01746_ _01920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09161_ cpu.last_addr\[6\] _04192_ _04196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09254__A1 cpu.PC\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06373_ _01435_ _01850_ _01851_ _01852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_16_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08112_ _03366_ _03369_ _03372_ _00235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09092_ _04142_ cpu.ROM_addr_buff\[4\] _04134_ _04143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06068__A1 _01364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05324_ cpu.regs\[2\]\[3\] _00832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_114_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08043_ _03311_ _03312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05815__A1 _01298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05255_ _00734_ _00768_ _00735_ _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05186_ cpu.br_rel_dest\[5\] _00701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_110_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09994_ _02450_ _04940_ _02458_ _04941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_50_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06240__A1 _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08945_ _00730_ _04020_ _04021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input22_I io_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08876_ _03929_ _03946_ _03970_ _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05971__I _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07827_ cpu.timer_div\[1\] _03119_ _03120_ cpu.timer_div\[5\] _03125_ _03126_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__05426__S0 _00856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07758_ _00806_ _03067_ _03058_ _03068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_66_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06709_ _02162_ _02184_ _02182_ _02185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07689_ _03018_ _00167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09428_ _04419_ _04447_ _04417_ _00477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_109_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09359_ _02052_ _04379_ _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output90_I net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08522__I _03678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10203_ _00098_ clknet_leaf_3_wb_clk_i cpu.regs\[13\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10134_ _00033_ clknet_leaf_102_wb_clk_i cpu.regs\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09781__C _04721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09353__I _04226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10065_ _01419_ _01272_ _05005_ _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_46_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08432__I _03626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05273__A2 cpu.ROM_spi_mode vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_84_Left_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06991_ _02037_ _02463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08730_ cpu.timer_top\[12\] _03849_ _03850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05942_ _01424_ _01425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08661_ _03800_ _03801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05873_ _01150_ _01357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_07612_ cpu.regs\[8\]\[2\] _02966_ _02969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07722__A1 cpu.regs\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_93_Left_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08592_ _03677_ cpu.toggle_ctr\[0\] cpu.toggle_ctr\[1\] _03755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_76_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07543_ _02014_ _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07474_ _02517_ _02882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_62_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06289__A1 net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09213_ _02614_ _01268_ _01863_ _04237_ _04238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__09227__A1 _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06425_ _01837_ _01902_ _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_17_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09144_ cpu.last_addr\[2\] _04177_ _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09078__I1 cpu.ROM_addr_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07089__I0 _02370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06356_ _01825_ _01834_ _01835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_16_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09075_ _04129_ _00442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05307_ cpu.regs\[1\]\[2\] _00816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06287_ _01724_ _01529_ _01752_ _01766_ _01767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_31_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08026_ cpu.spi.data_in_buff\[6\] _03198_ _03294_ cpu.spi.data_in_buff\[7\] _03299_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05238_ _00751_ _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05169_ _00684_ _00685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_73_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09977_ cpu.PORTA_DDR\[4\] _04926_ _04928_ _04920_ _04929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08928_ _04008_ _00416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_99_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08859_ cpu.timer_capture\[9\] _03943_ _03957_ _03951_ _03958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xclkbuf_leaf_58_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_58_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_95_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10076__A2 _01291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05327__I0 cpu.regs\[12\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09218__A1 _01153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05255__A2 _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09348__I _04319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06452__A1 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05876__I _01359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06204__A1 _00982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_14_0_wb_clk_i clknet_0_wb_clk_i clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_10117_ _00016_ clknet_leaf_1_wb_clk_i cpu.regs\[9\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10048_ _02440_ _04989_ _04990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10022__I net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06210_ _01181_ _01690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09209__B2 _01976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07190_ cpu.uart.divisor\[4\] _02613_ _02637_ _02640_ _02641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_54_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06141_ cpu.pwm_top\[3\] _01621_ _01177_ _01622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06072_ _01549_ _01552_ _01554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09900_ net79 _04869_ _04871_ _04862_ _04872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_111_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09831_ _03288_ _04815_ _04816_ _00511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__10584__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09762_ _04732_ _04759_ _04760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06974_ _02035_ _02037_ _02446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08713_ cpu.timer_div_counter\[6\] _03834_ _03838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05925_ _01125_ _01408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09693_ cpu.ROM_addr_buff\[6\] _04694_ _04695_ _04702_ _04703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09696__A1 _04147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer11 _00955_ net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_107_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08644_ _02812_ _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05856_ _01309_ _01340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_95_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05787_ _01270_ _01271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08575_ cpu.toggle_ctr\[8\] _03739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_1_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08337__I _02872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07526_ cpu.regs\[12\]\[0\] _02916_ _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_37_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07241__I _02655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07457_ _02865_ _02867_ _00739_ _00086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_64_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06408_ cpu.pwm_top\[6\] _01619_ _01408_ _01886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05485__A2 _00943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07388_ _02788_ _02782_ _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09127_ cpu.mem_cycle\[1\] _02029_ _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_72_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06339_ _00612_ _01685_ _01818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_105_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_105_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_118_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09058_ _02499_ _04116_ _04117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_118_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08009_ _03285_ _03199_ _03287_ _03093_ _03288_ _00217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_4_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_9_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05645__B _01107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output53_I net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10666_ _00560_ clknet_leaf_0_wb_clk_i cpu.regs\[15\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_97_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10597_ _00491_ clknet_leaf_69_wb_clk_i cpu.mem_cycle\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05228__A2 cpu.spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput80 net80 io_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput91 net91 sram_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05087__S1 _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07326__I _02638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_qcpu_98 io_oeb[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_37_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05710_ _01193_ _01194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_53_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06690_ cpu.regs\[1\]\[0\] _01954_ _02166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05641_ _01112_ _01083_ _01125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08360_ _03539_ _03570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06361__B1 _01839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05572_ _01054_ _01055_ _01056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07311_ _02739_ _02733_ _02740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_34_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_3_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_3_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08291_ _03516_ _03517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_102_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07242_ cpu.timer\[4\] _02685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_61_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07173_ _02621_ _02626_ _00043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06124_ cpu.uart.dout\[3\] _01194_ _01602_ _01604_ _01080_ _01605_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_42_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06416__A1 _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06055_ _01458_ _01536_ _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09814_ _04803_ _00507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_6_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09745_ _02438_ _04744_ _04746_ _00495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06957_ _02425_ _02428_ _00665_ _02429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09676_ cpu.last_addr\[12\] cpu.ROM_addr_buff\[12\] _04685_ _04686_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_05908_ _01390_ cpu.spi.divisor\[1\] _01189_ _01391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06888_ _00591_ _02358_ _02363_ _02364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05839_ cpu.C _01302_ _01304_ _01323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08627_ cpu.toggle_ctr\[13\] _03776_ _03778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_77_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08558_ cpu.toggle_ctr\[6\] _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08489_ _03665_ _03666_ _03667_ _00318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_65_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07509_ cpu.regs\[13\]\[3\] _02899_ _02905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10520_ _00415_ clknet_leaf_21_wb_clk_i cpu.timer_div\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_30_Left_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10451_ _00346_ clknet_leaf_4_wb_clk_i cpu.toggle_ctr\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10382_ _00277_ clknet_leaf_39_wb_clk_i cpu.uart.receive_buff\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_41_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07080__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_73_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_73_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_59_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_80_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06646__A1 cpu.regs\[1\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10649_ _00543_ clknet_leaf_59_wb_clk_i cpu.PORTA_DDR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_3_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer2 net119 net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_113_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08440__I _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09899__A1 _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07860_ cpu.timer_top\[4\] _02685_ _02679_ cpu.timer_top\[3\] _03158_ _03159_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09363__A3 cpu.PC\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07791_ _03093_ _03095_ _03096_ _03097_ _00190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06811_ _02286_ _02275_ _02287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_64_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09530_ _00790_ _04409_ _04545_ _04546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06895__I _00603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06742_ _00829_ _00933_ _02218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_39_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09461_ cpu.PC\[6\] _01019_ _04479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_104_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06673_ _02120_ _02148_ _02149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08412_ cpu.orig_IO_addr_buff\[0\] _03611_ _03612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09392_ _04373_ _04413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_19_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05624_ _01015_ _01106_ _01107_ _00844_ _01108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_08343_ cpu.uart.receive_div_counter\[4\] _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05152__A4 _00668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05555_ cpu.IO_addr_buff\[4\] _01039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08274_ cpu.uart.data_buff\[6\] _03491_ _03503_ _03504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06637__A1 _00634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07225_ cpu.timer_capture\[1\] _02656_ _02670_ _02664_ _02671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_61_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05486_ _00948_ _00972_ _00973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_27_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10085__C _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07156_ _02610_ _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_15_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06107_ _01587_ _01165_ _01166_ _01588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__07062__A1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07087_ _02546_ _02548_ _02551_ _02552_ _02553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06038_ cpu.toggle_top\[10\] _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_100_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_125_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09728_ cpu.startup_cycle\[6\] _04732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07989_ cpu.spi.div_counter\[5\] _03272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05471__S1 _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09659_ _04647_ _04669_ _00687_ _00486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_8_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05214__I _00668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_120_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_120_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_37_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_108_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10503_ _00398_ clknet_leaf_9_wb_clk_i cpu.timer_capture\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10434_ _00329_ clknet_leaf_11_wb_clk_i cpu.toggle_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10365_ _00260_ clknet_leaf_64_wb_clk_i cpu.uart.counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10296_ _00191_ clknet_leaf_52_wb_clk_i cpu.spi.dout\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05340_ cpu.PORTA_DDR\[5\] net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06619__A1 _02093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05271_ _00687_ _00783_ _00009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_113_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07010_ cpu.ROM_addr_buff\[11\] _02459_ _02455_ _02482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_3_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08961_ _02739_ _04028_ _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07912_ _03207_ _03095_ _03208_ _00200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08892_ _03982_ _03984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_110_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07843_ cpu.timer_top\[10\] _03142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05743__B _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07774_ _03081_ _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_79_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09513_ _02049_ _01018_ _04529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06725_ _02199_ _02200_ _02201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10103__A1 _01583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09444_ _02549_ _04351_ _04463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06656_ _02130_ _02131_ _02132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05607_ _01087_ _01090_ _01091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_74_Right_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09375_ _00766_ _04396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06587_ _00817_ _01287_ _02063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08326_ _03517_ _03542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05538_ _01018_ _01020_ _01021_ _01022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_7_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08257_ _03481_ _03488_ _03490_ _00263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_104_Left_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07283__A1 _02631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05469_ _00955_ _00956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_08188_ _03427_ _03433_ _00251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07208_ _01057_ _01078_ _01234_ _02610_ _02655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_62_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07139_ _02536_ _02540_ _02597_ _02493_ _02598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__07035__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_83_Right_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_76_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10150_ _00049_ clknet_leaf_31_wb_clk_i cpu.uart.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10081_ _01734_ _05012_ _05019_ _05021_ _05022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08535__A1 cpu.toggle_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_113_Left_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_92_Right_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09263__A2 _01002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10417_ _00312_ clknet_leaf_90_wb_clk_i cpu.orig_PC\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05828__B _01262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10348_ _00243_ clknet_leaf_33_wb_clk_i cpu.uart.div_counter\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10279_ _00174_ clknet_leaf_114_wb_clk_i cpu.regs\[4\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05563__B _01046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05760__A1 cpu.timer_capture\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06510_ _01982_ _01035_ _01985_ _01986_ _01204_ _01987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_48_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07490_ _01680_ _02888_ _02893_ _00093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06441_ _01331_ _01898_ _01916_ _01450_ _01918_ _01919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_118_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_100_Right_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_75_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09160_ _04147_ _04194_ _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06372_ _01846_ _01849_ _01851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_16_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08111_ _03094_ _03370_ _03371_ _03372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07265__A1 _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09091_ _02051_ _04136_ _04141_ _04142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05323_ _00830_ _00831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06068__A2 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08042_ _02872_ _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05254_ _00684_ _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05815__A2 _00712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05371__S0 _00856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05185_ _00687_ _00700_ _00011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09993_ _02031_ _02462_ _04940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08944_ _00754_ _00736_ _00746_ _04019_ _04020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_08875_ _02692_ _03947_ _03970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07826_ cpu.timer_div\[5\] _03120_ cpu.timer_div_counter\[7\] _01995_ _03124_ _03125_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__05426__S1 _00860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input15_I io_in[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07757_ _01480_ _02407_ _03066_ _03067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_94_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06708_ _02182_ _02183_ _02184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09493__A2 _04484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07688_ _03004_ cpu.regs\[5\]\[5\] _03009_ _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_94_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09427_ _04381_ _04442_ _04446_ _04447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06639_ _02065_ _02114_ _02115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09358_ _04296_ _04379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08309_ cpu.uart.receive_buff\[3\] _03523_ _03530_ cpu.uart.receive_buff\[4\] _03531_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09289_ _04309_ _04311_ _04312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_50_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05114__S0 _00630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10202_ _00097_ clknet_leaf_120_wb_clk_i cpu.regs\[14\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10133_ _00032_ clknet_leaf_101_wb_clk_i cpu.regs\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_89_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10064_ _04259_ _01290_ _05004_ _05005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05990__B2 _01322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07154__I _01008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07247__A1 cpu.timer_capture\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06990_ _02443_ _02462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input7_I io_in[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05941_ _01148_ _01424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08660_ _01067_ _02730_ _03800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05872_ _01012_ _01354_ _01355_ _01356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_07611_ _02918_ _02965_ _02968_ _00139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05733__A1 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08591_ cpu.toggle_clkdiv cpu.toggle_ctr\[1\] cpu.toggle_ctr\[0\] _03754_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_88_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07542_ _02926_ _00112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07473_ _02880_ _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09212_ _00909_ _00937_ _04236_ _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_06424_ _01825_ _01686_ _01828_ _01902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09143_ cpu.ROM_addr_buff\[2\] _04179_ _04182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06355_ _00597_ _01742_ _01834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05306_ cpu.regs\[4\]\[2\] cpu.regs\[5\]\[2\] cpu.regs\[6\]\[2\] cpu.regs\[7\]\[2\]
+ _00569_ _00574_ _00815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_32_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09074_ _04128_ cpu.ROM_addr_buff\[0\] _04023_ _04129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06286_ _01435_ _01756_ _01760_ _01322_ _01765_ _01766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_31_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08025_ _03296_ _03298_ _00223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05237_ _00750_ _00751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05168_ _00683_ _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08738__A1 _02727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09976_ _02634_ _04927_ _04928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05099_ cpu.regs\[1\]\[6\] _00618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08927_ cpu.timer_div\[3\] _04000_ _04007_ _04003_ _04008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08498__C _03653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05972__A1 _01015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08858_ _03167_ _03953_ _03954_ _03956_ _03957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07809_ _02516_ _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08910__A1 _02727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08789_ _02697_ _03894_ _03895_ _03897_ _03898_ _03899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_79_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_98_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_98_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_82_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_27_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_27_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_23_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09218__A2 _02796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08977__A1 cpu.uart.divisor\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06452__A2 _01296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07401__A1 _02592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10116_ _00015_ clknet_leaf_2_wb_clk_i cpu.regs\[9\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10047_ _02427_ _04735_ _04988_ _02433_ _04989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09154__A1 _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09457__A2 _00701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05132__I net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06140_ _01103_ _01621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06391__C _01121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06071_ _01549_ _01552_ _01553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_1_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09830_ _04811_ _02416_ _04806_ _04816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__06898__I _00619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09761_ _02420_ _04759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06973_ _02444_ _02445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05954__A1 _01435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09145__A1 _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08712_ cpu.timer_div_counter\[6\] _03834_ _03837_ _00371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05924_ cpu.pwm_top\[1\] _01251_ _01407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09692_ _04696_ _04699_ _04701_ _04702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05307__I cpu.regs\[1\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer12 _00955_ net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_107_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08643_ _03514_ _03787_ _03788_ _00351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05855_ _01338_ _01339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05182__A2 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05786_ _01267_ _01269_ _01270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08574_ _03721_ cpu.toggle_top\[7\] _03737_ _03738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_1_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07525_ _02913_ _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_37_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10088__C _04931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07456_ cpu.uart.receive_counter\[0\] _02864_ _02866_ _02867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_9_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06407_ cpu.timer_top\[14\] _01404_ _01621_ _01884_ _01885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_20_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07387_ _02802_ _02803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08959__A1 _02816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09126_ _04167_ _00455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_60_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07397__C _02763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06338_ _01774_ _01164_ _01815_ _01816_ _01817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_118_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_31_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09057_ _04114_ _04116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09620__A2 _01155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06269_ _01746_ _01748_ _01749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08008_ _02812_ _03288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_13_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09959_ _04914_ _04915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05645__C _01001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09912__I _04868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09687__A2 cpu.ROM_addr_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output46_I net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09439__A2 _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05661__B _01107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06122__A1 cpu.uart.divisor\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_70_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06048__I _00826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10665_ _00559_ clknet_leaf_3_wb_clk_i cpu.regs\[15\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_97_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10596_ _00490_ clknet_leaf_70_wb_clk_i cpu.mem_cycle\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput70 net70 io_out[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput81 net81 io_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput92 net92 sram_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07607__I _02963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10180__D _00075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_qcpu_99 io_oeb[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_77_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05640_ _01118_ _01122_ _01123_ _01124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_59_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06361__A1 _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05571_ _01043_ _01055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__05795__S0 _00864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_13_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07310_ _00925_ _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08290_ _03515_ net15 _03516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_85_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07241_ _02655_ _02684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer5_I _00875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07172_ _02622_ _02623_ _02625_ _02626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06123_ _01193_ _01603_ _01604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06054_ _01333_ _01430_ _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_115_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09813_ cpu.ROM_spi_dat_out\[6\] _04778_ _04802_ _04788_ _04803_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_6_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09744_ _03276_ _04745_ _04746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06956_ _02426_ _02427_ _02428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05907_ _01192_ _01388_ _01389_ _01390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09675_ cpu.last_addr\[11\] _04681_ _04685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06887_ _02362_ _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__08341__A2 _03518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05838_ _01321_ _01322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08626_ cpu.toggle_ctr\[13\] _03776_ _03777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_68_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05769_ cpu.pwm_top\[0\] _01251_ _01252_ _01253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_49_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08557_ cpu.toggle_ctr\[7\] _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_76_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08488_ _03649_ _03667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07508_ _01584_ _02900_ _02904_ _00100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07439_ cpu.uart.receive_div_counter\[14\] _02850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10450_ _00345_ clknet_leaf_4_wb_clk_i cpu.toggle_ctr\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09109_ _04155_ _00450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05500__I _00985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10381_ _00276_ clknet_leaf_43_wb_clk_i cpu.uart.receive_buff\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07604__A1 _01158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07080__A2 _02361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05091__A1 _00567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_42_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_42_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_87_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10648_ _00542_ clknet_leaf_60_wb_clk_i cpu.PORTA_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_70_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09596__A1 _00971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer3 net127 net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05410__I _00899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10579_ _00473_ clknet_leaf_90_wb_clk_i cpu.PC\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_51_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07790_ _02602_ _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08571__A2 cpu.toggle_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06810_ _02281_ _02280_ _02286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_64_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06741_ _00601_ net116 _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_39_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09460_ cpu.PC\[6\] _01019_ _04478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_104_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08411_ _03608_ _03611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05137__A2 cpu.base_address\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06672_ _02145_ _02147_ _02148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09391_ _02093_ _04409_ _04411_ _04412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_19_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05623_ _01013_ _01107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08342_ _03552_ _03555_ _00283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_117_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05554_ _00676_ _01038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08273_ _02642_ _03468_ _03503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06637__A2 _00976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05485_ _00940_ _00943_ _00972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07224_ _02667_ _02659_ _02660_ _02669_ _02670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_6_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07956__B _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07155_ _02609_ _00756_ _02610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09587__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07062__A2 _02361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07086_ _02044_ _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06106_ _01586_ _01587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06037_ _01485_ _01178_ _01517_ _01518_ _01367_ _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_07988_ _03271_ _00213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08562__A2 _01410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_114_Right_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09727_ cpu.startup_cycle\[0\] _04731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_06939_ net20 _02042_ _02407_ _02412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_97_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09658_ _04575_ _04665_ _04667_ _04668_ _04669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09589_ _03081_ _04601_ _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08609_ _03756_ _03765_ _03766_ _00339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_49_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10502_ _00397_ clknet_leaf_8_wb_clk_i cpu.timer_capture\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10433_ _00328_ clknet_leaf_11_wb_clk_i cpu.toggle_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10364_ _00259_ clknet_leaf_46_wb_clk_i cpu.uart.counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10295_ _00190_ clknet_leaf_49_wb_clk_i cpu.spi.dout\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05454__I3 cpu.regs\[11\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09502__A1 _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05270_ _00772_ _00695_ _00782_ _00783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_70_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09569__A1 _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08960_ _04033_ _00423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07911_ _02873_ cpu.spi.busy _03208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08891_ _03982_ _03983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_110_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07842_ _03139_ cpu.timer\[9\] cpu.timer\[8\] _03140_ _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07773_ cpu.PC\[11\] _03081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09512_ cpu.PC\[7\] cpu.br_rel_dest\[7\] _04528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_91_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06724_ _02163_ _02164_ _02166_ _02200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_65_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09443_ _04456_ _04460_ _04461_ _00767_ _04462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06655_ _00618_ _00934_ _02131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_87_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05606_ _01050_ _01040_ _01090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09374_ _02803_ _01587_ _04394_ _04395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08325_ _03532_ _03541_ _00280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06586_ _02046_ _02061_ _02062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05537_ _01009_ _00747_ _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_47_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08256_ cpu.uart.data_buff\[3\] _03484_ _03489_ _03490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08480__A1 _02570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05468_ _00004_ _00955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__05050__I _00570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08187_ cpu.uart.div_counter\[11\] _03405_ _03432_ _03408_ _03433_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07207_ _02654_ _00049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07138_ _00692_ _02540_ _02597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_61_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05399_ _00883_ _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_30_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07069_ cpu.rom_data_dist _02536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_30_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10080_ _01440_ _05010_ _05020_ _01548_ _01529_ _05021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_69_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09263__A3 _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09795__C _04788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08471__A1 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05895__I _01113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10416_ _00311_ clknet_leaf_90_wb_clk_i cpu.orig_PC\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09367__I _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10347_ _00242_ clknet_leaf_31_wb_clk_i cpu.uart.div_counter\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09971__A1 _03231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05588__A2 _00717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10278_ _00173_ clknet_leaf_111_wb_clk_i cpu.regs\[4\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_49_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06440_ _00654_ _01917_ _01918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06394__C _01871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06371_ _01846_ _01849_ _01850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08110_ _03196_ _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09090_ _04137_ _00591_ _04141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05322_ _00829_ _00830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08041_ cpu.uart.dout\[3\] _03309_ _03310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05253_ _00766_ _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_31_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05371__S1 _00860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10021__A1 _00778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05184_ cpu.instr_cycle\[3\] _00695_ _00698_ _00699_ _00700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_24_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09992_ _02470_ _00729_ _04939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09962__A1 cpu.PORTA_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08943_ _02606_ _01020_ _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08874_ _03969_ _00401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07525__I _02913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07825_ cpu.timer_div\[0\] _03121_ cpu.timer_div_counter\[2\] _03122_ _03123_ _03124_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_79_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07756_ net12 _03055_ _03065_ _02406_ _03066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__10088__A1 _01262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06707_ _02180_ _02181_ _02183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09426_ _04443_ _04423_ _04445_ _04413_ _04414_ _04446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_07687_ _03017_ _00166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05503__A2 _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06638_ _02063_ _02064_ _02113_ _02114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09357_ _04377_ _04378_ _03868_ _00475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06569_ _02044_ _02045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08308_ _03525_ _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09288_ _02781_ _01364_ _04310_ _04311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08239_ _03475_ _00260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_105_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10012__B2 cpu.ROM_addr_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10012__A1 cpu.ROM_addr_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10201_ _00096_ clknet_leaf_121_wb_clk_i cpu.regs\[14\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output76_I net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10132_ _00031_ clknet_leaf_101_wb_clk_i cpu.regs\[1\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05114__S1 _00631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10063_ _01263_ _04251_ _01099_ _01170_ _04213_ _05004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_89_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07170__I _00903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08692__A1 _03822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08995__A2 _01110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10003__A1 cpu.ROM_addr_buff\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05940_ _01421_ _01422_ _01173_ _01423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05871_ net26 _01012_ _01355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08590_ _03749_ _03753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07610_ cpu.regs\[8\]\[1\] _02966_ _02968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_109_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05733__A2 _01216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07541_ _01935_ cpu.regs\[12\]\[6\] _02913_ _02926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06930__A1 _01934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06930__B2 cpu.regs\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07472_ cpu.uart.receive_counter\[3\] cpu.uart.receive_counter\[2\] _02868_ _02880_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_72_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07730__I0 _03006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09211_ _00950_ _00986_ _01687_ _01785_ _04236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_06423_ _01898_ _01900_ _01901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09142_ _03378_ _04180_ _04181_ _00457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06354_ _01446_ _01832_ _01833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05305_ _00814_ net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_114_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_21_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09073_ _00790_ _02768_ _00728_ _04128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06285_ _01468_ _01762_ _01764_ _01765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_114_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08024_ cpu.spi.data_in_buff\[5\] _03198_ _03294_ cpu.spi.data_in_buff\[6\] _03298_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05236_ _00742_ _00749_ _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_25_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09935__A1 cpu.PORTB_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05167_ _00682_ _00683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09975_ _04914_ _04927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05098_ cpu.regs\[4\]\[6\] cpu.regs\[5\]\[6\] cpu.regs\[6\]\[6\] cpu.regs\[7\]\[6\]
+ _00615_ _00616_ _00617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08926_ _02742_ _03997_ _04007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08857_ _02668_ _03955_ _03956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07808_ _01691_ _03102_ _03110_ _00194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08788_ _03864_ _03898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05280__S0 _00785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07739_ _02034_ _02446_ _02581_ _03050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_67_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_60_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07477__A2 _01145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09409_ _04334_ _04422_ _04428_ _04345_ _04429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_23_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_67_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_67_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_90_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07165__I _02516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10115_ _00014_ clknet_leaf_2_wb_clk_i cpu.regs\[9\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10046_ _04743_ _04731_ _04988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05963__A2 _00929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_59_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06912__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05413__I _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09209__A3 _04230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06244__I _00596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06070_ _01550_ _01551_ _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_1 _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09917__A1 _04045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_105_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09760_ _04755_ _04751_ _04752_ _04758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06972_ _02032_ _02443_ _02444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09691_ cpu.last_addr\[2\] cpu.ROM_addr_buff\[2\] _04700_ _04701_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08711_ cpu.timer_div_counter\[6\] _03834_ _03836_ _03201_ _03837_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05923_ cpu.timer_top\[9\] _01179_ _01180_ _01406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_83_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08642_ cpu.pwm_counter\[1\] cpu.pwm_counter\[0\] cpu.pwm_counter\[2\] _03788_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__10480__CLK clknet_leaf_18_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09290__I _04270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer13 _02327_ net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05854_ _01337_ _01338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_89_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08573_ _03724_ _03735_ _03736_ _03737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05785_ _00656_ _01011_ _01268_ _01269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_88_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08656__A1 _02882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07524_ _02914_ _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07455_ cpu.uart.receiving net15 _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_91_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06406_ _01864_ _01616_ _01882_ _01883_ _01246_ _01884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_57_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07386_ cpu.PC\[3\] _02802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09125_ _04166_ cpu.ROM_addr_buff\[13\] _04159_ _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06337_ _00986_ _01278_ _01721_ _01816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_118_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09056_ _04114_ _04115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07631__A2 _02981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06268_ net94 _01747_ _01748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08007_ _03286_ _03287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05219_ _00708_ _00734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06199_ _01679_ _01680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_9_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09958_ _01042_ _04842_ _04914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08909_ cpu.spi.divisor\[7\] _03990_ _03994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05945__A2 _00799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09889_ _04863_ _00522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07147__A1 _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_114_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_114_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_56_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output39_I net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08647__A1 _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10664_ _00558_ clknet_leaf_3_wb_clk_i cpu.regs\[15\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10595_ _00489_ clknet_leaf_69_wb_clk_i cpu.mem_cycle\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05633__A1 _01081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput60 net60 io_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput71 net71 io_out[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput82 net82 io_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput93 net93 sram_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07138__A1 _00692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10029_ _02453_ _04967_ _04969_ _04971_ _04972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_86_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05570_ _00644_ _01054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_58_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05795__S1 _00865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07240_ _02683_ _00053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07861__A2 cpu.timer\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07171_ _02624_ _02616_ _02625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05872__A1 _01012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06122_ cpu.uart.divisor\[11\] _01220_ _01603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05624__A1 _01015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06053_ _01533_ _01534_ _01535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_100_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09812_ _04780_ _04801_ _04802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_6_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05318__I _00826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09743_ _02438_ _04744_ _04745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06955_ _00664_ _02427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07129__A1 _01015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05906_ cpu.uart.has_byte _01192_ _01389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09674_ cpu.ROM_addr_buff\[13\] _04683_ _04684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06886_ _02359_ _02361_ _02021_ _02362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_05837_ _00655_ _01320_ _01321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08625_ _03750_ _03775_ _03776_ _00345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_68_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08556_ cpu.toggle_ctr\[15\] _03717_ _03720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_81_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05768_ _01097_ _01252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07507_ cpu.regs\[13\]\[2\] _02901_ _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08487_ cpu.orig_PC\[9\] _03659_ _03666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05699_ _01054_ _01077_ _01036_ _01060_ _01183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_07438_ _02844_ _02848_ _02849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09054__A1 _00693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07369_ _02786_ _02778_ _02775_ _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09108_ _04154_ cpu.ROM_addr_buff\[8\] _04148_ _04155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_33_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10380_ _00275_ clknet_leaf_44_wb_clk_i cpu.uart.receive_buff\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09039_ _04084_ _04101_ _00434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_92_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07368__A1 _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07644__S _02978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05474__S0 _00956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06040__B2 _00909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06487__C _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_82_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_82_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_67_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_11_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_11_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_31_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10647_ _00541_ clknet_leaf_60_wb_clk_i cpu.PORTA_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_82_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09045__B2 _01957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer4 _02384_ net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10578_ _00472_ clknet_leaf_92_wb_clk_i cpu.Z vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_11_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08859__A1 cpu.timer_capture\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06740_ _02214_ _02215_ _02216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_39_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06671_ _02137_ _02146_ _02147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09989__B cpu.ROM_spi_mode vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08410_ _03609_ _03610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05622_ _01024_ _01065_ _01073_ _01105_ _01106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_80_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09390_ _04410_ _04386_ _04411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_19_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08341_ cpu.uart.receive_div_counter\[3\] _03518_ _03553_ _03554_ _03555_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_86_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05553_ _01036_ _01037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_74_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09284__A1 _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08272_ _03499_ _03501_ _03502_ _00266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_74_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05484_ _00970_ _00971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07223_ _02668_ _02661_ _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09036__A1 _01110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08912__I _03995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07154_ _01008_ _02609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06105_ cpu.br_rel_dest\[3\] _01586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_30_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07085_ _02550_ _02056_ _02551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06036_ cpu.pwm_top\[2\] _01251_ _01252_ _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05073__A2 _00592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07528__I _01481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07987_ cpu.spi.div_counter\[4\] _03264_ _03270_ _02753_ _03271_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09726_ _04673_ _04729_ _04730_ _02762_ _00492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06938_ _02410_ _02359_ _02411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09657_ _02513_ _04650_ _04227_ _04668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06869_ _02332_ _02344_ _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07522__A1 _02885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08608_ _03723_ _03762_ _03766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09588_ _02047_ _03071_ _04420_ _04601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_38_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08539_ cpu.toggle_ctr\[10\] _03703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10501_ _00396_ clknet_leaf_24_wb_clk_i cpu.timer\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10432_ _00327_ clknet_leaf_9_wb_clk_i cpu.toggle_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10363_ _00258_ clknet_leaf_64_wb_clk_i cpu.uart.counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08538__B1 _01256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10294_ _00189_ clknet_leaf_103_wb_clk_i cpu.regs\[2\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06013__A1 net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06252__A1 _01331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07910_ _02870_ _03207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08890_ _03200_ _03209_ _01051_ _02729_ _03982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_07841_ cpu.timer_top\[8\] _03140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07772_ _03069_ _03079_ _03080_ _00188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09511_ _04526_ _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06723_ _02197_ _02198_ _02199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_91_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09442_ _04333_ _04451_ _04461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06654_ _00804_ _01287_ _02130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05605_ _01088_ _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09257__A1 _04270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06585_ cpu.PC\[11\] _02047_ _02060_ _02061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09373_ _04339_ _04393_ _04394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08324_ _03537_ _03518_ _03540_ _03541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_74_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05536_ _01019_ _01020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05818__A1 _01162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08255_ _03111_ _03489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05467_ cpu.regs\[12\]\[4\] cpu.regs\[13\]\[4\] cpu.regs\[14\]\[4\] cpu.regs\[15\]\[4\]
+ net123 _00858_ _00954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_08186_ cpu.uart.div_counter\[11\] _03428_ _03432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07206_ _02650_ _02623_ _02653_ _02640_ _02654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_6_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05398_ _00881_ _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_42_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07137_ _02595_ _02587_ _02596_ _02589_ _00037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_113_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10414__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06243__A1 _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_18_Left_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07068_ _02391_ _02535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06019_ net8 _01371_ _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_97_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09709_ _02463_ _02538_ _04671_ _04717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_69_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_27_Left_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_87_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09248__A1 _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10415_ _00310_ clknet_leaf_90_wb_clk_i cpu.orig_PC\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_36_Left_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10346_ _00241_ clknet_leaf_32_wb_clk_i cpu.uart.div_counter\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07982__A1 _02882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10277_ _00172_ clknet_leaf_109_wb_clk_i cpu.regs\[4\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06021__B _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_45_Left_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_0_0_wb_clk_i clknet_0_wb_clk_i clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_118_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06370_ _01847_ _01835_ _01848_ _01849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_84_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05321_ cpu.regs\[1\]\[3\] _00829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08040_ _03300_ _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05252_ _00764_ _00765_ _00766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_54_Left_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_11_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05183_ cpu.TIE cpu.needs_timer_interrupt _00699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_51_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09991_ _04759_ _02429_ _02460_ _04938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_86_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08942_ _04018_ _00420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09507__B _04523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_63_Left_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08873_ cpu.timer_capture\[12\] _03965_ _03967_ _03968_ _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07725__A1 _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07824_ cpu.timer_div\[0\] _03121_ _03119_ cpu.timer_div\[1\] _03123_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07755_ _02552_ _03061_ _03064_ _03055_ _03065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_07686_ _03002_ cpu.regs\[5\]\[4\] _03010_ _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06706_ _02180_ _02181_ _02182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_clkbuf_leaf_50_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09425_ _02334_ _04409_ _04444_ _04445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06637_ _00634_ _00976_ _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09356_ _02789_ _04297_ _04378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06568_ _02043_ _02044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08307_ _03519_ _03529_ _00274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_72_Left_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05519_ _01003_ _01004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06499_ _01938_ _01939_ _01975_ _01976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_35_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09287_ cpu.PC\[0\] cpu.br_rel_dest\[0\] _04310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08238_ cpu.uart.counter\[3\] _03469_ _03471_ _03473_ _03474_ _03475_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_105_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05267__A2 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05996__I _01478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08169_ cpu.uart.div_counter\[7\] _03392_ _03414_ _03419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_10200_ _00095_ clknet_leaf_123_wb_clk_i cpu.regs\[14\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10131_ _00030_ clknet_leaf_101_wb_clk_i cpu.regs\[1\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output69_I net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10062_ cpu.orig_flags\[0\] _04073_ _04253_ _05002_ _05003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_89_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09469__A1 _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08141__A1 _03296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06016__B _01122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10329_ _00224_ clknet_leaf_52_wb_clk_i cpu.spi.data_in_buff\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05870_ _01297_ net90 _01353_ _01354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__09841__I net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07540_ _02925_ _00111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07471_ _02877_ _02866_ _02878_ _02879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_118_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09210_ _01939_ _01346_ _00711_ _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_06422_ _01899_ _01900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09141_ cpu.last_addr\[1\] _04177_ _04181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06353_ _01819_ _01830_ _01832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08192__I _03275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09072_ _04127_ _00441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09632__A1 _04327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05304_ _00566_ _00808_ _00813_ _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_32_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08023_ _03296_ _03297_ _00222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06284_ _01731_ _01763_ _01764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_102_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05235_ _00743_ _00658_ _00748_ _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_40_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08920__I _04002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05166_ _00649_ _00682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_40_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09974_ _04914_ _04926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05421__A2 _00909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05097_ _00575_ _00616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08925_ _03122_ _04000_ _04005_ _04006_ _00415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_input20_I io_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08856_ _03945_ _03955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07807_ cpu.spi.data_in_buff\[4\] _03107_ _03105_ _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05185__A1 _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08787_ _03856_ _03896_ _03897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05999_ _01481_ _01482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07738_ _02534_ _03048_ _03049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05280__S1 _00786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07669_ _01933_ _03006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_39_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09408_ _04425_ _04426_ _04427_ _04428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_23_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09339_ _00749_ _04361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_51_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_109_Right_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09623__A1 _04309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06437__A1 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_36_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_36_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10114_ _00013_ clknet_leaf_2_wb_clk_i cpu.regs\[9\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10045_ _02479_ _04986_ _04987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_59_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06912__A2 _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09610__B _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06676__A1 _02150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09090__A2 _00591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06971_ cpu.mem_cycle\[4\] _02443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09690_ cpu.last_addr\[1\] _04174_ _04700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08710_ _03131_ _03836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05922_ cpu.timer_top\[1\] _01240_ _01400_ _01403_ _01404_ _01405_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_83_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08641_ _03784_ _03783_ _03786_ _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05853_ _00655_ _01328_ _01337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_89_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer14 _02246_ net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_77_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05784_ _00704_ _00755_ _01268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08572_ _03721_ cpu.toggle_top\[7\] _03736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07523_ _02913_ _02914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07454_ cpu.uart.receive_counter\[0\] _02864_ _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_76_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06405_ cpu.timer_capture\[14\] _01233_ _01239_ _01883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07385_ _02392_ _02314_ _02800_ _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_32_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09124_ cpu.regs\[3\]\[5\] _03674_ _00727_ _04166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06336_ _01416_ _01785_ _01814_ _01589_ _01815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_17_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09055_ _02537_ _03050_ _04113_ _02493_ _04114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_06267_ _01744_ _01745_ _01747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08006_ _03197_ _03211_ _03286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05218_ _00729_ _00732_ _00733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__05642__A2 _01120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06198_ _01678_ _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05149_ cpu.mem_cycle\[5\] cpu.mem_cycle\[4\] cpu.mem_cycle\[3\] cpu.mem_cycle\[2\]
+ _00666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_09957_ _04913_ _00540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08908_ _02647_ _03989_ _03993_ _00411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09888_ net64 _04856_ _04860_ _04862_ _04863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_99_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08839_ _03176_ _03939_ _03860_ _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_56_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10663_ _00557_ clknet_leaf_61_wb_clk_i net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05330__A1 _00581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_97_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10594_ _00488_ clknet_leaf_79_wb_clk_i cpu.mem_cycle\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput61 net61 io_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput50 net50 io_oeb[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput72 net72 io_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput94 net94 sram_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput83 net83 sram_addr[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10028_ _00667_ _04970_ _04729_ _04971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_37_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07170_ _00903_ _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_26_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06121_ _01592_ _01383_ _01600_ _01601_ _01220_ _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_14_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06052_ _01530_ _00923_ _01534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__05624__A2 _01106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09811_ cpu.ROM_spi_dat_out\[5\] _02489_ _04785_ _04800_ _04801_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09742_ _04743_ _04734_ _02419_ _04744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_94_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06954_ _00662_ _02426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05905_ _01369_ _01386_ _01387_ _01388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09673_ cpu.last_addr\[13\] _04682_ _04683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06885_ _02360_ _02361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05836_ _01300_ _01320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08624_ cpu.toggle_ctr\[12\] _03774_ _03776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_77_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05767_ _01103_ _01251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08555_ _03713_ _03716_ _03718_ _03719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_81_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07506_ _01482_ _02900_ _02903_ _00099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05698_ _01181_ _01182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08486_ _03664_ _03657_ _03665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_13_0_wb_clk_i clknet_0_wb_clk_i clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07437_ _02845_ _02846_ cpu.uart.receive_div_counter\[14\] _02847_ _02848_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_92_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07368_ _01480_ _02764_ _02785_ _02786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06319_ _01224_ _01797_ _01798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09107_ _03045_ _04136_ _04153_ _04154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07299_ _01039_ _01038_ _02729_ _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_5_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09038_ _01039_ _04097_ _04099_ _04100_ _04101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_13_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output51_I net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05474__S1 _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06879__A1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09117__I0 cpu.regs\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05244__I _00757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10646_ _00540_ clknet_leaf_69_wb_clk_i cpu.PORTB_DDR\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xrebuffer5 _00875_ net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_106_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_51_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_51_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10577_ _00471_ clknet_leaf_58_wb_clk_i cpu.IE vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08223__C _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05419__I _00907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06670_ _02143_ _02144_ _02146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05621_ _01081_ _01086_ _01098_ _01104_ _01105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_59_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08340_ _02822_ _03548_ _03554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05552_ _01027_ _01036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08271_ cpu.uart.data_buff\[6\] _03497_ _03489_ _03502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05483_ _00969_ _00970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07222_ _00909_ _02668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_13_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07153_ cpu.uart.divisor\[0\] _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_89_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07809__I _02516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06104_ _01160_ _01584_ _01585_ _00015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07084_ _02549_ _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_14_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06035_ cpu.timer_top\[10\] _01179_ _01514_ _01516_ _01180_ _01517_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_23_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07986_ _03203_ _03268_ _03269_ _03270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09725_ _02031_ _04723_ _04730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06937_ _02409_ _02399_ _02410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05908__I0 _01390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09656_ _04594_ _04650_ _04666_ _04374_ _04667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08607_ _03723_ _03762_ _03765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06868_ _02336_ _02343_ _02344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09587_ _03082_ _04550_ _04600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06799_ _02269_ _02274_ _02275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05819_ _01111_ _00799_ _01303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05999__I _01481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08538_ cpu.toggle_ctr\[9\] _03701_ _01256_ cpu.toggle_ctr\[8\] _03702_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08469_ _02803_ _03651_ _03652_ _03653_ _00312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_108_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10500_ _00395_ clknet_leaf_8_wb_clk_i cpu.timer\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10431_ _00326_ clknet_leaf_9_wb_clk_i cpu.toggle_top\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10362_ _00257_ clknet_leaf_64_wb_clk_i cpu.uart.counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06261__A2 net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10293_ _00188_ clknet_leaf_103_wb_clk_i cpu.regs\[2\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05383__S0 _00856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10629_ _00523_ clknet_leaf_68_wb_clk_i net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_52_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07840_ cpu.timer_top\[9\] _03139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07771_ _00818_ _03069_ _03080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09510_ _04524_ _04500_ _04526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06722_ cpu.regs\[1\]\[0\] _00997_ _02198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_40_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09441_ _02549_ _01774_ _04459_ _04460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06653_ _02126_ _02127_ _02129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_115_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05604_ _01087_ _01085_ _01088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_65_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09372_ _04337_ _04338_ _04393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06584_ cpu.PC\[9\] _02059_ _02060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08323_ _03537_ _03539_ _03540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05535_ cpu.br_rel_dest\[6\] _01019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08254_ cpu.uart.data_buff\[2\] _03469_ _03487_ _03488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05466_ _00953_ net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08185_ _03427_ _03431_ _00250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07205_ _02652_ _02636_ _02653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05397_ _00863_ _00887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07136_ _01135_ _02585_ _02596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_113_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07067_ _02522_ _02534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_112_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06018_ _01492_ _01035_ _01498_ _01499_ _01371_ _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_11_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09193__A1 _03231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08940__A1 _02652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09708_ _02538_ _04673_ _02463_ _04716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07969_ cpu.spi.div_counter\[1\] _03256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05754__A1 _01046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_87_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09639_ _04649_ _04650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07259__A1 _02697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09929__I _04891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_41_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10239__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10414_ _00309_ clknet_4_9_0_wb_clk_i cpu.orig_PC\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05117__S0 _00630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10345_ _00240_ clknet_leaf_32_wb_clk_i cpu.uart.div_counter\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_70_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05588__A4 _01071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05993__A1 net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10276_ _00171_ clknet_leaf_110_wb_clk_i cpu.regs\[4\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_124_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05320_ cpu.regs\[4\]\[3\] cpu.regs\[5\]\[3\] cpu.regs\[6\]\[3\] cpu.regs\[7\]\[3\]
+ _00570_ _00827_ _00828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_71_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05251_ _00707_ _00651_ _00765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05182_ _00697_ net18 _00694_ _00698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_7_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09411__A2 _04068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07422__B2 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09990_ _03822_ _04937_ _00549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08941_ cpu.timer_div\[7\] _03996_ _04017_ _04015_ _04018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_50_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08872_ _03808_ _03968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07823_ cpu.timer_div\[2\] _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_07754_ _02351_ _03063_ _03064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09242__C _03920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06705_ _02140_ _02141_ _02181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07685_ _02987_ _03011_ _03016_ _00165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09424_ _04410_ _04423_ _04444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06636_ _02109_ _02111_ _02112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05342__I cpu.PORTA_DDR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09355_ _04328_ _04367_ _04376_ _04377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06567_ _00846_ _01001_ _01296_ _01071_ _02043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_118_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08306_ cpu.uart.receive_buff\[2\] _03523_ _03526_ cpu.uart.receive_buff\[3\] _03529_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09286_ _04308_ _04309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05518_ _00878_ _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06498_ _01315_ _01952_ _01970_ _01974_ _01975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_34_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08237_ _02619_ _03474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05449_ _00936_ _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07269__I _02707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08168_ _03391_ _03417_ _03393_ _03418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_108_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_108_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_15_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08099_ cpu.uart.counter\[3\] cpu.uart.counter\[2\] _03363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07119_ _02031_ _02462_ _02450_ _02582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_101_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10130_ _00029_ clknet_leaf_85_wb_clk_i cpu.instr_buff\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05975__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10061_ _04998_ _04254_ _05001_ _05002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05517__I _01001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09469__A2 _04349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07400__C _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07179__I _00952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10328_ _00223_ clknet_leaf_51_wb_clk_i cpu.spi.data_in_buff\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05966__A1 _01441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08904__A1 _02635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Left_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10259_ _00154_ clknet_leaf_12_wb_clk_i cpu.regs\[6\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09062__C _04050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07470_ cpu.uart.receive_counter\[2\] _02868_ _02878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_88_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06421_ _00628_ _01783_ _01899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09140_ cpu.ROM_addr_buff\[1\] _04179_ _04180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_6_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_6_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06352_ _01818_ _01830_ _01831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05329__S0 _00569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09071_ _00971_ _04115_ _04126_ _04124_ _04127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_44_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06283_ _01669_ _01761_ _01763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05303_ _00003_ _00810_ _00812_ _00813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08022_ cpu.spi.data_in_buff\[4\] _03291_ _03294_ cpu.spi.data_in_buff\[5\] _03297_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05234_ _00747_ _00748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05165_ _00681_ _00012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09973_ _04925_ _00544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_73_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05096_ _00598_ _00615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08924_ _02723_ _04006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09148__A1 cpu.ROM_addr_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08855_ _03942_ _03954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07806_ _01610_ _03102_ _03109_ _00193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08786_ _02691_ _03884_ _02697_ _03896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input13_I io_in[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07737_ _02325_ _03047_ _03048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05998_ _01480_ _01481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_95_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06134__A1 _01591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07668_ _03005_ _00159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_109_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09407_ _04425_ _04426_ _04341_ _04427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06619_ _02093_ _01288_ _02094_ _02095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07599_ _02017_ _02960_ _00134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09338_ cpu.orig_PC\[2\] _04359_ _04360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_51_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09269_ _04291_ _04286_ _04290_ _04293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_50_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09428__B _04417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output81_I net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10113_ _02014_ _05036_ _05044_ _00565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08986__C _04050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_76_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_76_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10044_ _00693_ _04985_ _02481_ _04986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_59_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06373__A1 _01435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09862__A2 _02729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09389__I _04319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06541__I _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05939__A1 cpu.Z vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06970_ _02028_ _02442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_67_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input5_I io_in[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05921_ _01246_ _01404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08640_ cpu.pwm_counter\[2\] _03786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09550__A1 _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05852_ _01335_ _01336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06364__B2 _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06364__A1 _01438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05783_ _01016_ _01267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08571_ _03723_ cpu.toggle_top\[6\] cpu.toggle_top\[5\] _03725_ _03734_ _03735_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09801__B _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06116__A1 net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07522_ _02885_ _02912_ _02913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_07453_ cpu.uart.receiving _02863_ _02864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06404_ cpu.timer_capture\[6\] _01690_ _01879_ _01881_ _01242_ _01882_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_64_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09123_ _04165_ _00454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07384_ _02311_ _02799_ _02313_ _02800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_29_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06335_ _01414_ _01813_ _01814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09054_ _00693_ _03050_ _04113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06266_ _01724_ _01744_ _01745_ _01746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_32_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08005_ net16 _03285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05217_ _00668_ _00730_ _00731_ _00688_ _00732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_102_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06197_ _01588_ _01632_ _01677_ _01479_ _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_05148_ _00662_ _00663_ _00664_ _00665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_110_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09956_ cpu.PORTB_DDR\[7\] _04903_ _04912_ _04908_ _04913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05079_ _00575_ _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09887_ _04861_ _04862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08907_ cpu.spi.divisor\[6\] _03990_ _03993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08838_ cpu.timer\[15\] _03938_ _03939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_56_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08769_ cpu.timer\[3\] _03876_ _03880_ _03858_ _03881_ _03882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_68_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06107__A1 _01587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_36_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09002__I _04068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_123_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_123_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10662_ _00556_ clknet_4_10_0_wb_clk_i cpu.C vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05530__I _01013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10593_ _00487_ clknet_leaf_70_wb_clk_i cpu.mem_cycle\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_97_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05633__A3 _01114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09080__I0 _00818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput51 net51 io_oeb[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput40 net40 io_oeb[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput73 net73 io_out[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput62 net62 io_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput84 net84 sram_addr[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput95 net95 sram_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10027_ _02464_ _02582_ _04970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_90_Left_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05705__I _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07192__I _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06120_ net9 _01204_ _01205_ _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_42_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06051_ _01532_ _01533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_117_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_99_Right_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08023__A1 _03296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09810_ _02420_ _04750_ _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08574__A2 cpu.toggle_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09741_ cpu.startup_cycle\[1\] _04743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06953_ _02421_ _02424_ _02425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09582__I _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05904_ cpu.uart.dout\[1\] _00012_ _01387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09523__A1 _01002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09672_ cpu.last_addr\[12\] cpu.last_addr\[11\] _04681_ _04682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06884_ _00743_ _01267_ _01022_ _02360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_27_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05835_ _01170_ _01318_ _01319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08623_ cpu.toggle_ctr\[12\] _03774_ _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_68_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05766_ cpu.timer_top\[8\] _01179_ _01180_ _01249_ _01250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_08554_ cpu.toggle_ctr\[15\] _03717_ _03714_ cpu.toggle_ctr\[14\] _03718_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_81_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07505_ cpu.regs\[13\]\[1\] _02901_ _02903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05697_ _01094_ _01062_ _01181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08485_ _03060_ _03664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_107_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07436_ cpu.uart.divisor\[14\] _02847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__05350__I cpu.PORTB_DDR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07367_ _02521_ _02780_ _02784_ _02785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_33_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06318_ cpu.uart.divisor\[13\] _01489_ _01797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09106_ _04137_ cpu.regs\[3\]\[0\] _04153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07298_ _02609_ _00757_ _02729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_09037_ _04081_ _04100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07277__I _00776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06249_ _01728_ _01727_ _01729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09939_ _04900_ _00535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_output44_I net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06879__A2 _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09117__I1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08057__B _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10645_ _00539_ clknet_leaf_60_wb_clk_i cpu.PORTB_DDR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08253__A1 _00904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10576_ _00470_ clknet_leaf_57_wb_clk_i cpu.TIE vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer6 _02315_ net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_20_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_20_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09505__A1 _02570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05435__I _00923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_30_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05620_ _01100_ _01102_ _01103_ _01104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_86_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_19_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07819__A1 cpu.timer_div\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05551_ _01034_ _01035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_80_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08270_ cpu.uart.data_buff\[5\] _03491_ _03500_ _03501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05482_ cpu.base_address\[3\] _00969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_27_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07221_ _02666_ _02667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_30_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08244__A1 _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07047__A2 _02514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07152_ _02595_ _02600_ _02607_ _02603_ _00041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_42_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06103_ cpu.regs\[9\]\[2\] _01361_ _01585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07083_ cpu.PC\[5\] _02549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06034_ _01179_ _01515_ _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09744__A1 _03276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07985_ cpu.spi.div_counter\[4\] _03251_ _03269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09724_ _04169_ _04674_ _04729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05345__I cpu.PORTA_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06936_ _02395_ _02408_ _02396_ _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09655_ _00604_ _04596_ _04666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06867_ _02337_ _02342_ _02343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08606_ _03764_ _00338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05818_ _01162_ _00800_ _01302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_96_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09586_ _04574_ _04599_ _04523_ _00483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06798_ _02270_ _00976_ _02273_ _02274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05749_ _01232_ _01233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08537_ cpu.toggle_top\[9\] _03701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_37_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08468_ _02761_ _03653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07419_ cpu.uart.receive_div_counter\[8\] _02830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08399_ cpu.uart.receive_div_counter\[15\] _03597_ _03601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10430_ _00325_ clknet_leaf_9_wb_clk_i cpu.toggle_top\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10361_ _00256_ clknet_leaf_47_wb_clk_i cpu.uart.has_byte vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09983__A1 _02646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10292_ _00187_ clknet_leaf_107_wb_clk_i cpu.regs\[2\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07746__B1 _03054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_114_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05383__S1 _00860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10628_ _00522_ clknet_leaf_68_wb_clk_i net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07029__A2 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10559_ _00453_ clknet_leaf_87_wb_clk_i cpu.ROM_addr_buff\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08250__B _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07770_ _01582_ _03078_ _02023_ _03079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05165__I _00681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06721_ _00804_ _00964_ _02197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09440_ _04425_ _04457_ _04458_ _04459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06652_ _02126_ _02127_ _02128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06712__A1 cpu.regs\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05603_ _01026_ _01028_ _01087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_65_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09371_ _04273_ _04392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05071__S0 _00571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06583_ _02048_ _02058_ _02059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08322_ _03538_ _03539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05534_ cpu.br_rel_dest\[7\] _01018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08253_ _00904_ _03486_ _03487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07204_ _02651_ _02652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05465_ _00928_ _00939_ _00952_ _00953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_62_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08184_ cpu.uart.div_counter\[10\] _03389_ _03429_ _03430_ _03431_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05396_ _00880_ _00885_ _00886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07135_ _02514_ _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07066_ _02017_ _02521_ _02532_ _02533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06017_ net61 _01069_ _01216_ _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_76_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05451__A1 _00715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09256__B _04279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07968_ _02874_ _03255_ _00209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05203__A1 _00711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09707_ _02027_ _04713_ _04715_ _03920_ _00488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_4_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06919_ _02380_ _02378_ _02393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07899_ cpu.spi.counter\[0\] _03196_ _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_69_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07290__I _02723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09638_ _04648_ _04649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05803__I _01286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09569_ _04333_ _04576_ _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09956__A1 cpu.PORTB_DDR\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10413_ _00308_ clknet_leaf_56_wb_clk_i cpu.orig_flags\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10344_ _00239_ clknet_leaf_64_wb_clk_i cpu.uart.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05117__S1 _00631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10275_ _00170_ clknet_leaf_109_wb_clk_i cpu.regs\[4\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_49_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05250_ _00706_ _00764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05181_ _00696_ _00697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08940_ _02652_ _04009_ _04017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08871_ _03136_ _03953_ _03954_ _03966_ _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07186__A1 _02635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07822_ cpu.timer_div_counter\[0\] _03121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_07753_ net117 _03062_ _03063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06704_ _02177_ _02178_ _02179_ _02180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07684_ cpu.regs\[5\]\[3\] _03010_ _03016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09423_ _02512_ _04443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06635_ _02110_ _02094_ _02111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__05623__I _01013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09354_ _04368_ _04332_ _04372_ _04374_ _04375_ _04376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_47_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08305_ _03519_ _03528_ _00273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07978__C _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06566_ _02041_ _02042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09285_ _00970_ _04272_ _04308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06497_ _01441_ _01947_ _01972_ _01973_ _01974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_05517_ _01001_ _01002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08236_ _03472_ _03473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05448_ _00935_ _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09938__A1 cpu.PORTB_DDR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08167_ _03340_ _03414_ _03417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_90_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07994__B _03276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05672__B2 _01155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07118_ _02026_ _02442_ _02581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05379_ cpu.regs\[12\]\[0\] cpu.regs\[13\]\[0\] cpu.regs\[14\]\[0\] cpu.regs\[15\]\[0\]
+ _00864_ _00865_ _00869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_08098_ cpu.uart.counter\[0\] cpu.uart.counter\[1\] _03362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_101_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07049_ _02516_ _02517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10060_ _04244_ _04999_ _05000_ _05001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05975__A2 _00907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05283__S0 _00785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08844__I _03942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05415__A1 _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10327_ _00222_ clknet_leaf_50_wb_clk_i cpu.spi.data_in_buff\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05708__I _01079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10258_ _00153_ clknet_leaf_118_wb_clk_i cpu.regs\[7\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10189_ _00084_ clknet_leaf_14_wb_clk_i _00002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_109_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05443__I _00930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06420_ _00628_ _01784_ _01898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07340__A1 _02580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08754__I _03859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06351_ _01730_ _01738_ _01820_ _01830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09070_ _02514_ _04116_ _04126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06282_ _01669_ _01730_ _01761_ _01762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__05329__S1 _00827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05302_ _00580_ _00811_ _00812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08021_ _02873_ _03296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08840__A1 cpu.timer_capture\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05233_ _00744_ _00746_ _00718_ _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_4_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05164_ _00647_ _00680_ _00681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09972_ cpu.PORTA_DDR\[3\] _04915_ _04924_ _04920_ _04925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05095_ _00567_ _00614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_0_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08923_ _02675_ _03997_ _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_110_Left_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08929__I _03995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07833__I cpu.TIE vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08854_ _03945_ _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09534__B _04523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07805_ cpu.spi.data_in_buff\[3\] _03107_ _03105_ _03109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08785_ cpu.timer\[6\] cpu.timer\[5\] _03884_ _03895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_05997_ _01366_ _01423_ _01477_ _01479_ _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_07736_ _02265_ _02323_ _02324_ _03047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_79_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05353__I cpu.base_address\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07331__A1 _02755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07667_ _03004_ cpu.regs\[6\]\[5\] _02994_ _03005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09406_ _04418_ _01683_ _04426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06618_ _02090_ _02091_ _02094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07598_ _01680_ _02961_ _00133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05893__A1 _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06549_ cpu.mem_cycle\[1\] _02025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_63_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09337_ _04073_ _04359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_51_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09268_ _04286_ _04290_ _04291_ _04292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08219_ _03452_ _03454_ _03453_ _03457_ _03458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06117__C _01216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05645__A1 _01111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07634__A2 _02981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09199_ _00779_ _04216_ _04217_ _04224_ _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_95_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10581__D _00475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10112_ cpu.regs\[15\]\[7\] _05034_ _05044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10043_ _00690_ _04710_ _04714_ _04985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08898__A1 _02627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07570__A1 _01158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05263__I _00776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_45_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_45_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07322__A1 cpu.toggle_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09378__A2 _00735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07389__A1 _02803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06061__A1 _01364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05920_ _01401_ _01402_ _01240_ _01403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__08749__I _03864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05851_ _01142_ _01334_ _01335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_83_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08570_ _03729_ _03732_ _03733_ _03734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05173__I _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05782_ _01175_ _01255_ _01258_ _01261_ _01265_ _01266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_16_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07521_ _02911_ _02912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_76_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07452_ _02862_ _02863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_92_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06403_ _01612_ _01880_ _01881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07383_ _02307_ _02310_ _02799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09122_ _04164_ cpu.ROM_addr_buff\[12\] _04159_ _04165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_57_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06334_ _01174_ _01811_ _01812_ _01261_ _00986_ _01813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_8_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09053_ _04102_ _04112_ _00437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06265_ _01586_ net93 _01745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_115_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08004_ _02874_ _03284_ _00216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05216_ cpu.IE cpu.needs_interrupt _00699_ _00731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06196_ net29 _01676_ _01580_ _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05147_ cpu.startup_cycle\[3\] cpu.startup_cycle\[2\] _00664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_12_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05348__I cpu.PORTB_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09955_ _04052_ _04904_ _04912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05078_ _00571_ _00598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09886_ _02501_ _04861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08906_ _02643_ _03989_ _03992_ _00410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08837_ _03933_ _03861_ _03934_ _03938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_56_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06355__A2 _01742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08768_ _03864_ _03881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_68_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08699_ cpu.timer_div_counter\[0\] cpu.timer_div_counter\[1\] cpu.timer_div_counter\[2\]
+ _03829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_67_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07304__A1 _01256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_0_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07719_ _01359_ _03035_ _03037_ _00178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10661_ _00555_ clknet_leaf_71_wb_clk_i net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_36_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10592_ _00486_ clknet_leaf_95_wb_clk_i cpu.PC\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_97_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09080__I1 _02789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06043__A1 _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput52 net52 io_oeb[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput41 net41 io_oeb[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput74 net74 io_out[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput63 net63 io_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput85 net85 sram_addr[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput96 net96 sram_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10026_ _02451_ _04968_ _02454_ _02465_ _04969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_clkbuf_leaf_20_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07394__I1 _02093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05721__I _01199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07648__I _02013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06050_ _01530_ _00923_ _01532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_117_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09068__C _04124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07584__S _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09740_ _04222_ _04742_ _00494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06952_ _02423_ _02424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07782__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
.ends

