magic
tech gf180mcuD
magscale 1 10
timestamp 1753968227
<< metal1 >>
rect 30650 47966 30662 48018
rect 30714 48015 30726 48018
rect 31826 48015 31838 48018
rect 30714 47969 31838 48015
rect 30714 47966 30726 47969
rect 31826 47966 31838 47969
rect 31890 47966 31902 48018
rect 43362 47966 43374 48018
rect 43426 48015 43438 48018
rect 43810 48015 43822 48018
rect 43426 47969 43822 48015
rect 43426 47966 43438 47969
rect 43810 47966 43822 47969
rect 43874 47966 43886 48018
rect 1344 47850 49616 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 49616 47850
rect 1344 47764 49616 47798
rect 14366 47682 14418 47694
rect 14366 47618 14418 47630
rect 19014 47570 19066 47582
rect 30662 47570 30714 47582
rect 38838 47570 38890 47582
rect 14802 47518 14814 47570
rect 14866 47518 14878 47570
rect 22418 47518 22430 47570
rect 22482 47518 22494 47570
rect 32610 47518 32622 47570
rect 32674 47518 32686 47570
rect 35970 47518 35982 47570
rect 36034 47518 36046 47570
rect 19014 47506 19066 47518
rect 30662 47506 30714 47518
rect 38838 47506 38890 47518
rect 39286 47570 39338 47582
rect 46386 47518 46398 47570
rect 46450 47518 46462 47570
rect 39286 47506 39338 47518
rect 11790 47458 11842 47470
rect 11790 47394 11842 47406
rect 13246 47458 13298 47470
rect 19182 47458 19234 47470
rect 26238 47458 26290 47470
rect 13246 47394 13298 47406
rect 14110 47350 14122 47402
rect 14174 47350 14186 47402
rect 14914 47391 14926 47443
rect 14978 47391 14990 47443
rect 15138 47406 15150 47458
rect 15202 47406 15214 47458
rect 21186 47406 21198 47458
rect 21250 47406 21262 47458
rect 22754 47406 22766 47458
rect 22818 47406 22830 47458
rect 23090 47406 23102 47458
rect 23154 47406 23166 47458
rect 19182 47394 19234 47406
rect 22586 47350 22598 47402
rect 22650 47350 22662 47402
rect 24658 47362 24670 47414
rect 24722 47362 24734 47414
rect 24882 47406 24894 47458
rect 24946 47406 24958 47458
rect 26238 47394 26290 47406
rect 26350 47458 26402 47470
rect 28366 47458 28418 47470
rect 30830 47458 30882 47470
rect 37326 47458 37378 47470
rect 26618 47406 26630 47458
rect 26682 47406 26694 47458
rect 29230 47406 29242 47458
rect 29294 47406 29306 47458
rect 32162 47406 32174 47458
rect 32226 47406 32238 47458
rect 26350 47394 26402 47406
rect 28366 47394 28418 47406
rect 30830 47394 30882 47406
rect 32498 47362 32510 47414
rect 32562 47362 32574 47414
rect 35186 47378 35198 47430
rect 35250 47378 35262 47430
rect 36082 47362 36094 47414
rect 36146 47362 36158 47414
rect 36306 47406 36318 47458
rect 36370 47406 36382 47458
rect 37326 47394 37378 47406
rect 38278 47458 38330 47470
rect 38278 47394 38330 47406
rect 39678 47458 39730 47470
rect 47294 47458 47346 47470
rect 49310 47458 49362 47470
rect 40450 47406 40462 47458
rect 40514 47406 40526 47458
rect 42802 47406 42814 47458
rect 42866 47406 42878 47458
rect 43810 47406 43822 47458
rect 43874 47406 43886 47458
rect 39678 47394 39730 47406
rect 45826 47378 45838 47430
rect 45890 47378 45902 47430
rect 46498 47362 46510 47414
rect 46562 47362 46574 47414
rect 46722 47406 46734 47458
rect 46786 47406 46798 47458
rect 47954 47406 47966 47458
rect 48018 47406 48030 47458
rect 47294 47394 47346 47406
rect 49310 47394 49362 47406
rect 29486 47346 29538 47358
rect 11454 47234 11506 47246
rect 11454 47170 11506 47182
rect 19518 47234 19570 47246
rect 19518 47170 19570 47182
rect 20918 47234 20970 47246
rect 20918 47170 20970 47182
rect 21366 47234 21418 47246
rect 21366 47170 21418 47182
rect 21926 47234 21978 47246
rect 21926 47170 21978 47182
rect 23270 47234 23322 47246
rect 24770 47238 24782 47290
rect 24834 47238 24846 47290
rect 29486 47282 29538 47294
rect 42366 47346 42418 47358
rect 42366 47282 42418 47294
rect 42982 47290 43034 47302
rect 23270 47170 23322 47182
rect 30214 47234 30266 47246
rect 30214 47170 30266 47182
rect 31166 47234 31218 47246
rect 31166 47170 31218 47182
rect 33742 47234 33794 47246
rect 33742 47170 33794 47182
rect 36934 47234 36986 47246
rect 36934 47170 36986 47182
rect 37662 47234 37714 47246
rect 42982 47226 43034 47238
rect 47630 47234 47682 47246
rect 37662 47170 37714 47182
rect 47630 47170 47682 47182
rect 48134 47234 48186 47246
rect 48134 47170 48186 47182
rect 48974 47234 49026 47246
rect 48974 47170 49026 47182
rect 1344 47066 49616 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 49616 47066
rect 1344 46980 49616 47014
rect 40238 46842 40290 46854
rect 22878 46786 22930 46798
rect 22878 46722 22930 46734
rect 23438 46786 23490 46798
rect 23438 46722 23490 46734
rect 25342 46786 25394 46798
rect 40238 46778 40290 46790
rect 25342 46722 25394 46734
rect 10222 46674 10274 46686
rect 13358 46674 13410 46686
rect 10994 46622 11006 46674
rect 11058 46622 11070 46674
rect 10222 46610 10274 46622
rect 13358 46610 13410 46622
rect 13470 46674 13522 46686
rect 13470 46610 13522 46622
rect 14030 46674 14082 46686
rect 19966 46674 20018 46686
rect 14802 46622 14814 46674
rect 14866 46622 14878 46674
rect 17602 46622 17614 46674
rect 17666 46622 17678 46674
rect 14030 46610 14082 46622
rect 19966 46610 20018 46622
rect 20190 46674 20242 46686
rect 24558 46674 24610 46686
rect 20962 46622 20974 46674
rect 21026 46622 21038 46674
rect 23669 46622 23681 46674
rect 23733 46622 23745 46674
rect 25573 46653 25585 46705
rect 25637 46653 25649 46705
rect 31446 46703 31498 46715
rect 26462 46674 26514 46686
rect 20190 46610 20242 46622
rect 24558 46610 24610 46622
rect 26462 46610 26514 46622
rect 27582 46674 27634 46686
rect 27582 46610 27634 46622
rect 30270 46674 30322 46686
rect 30270 46610 30322 46622
rect 30382 46674 30434 46686
rect 30382 46610 30434 46622
rect 30606 46674 30658 46686
rect 32062 46674 32114 46686
rect 36318 46674 36370 46686
rect 31446 46639 31498 46651
rect 31714 46622 31726 46674
rect 31778 46622 31790 46674
rect 32946 46622 32958 46674
rect 33010 46622 33022 46674
rect 35522 46622 35534 46674
rect 35586 46622 35598 46674
rect 30606 46610 30658 46622
rect 32062 46610 32114 46622
rect 36318 46610 36370 46622
rect 39342 46674 39394 46686
rect 40002 46622 40014 46674
rect 40066 46622 40078 46674
rect 40226 46637 40238 46689
rect 40290 46637 40302 46689
rect 41470 46674 41522 46686
rect 41738 46678 41750 46730
rect 41802 46678 41814 46730
rect 41918 46674 41970 46686
rect 45278 46674 45330 46686
rect 41570 46622 41582 46674
rect 41634 46622 41646 46674
rect 44482 46622 44494 46674
rect 44546 46622 44558 46674
rect 39342 46610 39394 46622
rect 41470 46610 41522 46622
rect 41918 46610 41970 46622
rect 45278 46610 45330 46622
rect 45390 46674 45442 46686
rect 45390 46610 45442 46622
rect 48638 46674 48690 46686
rect 48638 46610 48690 46622
rect 48974 46562 49026 46574
rect 12898 46510 12910 46562
rect 12962 46510 12974 46562
rect 16706 46510 16718 46562
rect 16770 46510 16782 46562
rect 29474 46510 29486 46562
rect 29538 46510 29550 46562
rect 31266 46510 31278 46562
rect 31330 46510 31342 46562
rect 33618 46510 33630 46562
rect 33682 46510 33694 46562
rect 36642 46510 36654 46562
rect 36706 46510 36718 46562
rect 38546 46510 38558 46562
rect 38610 46510 38622 46562
rect 42578 46510 42590 46562
rect 42642 46510 42654 46562
rect 46162 46510 46174 46562
rect 46226 46510 46238 46562
rect 48066 46510 48078 46562
rect 48130 46510 48142 46562
rect 48974 46498 49026 46510
rect 17446 46450 17498 46462
rect 13738 46398 13750 46450
rect 13802 46398 13814 46450
rect 17446 46386 17498 46398
rect 19630 46450 19682 46462
rect 32398 46450 32450 46462
rect 30874 46398 30886 46450
rect 30938 46398 30950 46450
rect 19630 46386 19682 46398
rect 32398 46386 32450 46398
rect 33126 46450 33178 46462
rect 33126 46386 33178 46398
rect 41190 46450 41242 46462
rect 41190 46386 41242 46398
rect 1344 46282 49616 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 49616 46282
rect 1344 46196 49616 46230
rect 43822 46114 43874 46126
rect 40350 46058 40402 46070
rect 43822 46050 43874 46062
rect 11442 45950 11454 46002
rect 11506 45950 11518 46002
rect 18722 45950 18734 46002
rect 18786 45950 18798 46002
rect 22642 45950 22654 46002
rect 22706 45950 22718 46002
rect 24434 45950 24446 46002
rect 24498 45950 24510 46002
rect 29586 45950 29598 46002
rect 29650 45950 29662 46002
rect 30818 45950 30830 46002
rect 30882 45950 30894 46002
rect 37650 45950 37662 46002
rect 37714 45950 37726 46002
rect 40350 45994 40402 46006
rect 41346 45950 41358 46002
rect 41410 45950 41422 46002
rect 12014 45890 12066 45902
rect 14702 45890 14754 45902
rect 9538 45838 9550 45890
rect 9602 45838 9614 45890
rect 11106 45838 11118 45890
rect 11170 45838 11182 45890
rect 11330 45794 11342 45846
rect 11394 45794 11406 45846
rect 12014 45826 12066 45838
rect 12338 45811 12350 45863
rect 12402 45811 12414 45863
rect 12562 45838 12574 45890
rect 12626 45838 12638 45890
rect 13582 45778 13634 45790
rect 13813 45782 13825 45834
rect 13877 45782 13889 45834
rect 14702 45826 14754 45838
rect 14926 45890 14978 45902
rect 17950 45890 18002 45902
rect 15698 45838 15710 45890
rect 15762 45838 15774 45890
rect 14926 45826 14978 45838
rect 17950 45826 18002 45838
rect 21310 45890 21362 45902
rect 23662 45890 23714 45902
rect 21310 45826 21362 45838
rect 22754 45794 22766 45846
rect 22818 45794 22830 45846
rect 23090 45838 23102 45890
rect 23154 45838 23166 45890
rect 23662 45826 23714 45838
rect 26350 45890 26402 45902
rect 26350 45826 26402 45838
rect 27694 45890 27746 45902
rect 28646 45890 28698 45902
rect 30046 45890 30098 45902
rect 27794 45838 27806 45890
rect 27858 45838 27870 45890
rect 29138 45838 29150 45890
rect 29202 45838 29214 45890
rect 29430 45860 29482 45872
rect 27694 45826 27746 45838
rect 28646 45826 28698 45838
rect 36878 45890 36930 45902
rect 41806 45890 41858 45902
rect 30046 45826 30098 45838
rect 33506 45810 33518 45862
rect 33570 45810 33582 45862
rect 40450 45838 40462 45890
rect 40514 45838 40526 45890
rect 40786 45838 40798 45890
rect 40850 45838 40862 45890
rect 41234 45838 41246 45890
rect 41298 45838 41310 45890
rect 36878 45826 36930 45838
rect 41458 45811 41470 45863
rect 41522 45811 41534 45863
rect 41806 45826 41858 45838
rect 42142 45890 42194 45902
rect 42142 45826 42194 45838
rect 42702 45890 42754 45902
rect 45950 45890 46002 45902
rect 45042 45838 45054 45890
rect 45106 45838 45118 45890
rect 45266 45838 45278 45890
rect 45330 45838 45342 45890
rect 42702 45826 42754 45838
rect 29430 45796 29482 45808
rect 12114 45670 12126 45722
rect 12178 45670 12190 45722
rect 13582 45714 13634 45726
rect 17614 45778 17666 45790
rect 17614 45714 17666 45726
rect 20638 45778 20690 45790
rect 20638 45714 20690 45726
rect 32734 45778 32786 45790
rect 32734 45714 32786 45726
rect 39566 45778 39618 45790
rect 43566 45782 43578 45834
rect 43630 45782 43642 45834
rect 45602 45782 45614 45834
rect 45666 45782 45678 45834
rect 45950 45826 46002 45838
rect 46398 45890 46450 45902
rect 47170 45838 47182 45890
rect 47234 45838 47246 45890
rect 46398 45826 46450 45838
rect 39566 45714 39618 45726
rect 49086 45778 49138 45790
rect 27358 45666 27410 45678
rect 27358 45602 27410 45614
rect 27974 45666 28026 45678
rect 27974 45602 28026 45614
rect 36486 45666 36538 45678
rect 36486 45602 36538 45614
rect 44886 45666 44938 45678
rect 46050 45670 46062 45722
rect 46114 45670 46126 45722
rect 49086 45714 49138 45726
rect 44886 45602 44938 45614
rect 1344 45498 49616 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 49616 45498
rect 1344 45412 49616 45446
rect 38894 45330 38946 45342
rect 12126 45218 12178 45230
rect 30706 45222 30718 45274
rect 30770 45222 30782 45274
rect 38894 45266 38946 45278
rect 39958 45330 40010 45342
rect 39958 45266 40010 45278
rect 40406 45330 40458 45342
rect 40406 45266 40458 45278
rect 12126 45154 12178 45166
rect 37494 45218 37546 45230
rect 47506 45222 47518 45274
rect 47570 45222 47582 45274
rect 13694 45145 13746 45157
rect 9438 45106 9490 45118
rect 9438 45042 9490 45054
rect 13470 45106 13522 45118
rect 13694 45081 13746 45093
rect 14018 45054 14030 45106
rect 14082 45054 14094 45106
rect 14578 45098 14590 45150
rect 14642 45098 14654 45150
rect 14802 45054 14814 45106
rect 14866 45054 14878 45106
rect 15362 45054 15374 45106
rect 15426 45054 15438 45106
rect 15586 45098 15598 45150
rect 15650 45098 15662 45150
rect 31054 45145 31106 45157
rect 17726 45106 17778 45118
rect 16930 45054 16942 45106
rect 16994 45054 17006 45106
rect 13470 45042 13522 45054
rect 17726 45042 17778 45054
rect 17838 45106 17890 45118
rect 17838 45042 17890 45054
rect 18398 45106 18450 45118
rect 18398 45042 18450 45054
rect 21534 45106 21586 45118
rect 22306 45054 22318 45106
rect 22370 45054 22382 45106
rect 25218 45054 25230 45106
rect 25282 45054 25294 45106
rect 25554 45069 25566 45121
rect 25618 45069 25630 45121
rect 25902 45106 25954 45118
rect 26674 45054 26686 45106
rect 26738 45054 26750 45106
rect 30594 45054 30606 45106
rect 30658 45054 30670 45106
rect 36206 45141 36258 45153
rect 31054 45081 31106 45093
rect 31278 45106 31330 45118
rect 21534 45042 21586 45054
rect 25902 45042 25954 45054
rect 31278 45042 31330 45054
rect 31726 45106 31778 45118
rect 31726 45042 31778 45054
rect 31950 45106 32002 45118
rect 32958 45106 33010 45118
rect 32218 45054 32230 45106
rect 32282 45054 32294 45106
rect 33730 45054 33742 45106
rect 33794 45054 33806 45106
rect 36306 45110 36318 45162
rect 36370 45110 36382 45162
rect 36542 45134 36594 45146
rect 36206 45077 36258 45089
rect 36754 45110 36766 45162
rect 36818 45110 36830 45162
rect 37494 45154 37546 45166
rect 38334 45162 38386 45174
rect 37774 45134 37826 45146
rect 36542 45070 36594 45082
rect 37046 45106 37098 45118
rect 37774 45070 37826 45082
rect 37998 45134 38050 45146
rect 38210 45110 38222 45162
rect 38274 45110 38286 45162
rect 45726 45141 45778 45153
rect 38334 45098 38386 45110
rect 38558 45106 38610 45118
rect 37998 45070 38050 45082
rect 31950 45042 32002 45054
rect 32958 45042 33010 45054
rect 37046 45042 37098 45054
rect 38558 45042 38610 45054
rect 40910 45106 40962 45118
rect 41774 45054 41786 45106
rect 41838 45054 41850 45106
rect 42690 45054 42702 45106
rect 42754 45054 42766 45106
rect 43250 45081 43262 45133
rect 43314 45081 43326 45133
rect 45826 45110 45838 45162
rect 45890 45110 45902 45162
rect 46062 45134 46114 45146
rect 45726 45077 45778 45089
rect 46274 45110 46286 45162
rect 46338 45110 46350 45162
rect 47742 45145 47794 45157
rect 46062 45070 46114 45082
rect 47282 45054 47294 45106
rect 47346 45054 47358 45106
rect 47742 45081 47794 45093
rect 47966 45106 48018 45118
rect 40910 45042 40962 45054
rect 47966 45042 48018 45054
rect 48638 45106 48690 45118
rect 48638 45042 48690 45054
rect 48862 45106 48914 45118
rect 49130 45054 49142 45106
rect 49194 45054 49206 45106
rect 48862 45042 48914 45054
rect 12742 44994 12794 45006
rect 29542 44994 29594 45006
rect 39510 44994 39562 45006
rect 10210 44942 10222 44994
rect 10274 44942 10286 44994
rect 13906 44942 13918 44994
rect 13970 44942 13982 44994
rect 14466 44942 14478 44994
rect 14530 44942 14542 44994
rect 15698 44942 15710 44994
rect 15762 44942 15774 44994
rect 19170 44942 19182 44994
rect 19234 44942 19246 44994
rect 21074 44942 21086 44994
rect 21138 44942 21150 44994
rect 24210 44942 24222 44994
rect 24274 44942 24286 44994
rect 25666 44942 25678 44994
rect 25730 44942 25742 44994
rect 28578 44942 28590 44994
rect 28642 44942 28654 44994
rect 35634 44942 35646 44994
rect 35698 44942 35710 44994
rect 12742 44930 12794 44942
rect 29542 44930 29594 44942
rect 39510 44930 39562 44942
rect 16774 44882 16826 44894
rect 42030 44882 42082 44894
rect 17434 44830 17446 44882
rect 17498 44830 17510 44882
rect 16774 44818 16826 44830
rect 42030 44818 42082 44830
rect 42534 44882 42586 44894
rect 42534 44818 42586 44830
rect 46566 44882 46618 44894
rect 46566 44818 46618 44830
rect 1344 44714 49616 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 49616 44714
rect 1344 44628 49616 44662
rect 9102 44546 9154 44558
rect 9102 44482 9154 44494
rect 19070 44546 19122 44558
rect 34638 44546 34690 44558
rect 19070 44482 19122 44494
rect 30606 44490 30658 44502
rect 24782 44434 24834 44446
rect 7410 44382 7422 44434
rect 7474 44382 7486 44434
rect 12450 44382 12462 44434
rect 12514 44382 12526 44434
rect 15810 44382 15822 44434
rect 15874 44382 15886 44434
rect 24782 44370 24834 44382
rect 28534 44434 28586 44446
rect 34638 44482 34690 44494
rect 37998 44546 38050 44558
rect 43486 44546 43538 44558
rect 42522 44494 42534 44546
rect 42586 44494 42598 44546
rect 37998 44482 38050 44494
rect 43486 44482 43538 44494
rect 44046 44546 44098 44558
rect 44046 44482 44098 44494
rect 44830 44490 44882 44502
rect 45658 44494 45670 44546
rect 45722 44494 45734 44546
rect 30606 44426 30658 44438
rect 35758 44434 35810 44446
rect 28534 44370 28586 44382
rect 36978 44382 36990 44434
rect 37042 44382 37054 44434
rect 40450 44382 40462 44434
rect 40514 44382 40526 44434
rect 41458 44382 41470 44434
rect 41522 44382 41534 44434
rect 44830 44426 44882 44438
rect 46386 44382 46398 44434
rect 46450 44382 46462 44434
rect 47730 44382 47742 44434
rect 47794 44382 47806 44434
rect 35758 44370 35810 44382
rect 9438 44322 9490 44334
rect 17054 44322 17106 44334
rect 7522 44226 7534 44278
rect 7586 44226 7598 44278
rect 7858 44270 7870 44322
rect 7922 44270 7934 44322
rect 9874 44270 9886 44322
rect 9938 44270 9950 44322
rect 9438 44258 9490 44270
rect 12114 44242 12126 44294
rect 12178 44242 12190 44294
rect 12562 44226 12574 44278
rect 12626 44226 12638 44278
rect 12898 44270 12910 44322
rect 12962 44270 12974 44322
rect 13346 44270 13358 44322
rect 13410 44270 13422 44322
rect 13794 44270 13806 44322
rect 13858 44270 13870 44322
rect 14914 44270 14926 44322
rect 14978 44270 14990 44322
rect 15922 44226 15934 44278
rect 15986 44226 15998 44278
rect 16146 44270 16158 44322
rect 16210 44270 16222 44322
rect 19406 44322 19458 44334
rect 17054 44258 17106 44270
rect 17614 44294 17666 44306
rect 17614 44230 17666 44242
rect 17838 44294 17890 44306
rect 17838 44230 17890 44242
rect 18062 44294 18114 44306
rect 18218 44254 18230 44306
rect 18282 44254 18294 44306
rect 19406 44258 19458 44270
rect 19686 44322 19738 44334
rect 23438 44322 23490 44334
rect 19686 44258 19738 44270
rect 19966 44294 20018 44306
rect 18062 44230 18114 44242
rect 20526 44287 20578 44299
rect 19966 44230 20018 44242
rect 17334 44210 17386 44222
rect 20178 44214 20190 44266
rect 20242 44214 20254 44266
rect 20402 44214 20414 44266
rect 20466 44214 20478 44266
rect 21746 44242 21758 44294
rect 21810 44242 21822 44294
rect 23438 44258 23490 44270
rect 24446 44322 24498 44334
rect 29038 44322 29090 44334
rect 24994 44270 25006 44322
rect 25058 44270 25070 44322
rect 28030 44294 28082 44306
rect 24446 44258 24498 44270
rect 27694 44266 27746 44278
rect 20526 44223 20578 44235
rect 24658 44214 24670 44266
rect 24722 44214 24734 44266
rect 27794 44214 27806 44266
rect 27858 44214 27870 44266
rect 28030 44230 28082 44242
rect 28254 44294 28306 44306
rect 29038 44258 29090 44270
rect 29262 44322 29314 44334
rect 32622 44322 32674 44334
rect 29530 44270 29542 44322
rect 29594 44270 29606 44322
rect 30146 44270 30158 44322
rect 30210 44270 30222 44322
rect 30482 44270 30494 44322
rect 30546 44270 30558 44322
rect 31154 44270 31166 44322
rect 31218 44270 31230 44322
rect 31726 44294 31778 44306
rect 29262 44258 29314 44270
rect 31390 44266 31442 44278
rect 28254 44230 28306 44242
rect 27694 44202 27746 44214
rect 31390 44202 31442 44214
rect 31558 44266 31610 44278
rect 31726 44230 31778 44242
rect 32006 44287 32058 44299
rect 32622 44258 32674 44270
rect 32734 44322 32786 44334
rect 32734 44258 32786 44270
rect 33518 44322 33570 44334
rect 37662 44322 37714 44334
rect 34382 44270 34394 44322
rect 34446 44270 34458 44322
rect 35198 44284 35250 44296
rect 33518 44258 33570 44270
rect 32006 44223 32058 44235
rect 35522 44270 35534 44322
rect 35586 44270 35598 44322
rect 31558 44202 31610 44214
rect 32230 44210 32282 44222
rect 35198 44220 35250 44232
rect 35926 44266 35978 44278
rect 36082 44270 36094 44322
rect 36146 44270 36158 44322
rect 37090 44226 37102 44278
rect 37154 44226 37166 44278
rect 37314 44270 37326 44322
rect 37378 44270 37390 44322
rect 37662 44258 37714 44270
rect 41246 44322 41298 44334
rect 42814 44322 42866 44334
rect 41794 44270 41806 44322
rect 41858 44270 41870 44322
rect 41246 44258 41298 44270
rect 17334 44146 17386 44158
rect 33002 44158 33014 44210
rect 33066 44158 33078 44210
rect 35926 44202 35978 44214
rect 38558 44210 38610 44222
rect 41626 44214 41638 44266
rect 41690 44214 41702 44266
rect 42814 44258 42866 44270
rect 42926 44322 42978 44334
rect 42926 44258 42978 44270
rect 43150 44322 43202 44334
rect 43150 44258 43202 44270
rect 44382 44322 44434 44334
rect 45950 44322 46002 44334
rect 44930 44270 44942 44322
rect 44994 44270 45006 44322
rect 45266 44270 45278 44322
rect 45330 44270 45342 44322
rect 44382 44258 44434 44270
rect 45950 44258 46002 44270
rect 46062 44322 46114 44334
rect 46062 44258 46114 44270
rect 46498 44255 46510 44307
rect 46562 44255 46574 44307
rect 46834 44270 46846 44322
rect 46898 44270 46910 44322
rect 47282 44270 47294 44322
rect 47346 44270 47358 44322
rect 47618 44255 47630 44307
rect 47682 44255 47694 44307
rect 48290 44270 48302 44322
rect 48354 44270 48366 44322
rect 32230 44146 32282 44158
rect 38558 44146 38610 44158
rect 13526 44098 13578 44110
rect 13526 44034 13578 44046
rect 13974 44098 14026 44110
rect 13974 44034 14026 44046
rect 16718 44098 16770 44110
rect 16718 44034 16770 44046
rect 18678 44098 18730 44110
rect 18678 44034 18730 44046
rect 27414 44098 27466 44110
rect 27414 44034 27466 44046
rect 30998 44098 31050 44110
rect 30998 44034 31050 44046
rect 36262 44098 36314 44110
rect 36262 44034 36314 44046
rect 1344 43930 49616 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 49616 43930
rect 1344 43844 49616 43878
rect 43094 43706 43146 43718
rect 11330 43654 11342 43706
rect 11394 43654 11406 43706
rect 21970 43654 21982 43706
rect 22034 43654 22046 43706
rect 22766 43650 22818 43662
rect 19910 43594 19962 43606
rect 6190 43538 6242 43550
rect 9998 43538 10050 43550
rect 6962 43486 6974 43538
rect 7026 43486 7038 43538
rect 10546 43486 10558 43538
rect 10610 43486 10622 43538
rect 10770 43530 10782 43582
rect 10834 43530 10846 43582
rect 11666 43542 11678 43594
rect 11730 43542 11742 43594
rect 11902 43538 11954 43550
rect 11330 43486 11342 43538
rect 11394 43486 11406 43538
rect 6190 43474 6242 43486
rect 9998 43474 10050 43486
rect 11902 43474 11954 43486
rect 12798 43538 12850 43550
rect 12798 43474 12850 43486
rect 12910 43538 12962 43550
rect 12910 43474 12962 43486
rect 13694 43538 13746 43550
rect 13694 43474 13746 43486
rect 13806 43538 13858 43550
rect 13806 43474 13858 43486
rect 14030 43538 14082 43550
rect 16718 43538 16770 43550
rect 14802 43486 14814 43538
rect 14866 43486 14878 43538
rect 14030 43474 14082 43486
rect 16718 43474 16770 43486
rect 17278 43538 17330 43550
rect 17278 43474 17330 43486
rect 17502 43538 17554 43550
rect 19406 43538 19458 43550
rect 18162 43486 18174 43538
rect 18226 43486 18238 43538
rect 18498 43486 18510 43538
rect 18562 43486 18574 43538
rect 20601 43594 20653 43606
rect 19910 43530 19962 43542
rect 20190 43566 20242 43578
rect 20190 43502 20242 43514
rect 20414 43566 20466 43578
rect 21858 43542 21870 43594
rect 21922 43542 21934 43594
rect 22766 43586 22818 43598
rect 28422 43650 28474 43662
rect 20601 43530 20653 43542
rect 22094 43538 22146 43550
rect 22997 43542 23009 43594
rect 23061 43542 23073 43594
rect 20414 43502 20466 43514
rect 21522 43486 21534 43538
rect 21586 43486 21598 43538
rect 17502 43474 17554 43486
rect 19406 43474 19458 43486
rect 22094 43474 22146 43486
rect 23886 43538 23938 43550
rect 24378 43542 24390 43594
rect 24442 43542 24454 43594
rect 28422 43586 28474 43598
rect 33406 43650 33458 43662
rect 43094 43642 43146 43654
rect 25230 43538 25282 43550
rect 28690 43542 28702 43594
rect 28754 43542 28766 43594
rect 28926 43566 28978 43578
rect 24546 43486 24558 43538
rect 24610 43486 24622 43538
rect 28926 43502 28978 43514
rect 29150 43566 29202 43578
rect 29150 43502 29202 43514
rect 29262 43573 29314 43585
rect 29262 43509 29314 43521
rect 29822 43538 29874 43550
rect 30270 43538 30322 43550
rect 23886 43474 23938 43486
rect 25230 43474 25282 43486
rect 29822 43474 29874 43486
rect 29990 43482 30042 43494
rect 30146 43486 30158 43538
rect 30210 43486 30222 43538
rect 19686 43426 19738 43438
rect 8866 43374 8878 43426
rect 8930 43374 8942 43426
rect 10882 43374 10894 43426
rect 10946 43374 10958 43426
rect 9662 43314 9714 43326
rect 18386 43318 18398 43370
rect 18450 43318 18462 43370
rect 19686 43362 19738 43374
rect 21030 43426 21082 43438
rect 30270 43474 30322 43486
rect 31166 43538 31218 43550
rect 31166 43474 31218 43486
rect 31502 43538 31554 43550
rect 31826 43542 31838 43594
rect 31890 43542 31902 43594
rect 33406 43586 33458 43598
rect 35385 43594 35437 43606
rect 44326 43594 44378 43606
rect 33070 43538 33122 43550
rect 32162 43486 32174 43538
rect 32226 43486 32238 43538
rect 33518 43538 33570 43550
rect 34738 43542 34750 43594
rect 34802 43542 34814 43594
rect 34974 43566 35026 43578
rect 31502 43474 31554 43486
rect 33070 43474 33122 43486
rect 33238 43482 33290 43494
rect 24210 43374 24222 43426
rect 24274 43374 24286 43426
rect 26002 43374 26014 43426
rect 26066 43374 26078 43426
rect 27906 43374 27918 43426
rect 27970 43374 27982 43426
rect 29990 43418 30042 43430
rect 30550 43426 30602 43438
rect 21030 43362 21082 43374
rect 30550 43362 30602 43374
rect 31838 43426 31890 43438
rect 34974 43502 35026 43514
rect 35142 43573 35194 43585
rect 35385 43530 35437 43542
rect 36542 43538 36594 43550
rect 40462 43538 40514 43550
rect 35142 43509 35194 43521
rect 35746 43486 35758 43538
rect 35810 43486 35822 43538
rect 36082 43486 36094 43538
rect 36146 43486 36158 43538
rect 37314 43486 37326 43538
rect 37378 43486 37390 43538
rect 40786 43486 40798 43538
rect 40850 43486 40862 43538
rect 41458 43516 41470 43568
rect 41522 43516 41534 43568
rect 41682 43542 41694 43594
rect 41746 43542 41758 43594
rect 42914 43486 42926 43538
rect 42978 43486 42990 43538
rect 43698 43514 43710 43566
rect 43762 43514 43774 43566
rect 44158 43538 44210 43550
rect 43922 43486 43934 43538
rect 43986 43486 43998 43538
rect 44326 43530 44378 43542
rect 44606 43594 44658 43606
rect 44606 43530 44658 43542
rect 44718 43566 44770 43578
rect 44930 43542 44942 43594
rect 44994 43542 45006 43594
rect 45154 43542 45166 43594
rect 45218 43542 45230 43594
rect 44718 43502 44770 43514
rect 45726 43538 45778 43550
rect 33518 43474 33570 43486
rect 36542 43474 36594 43486
rect 40462 43474 40514 43486
rect 41962 43430 41974 43482
rect 42026 43430 42038 43482
rect 44158 43474 44210 43486
rect 45726 43474 45778 43486
rect 45950 43538 46002 43550
rect 45950 43474 46002 43486
rect 47294 43538 47346 43550
rect 47506 43486 47518 43538
rect 47570 43486 47582 43538
rect 47842 43501 47854 43553
rect 47906 43501 47918 43553
rect 48638 43538 48690 43550
rect 47294 43474 47346 43486
rect 48638 43474 48690 43486
rect 33238 43418 33290 43430
rect 31838 43362 31890 43374
rect 35646 43370 35698 43382
rect 39218 43374 39230 43426
rect 39282 43374 39294 43426
rect 19070 43314 19122 43326
rect 12506 43262 12518 43314
rect 12570 43262 12582 43314
rect 13402 43262 13414 43314
rect 13466 43262 13478 43314
rect 17770 43262 17782 43314
rect 17834 43262 17846 43314
rect 9662 43250 9714 43262
rect 19070 43250 19122 43262
rect 33798 43314 33850 43326
rect 33798 43250 33850 43262
rect 34470 43314 34522 43326
rect 40966 43370 41018 43382
rect 47954 43374 47966 43426
rect 48018 43374 48030 43426
rect 35646 43306 35698 43318
rect 40126 43314 40178 43326
rect 34470 43250 34522 43262
rect 40966 43306 41018 43318
rect 42254 43314 42306 43326
rect 40126 43250 40178 43262
rect 42254 43250 42306 43262
rect 45446 43314 45498 43326
rect 46958 43314 47010 43326
rect 46218 43262 46230 43314
rect 46282 43262 46294 43314
rect 45446 43250 45498 43262
rect 46958 43250 47010 43262
rect 48974 43314 49026 43326
rect 48974 43250 49026 43262
rect 1344 43146 49616 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 49616 43146
rect 1344 43060 49616 43094
rect 7198 42978 7250 42990
rect 7198 42914 7250 42926
rect 14590 42978 14642 42990
rect 14590 42914 14642 42926
rect 16046 42978 16098 42990
rect 16046 42914 16098 42926
rect 25454 42978 25506 42990
rect 37830 42978 37882 42990
rect 29530 42926 29542 42978
rect 29594 42926 29606 42978
rect 30314 42926 30326 42978
rect 30378 42926 30390 42978
rect 25454 42914 25506 42926
rect 37830 42914 37882 42926
rect 38446 42978 38498 42990
rect 38446 42914 38498 42926
rect 42030 42978 42082 42990
rect 42030 42914 42082 42926
rect 44102 42978 44154 42990
rect 44102 42914 44154 42926
rect 18722 42814 18734 42866
rect 18786 42814 18798 42866
rect 32790 42810 32842 42822
rect 35298 42814 35310 42866
rect 35362 42814 35374 42866
rect 47170 42814 47182 42866
rect 47234 42814 47246 42866
rect 8318 42754 8370 42766
rect 7429 42702 7441 42754
rect 7493 42702 7505 42754
rect 8318 42690 8370 42702
rect 8766 42754 8818 42766
rect 12238 42754 12290 42766
rect 13470 42754 13522 42766
rect 17950 42754 18002 42766
rect 21646 42754 21698 42766
rect 25790 42754 25842 42766
rect 27414 42754 27466 42766
rect 9538 42702 9550 42754
rect 9602 42702 9614 42754
rect 12898 42702 12910 42754
rect 12962 42702 12974 42754
rect 14334 42702 14346 42754
rect 14398 42702 14410 42754
rect 8766 42690 8818 42702
rect 12238 42690 12290 42702
rect 11454 42642 11506 42654
rect 12562 42646 12574 42698
rect 12626 42646 12638 42698
rect 13470 42690 13522 42702
rect 15362 42674 15374 42726
rect 15426 42674 15438 42726
rect 21186 42702 21198 42754
rect 21250 42702 21262 42754
rect 22418 42702 22430 42754
rect 22482 42702 22494 42754
rect 24770 42702 24782 42754
rect 24834 42702 24846 42754
rect 25890 42702 25902 42754
rect 25954 42702 25966 42754
rect 29038 42754 29090 42766
rect 17950 42690 18002 42702
rect 21646 42690 21698 42702
rect 25790 42690 25842 42702
rect 27414 42690 27466 42702
rect 27694 42726 27746 42738
rect 27694 42662 27746 42674
rect 27918 42726 27970 42738
rect 27918 42662 27970 42674
rect 28142 42726 28194 42738
rect 28142 42662 28194 42674
rect 28254 42698 28306 42710
rect 11454 42578 11506 42590
rect 20638 42642 20690 42654
rect 12114 42534 12126 42586
rect 12178 42534 12190 42586
rect 20638 42578 20690 42590
rect 24334 42642 24386 42654
rect 29038 42690 29090 42702
rect 29262 42754 29314 42766
rect 29262 42690 29314 42702
rect 29822 42754 29874 42766
rect 29822 42690 29874 42702
rect 30046 42754 30098 42766
rect 30046 42690 30098 42702
rect 31166 42754 31218 42766
rect 32510 42754 32562 42766
rect 31166 42690 31218 42702
rect 31390 42715 31442 42727
rect 31826 42702 31838 42754
rect 31890 42702 31902 42754
rect 32790 42746 32842 42758
rect 32958 42754 33010 42766
rect 32510 42690 32562 42702
rect 32958 42690 33010 42702
rect 34078 42754 34130 42766
rect 35982 42754 36034 42766
rect 34078 42690 34130 42702
rect 35030 42698 35082 42710
rect 31390 42651 31442 42663
rect 28254 42634 28306 42646
rect 32230 42642 32282 42654
rect 24334 42578 24386 42590
rect 24950 42586 25002 42598
rect 21366 42530 21418 42542
rect 31266 42534 31278 42586
rect 31330 42534 31342 42586
rect 32230 42578 32282 42590
rect 32622 42642 32674 42654
rect 34514 42646 34526 42698
rect 34578 42646 34590 42698
rect 34738 42646 34750 42698
rect 34802 42646 34814 42698
rect 35410 42687 35422 42739
rect 35474 42687 35486 42739
rect 35634 42702 35646 42754
rect 35698 42702 35710 42754
rect 38110 42754 38162 42766
rect 37102 42726 37154 42738
rect 35982 42690 36034 42702
rect 36990 42698 37042 42710
rect 35030 42634 35082 42646
rect 37550 42726 37602 42738
rect 37102 42662 37154 42674
rect 37314 42646 37326 42698
rect 37378 42646 37390 42698
rect 38110 42690 38162 42702
rect 38782 42754 38834 42766
rect 38782 42690 38834 42702
rect 39790 42754 39842 42766
rect 40910 42754 40962 42766
rect 42366 42754 42418 42766
rect 40338 42702 40350 42754
rect 40402 42702 40414 42754
rect 41774 42702 41786 42754
rect 41838 42702 41850 42754
rect 39790 42690 39842 42702
rect 40910 42690 40962 42702
rect 42366 42690 42418 42702
rect 42590 42754 42642 42766
rect 42590 42690 42642 42702
rect 43374 42754 43426 42766
rect 43374 42690 43426 42702
rect 43822 42754 43874 42766
rect 37550 42662 37602 42674
rect 43530 42646 43542 42698
rect 43594 42646 43606 42698
rect 43822 42690 43874 42702
rect 45166 42754 45218 42766
rect 46398 42754 46450 42766
rect 45166 42690 45218 42702
rect 45390 42715 45442 42727
rect 45714 42702 45726 42754
rect 45778 42702 45790 42754
rect 46398 42690 46450 42702
rect 36990 42634 37042 42646
rect 43710 42642 43762 42654
rect 45390 42651 45442 42663
rect 42858 42590 42870 42642
rect 42922 42590 42934 42642
rect 32622 42578 32674 42590
rect 24950 42522 25002 42534
rect 36318 42530 36370 42542
rect 21366 42466 21418 42478
rect 36318 42466 36370 42478
rect 39118 42530 39170 42542
rect 40450 42534 40462 42586
rect 40514 42534 40526 42586
rect 43710 42578 43762 42590
rect 49086 42642 49138 42654
rect 45602 42534 45614 42586
rect 45666 42534 45678 42586
rect 49086 42578 49138 42590
rect 39118 42466 39170 42478
rect 1344 42362 49616 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 49616 42362
rect 1344 42276 49616 42310
rect 9998 42194 10050 42206
rect 9998 42130 10050 42142
rect 34694 42194 34746 42206
rect 11218 42086 11230 42138
rect 11282 42086 11294 42138
rect 34694 42130 34746 42142
rect 18958 42082 19010 42094
rect 13582 42026 13634 42038
rect 5854 41970 5906 41982
rect 5854 41906 5906 41918
rect 6414 41970 6466 41982
rect 6414 41906 6466 41918
rect 6638 41970 6690 41982
rect 7198 41970 7250 41982
rect 6906 41918 6918 41970
rect 6970 41918 6982 41970
rect 6638 41906 6690 41918
rect 7198 41906 7250 41918
rect 7422 41970 7474 41982
rect 7746 41933 7758 41985
rect 7810 41933 7822 41985
rect 8878 41970 8930 41982
rect 8082 41918 8094 41970
rect 8146 41918 8158 41970
rect 7422 41906 7474 41918
rect 8878 41906 8930 41918
rect 9102 41970 9154 41982
rect 9102 41906 9154 41918
rect 10334 41970 10386 41982
rect 11554 41974 11566 42026
rect 11618 41974 11630 42026
rect 11790 41970 11842 41982
rect 10882 41918 10894 41970
rect 10946 41918 10958 41970
rect 11218 41918 11230 41970
rect 11282 41918 11294 41970
rect 12334 41956 12346 42008
rect 12398 41956 12410 42008
rect 13010 41918 13022 41970
rect 13074 41918 13086 41970
rect 13582 41962 13634 41974
rect 13694 41998 13746 42010
rect 13694 41934 13746 41946
rect 13918 41998 13970 42010
rect 14130 41974 14142 42026
rect 14194 41974 14206 42026
rect 15598 42005 15650 42017
rect 13918 41934 13970 41946
rect 15598 41941 15650 41953
rect 15710 41998 15762 42010
rect 15710 41934 15762 41946
rect 15934 41998 15986 42010
rect 16146 41974 16158 42026
rect 16210 41974 16222 42026
rect 17390 42005 17442 42017
rect 15934 41934 15986 41946
rect 16438 41970 16490 41982
rect 17490 41974 17502 42026
rect 17554 41974 17566 42026
rect 17714 41974 17726 42026
rect 17778 41974 17790 42026
rect 17938 41974 17950 42026
rect 18002 41974 18014 42026
rect 18958 42018 19010 42030
rect 19798 42082 19850 42094
rect 29542 42082 29594 42094
rect 19798 42018 19850 42030
rect 20246 42026 20298 42038
rect 17390 41941 17442 41953
rect 18622 41970 18674 41982
rect 10334 41906 10386 41918
rect 11790 41906 11842 41918
rect 16438 41906 16490 41918
rect 19070 41970 19122 41982
rect 20066 41974 20078 42026
rect 20130 41974 20142 42026
rect 20713 42026 20765 42038
rect 22250 42030 22262 42082
rect 22314 42030 22326 42082
rect 18622 41906 18674 41918
rect 18790 41914 18842 41926
rect 20246 41962 20298 41974
rect 20526 41998 20578 42010
rect 29542 42018 29594 42030
rect 35590 42082 35642 42094
rect 35590 42018 35642 42030
rect 42030 42082 42082 42094
rect 29766 42005 29818 42017
rect 20713 41962 20765 41974
rect 21646 41970 21698 41982
rect 20526 41934 20578 41946
rect 19070 41906 19122 41918
rect 21646 41906 21698 41918
rect 21982 41970 22034 41982
rect 21982 41906 22034 41918
rect 22542 41970 22594 41982
rect 22542 41906 22594 41918
rect 22766 41970 22818 41982
rect 26462 41970 26514 41982
rect 23762 41918 23774 41970
rect 23826 41918 23838 41970
rect 25218 41918 25230 41970
rect 25282 41918 25294 41970
rect 28466 41945 28478 41997
rect 28530 41945 28542 41997
rect 29766 41941 29818 41953
rect 30046 41998 30098 42010
rect 30046 41934 30098 41946
rect 30270 41998 30322 42010
rect 35870 41998 35922 42010
rect 30270 41934 30322 41946
rect 30426 41934 30438 41986
rect 30490 41934 30502 41986
rect 31502 41970 31554 41982
rect 30706 41918 30718 41970
rect 30770 41918 30782 41970
rect 31042 41918 31054 41970
rect 31106 41918 31118 41970
rect 22766 41906 22818 41918
rect 26462 41906 26514 41918
rect 31502 41906 31554 41918
rect 31726 41970 31778 41982
rect 31726 41906 31778 41918
rect 33742 41970 33794 41982
rect 34850 41918 34862 41970
rect 34914 41918 34926 41970
rect 36082 41974 36094 42026
rect 36146 41974 36158 42026
rect 36306 41974 36318 42026
rect 36370 41974 36382 42026
rect 36430 42005 36482 42017
rect 35870 41934 35922 41946
rect 36430 41941 36482 41953
rect 36654 41970 36706 41982
rect 39678 41970 39730 41982
rect 37426 41918 37438 41970
rect 37490 41918 37502 41970
rect 33742 41906 33794 41918
rect 36654 41906 36706 41918
rect 39678 41906 39730 41918
rect 40910 41970 40962 41982
rect 41774 41974 41786 42026
rect 41838 41974 41850 42026
rect 42030 42018 42082 42030
rect 40910 41906 40962 41918
rect 42478 41970 42530 41982
rect 42478 41906 42530 41918
rect 42590 41970 42642 41982
rect 43486 41970 43538 41982
rect 42858 41918 42870 41970
rect 42922 41918 42934 41970
rect 42590 41906 42642 41918
rect 43486 41906 43538 41918
rect 43822 41970 43874 41982
rect 44034 41974 44046 42026
rect 44098 41974 44110 42026
rect 44482 41918 44494 41970
rect 44546 41918 44558 41970
rect 44706 41918 44718 41970
rect 44770 41918 44782 41970
rect 45154 41918 45166 41970
rect 45218 41918 45230 41970
rect 45826 41945 45838 41997
rect 45890 41945 45902 41997
rect 48638 41970 48690 41982
rect 47954 41918 47966 41970
rect 48018 41918 48030 41970
rect 43822 41906 43874 41918
rect 48638 41906 48690 41918
rect 7634 41806 7646 41858
rect 7698 41806 7710 41858
rect 18790 41850 18842 41862
rect 21142 41858 21194 41870
rect 10726 41802 10778 41814
rect 5518 41746 5570 41758
rect 12786 41750 12798 41802
rect 12850 41750 12862 41802
rect 21142 41794 21194 41806
rect 28982 41858 29034 41870
rect 28982 41794 29034 41806
rect 35254 41858 35306 41870
rect 39330 41806 39342 41858
rect 39394 41806 39406 41858
rect 44258 41806 44270 41858
rect 44322 41806 44334 41858
rect 6122 41694 6134 41746
rect 6186 41694 6198 41746
rect 8586 41694 8598 41746
rect 8650 41694 8662 41746
rect 10726 41738 10778 41750
rect 14422 41746 14474 41758
rect 5518 41682 5570 41694
rect 14422 41682 14474 41694
rect 18230 41746 18282 41758
rect 18230 41682 18282 41694
rect 19350 41746 19402 41758
rect 19350 41682 19402 41694
rect 23942 41746 23994 41758
rect 23942 41682 23994 41694
rect 25398 41746 25450 41758
rect 30930 41750 30942 41802
rect 30994 41750 31006 41802
rect 35254 41794 35306 41806
rect 34078 41746 34130 41758
rect 31994 41694 32006 41746
rect 32058 41694 32070 41746
rect 25398 41682 25450 41694
rect 34078 41682 34130 41694
rect 40014 41746 40066 41758
rect 40014 41682 40066 41694
rect 44886 41746 44938 41758
rect 44886 41682 44938 41694
rect 45334 41746 45386 41758
rect 45334 41682 45386 41694
rect 48974 41746 49026 41758
rect 48974 41682 49026 41694
rect 1344 41578 49616 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 49616 41578
rect 1344 41492 49616 41526
rect 10614 41410 10666 41422
rect 10222 41354 10274 41366
rect 10614 41346 10666 41358
rect 17502 41410 17554 41422
rect 40462 41410 40514 41422
rect 17502 41346 17554 41358
rect 31390 41354 31442 41366
rect 6290 41246 6302 41298
rect 6354 41246 6366 41298
rect 10222 41290 10274 41302
rect 40462 41346 40514 41358
rect 43094 41410 43146 41422
rect 43094 41346 43146 41358
rect 15474 41246 15486 41298
rect 15538 41246 15550 41298
rect 16034 41246 16046 41298
rect 16098 41246 16110 41298
rect 29530 41246 29542 41298
rect 29594 41246 29606 41298
rect 31390 41290 31442 41302
rect 45502 41298 45554 41310
rect 35186 41246 35198 41298
rect 35250 41246 35262 41298
rect 45502 41234 45554 41246
rect 5518 41186 5570 41198
rect 5518 41122 5570 41134
rect 8542 41186 8594 41198
rect 8542 41122 8594 41134
rect 8766 41186 8818 41198
rect 11678 41186 11730 41198
rect 16830 41186 16882 41198
rect 17110 41186 17162 41198
rect 9874 41134 9886 41186
rect 9938 41134 9950 41186
rect 10098 41134 10110 41186
rect 10162 41134 10174 41186
rect 10434 41134 10446 41186
rect 10498 41134 10510 41186
rect 10882 41134 10894 41186
rect 10946 41134 10958 41186
rect 8766 41122 8818 41134
rect 11678 41122 11730 41134
rect 8206 41074 8258 41086
rect 12542 41078 12554 41130
rect 12606 41078 12618 41130
rect 13458 41101 13470 41153
rect 13522 41101 13534 41153
rect 13794 41101 13806 41153
rect 13858 41101 13870 41153
rect 12798 41074 12850 41086
rect 14298 41078 14310 41130
rect 14362 41078 14374 41130
rect 14552 41094 14564 41146
rect 14616 41094 14628 41146
rect 15026 41134 15038 41186
rect 15090 41134 15102 41186
rect 15362 41090 15374 41142
rect 15426 41090 15438 41142
rect 16146 41119 16158 41171
rect 16210 41119 16222 41171
rect 16482 41134 16494 41186
rect 16546 41134 16558 41186
rect 16930 41134 16942 41186
rect 16994 41134 17006 41186
rect 16830 41122 16882 41134
rect 17110 41122 17162 41134
rect 19966 41186 20018 41198
rect 22878 41186 22930 41198
rect 23774 41186 23826 41198
rect 21858 41134 21870 41186
rect 21922 41134 21934 41186
rect 23538 41134 23550 41186
rect 23602 41134 23614 41186
rect 19966 41122 20018 41134
rect 22878 41122 22930 41134
rect 9034 41022 9046 41074
rect 9098 41022 9110 41074
rect 8206 41010 8258 41022
rect 12798 41010 12850 41022
rect 14702 41074 14754 41086
rect 23202 41078 23214 41130
rect 23266 41078 23278 41130
rect 23774 41122 23826 41134
rect 24446 41186 24498 41198
rect 29038 41186 29090 41198
rect 25218 41134 25230 41186
rect 25282 41134 25294 41186
rect 27918 41158 27970 41170
rect 24446 41122 24498 41134
rect 28478 41130 28530 41142
rect 27918 41094 27970 41106
rect 14702 41010 14754 41022
rect 27134 41074 27186 41086
rect 11062 40962 11114 40974
rect 11062 40898 11114 40910
rect 18118 40962 18170 40974
rect 18118 40898 18170 40910
rect 19630 40962 19682 40974
rect 19630 40898 19682 40910
rect 20358 40962 20410 40974
rect 20358 40898 20410 40910
rect 20806 40962 20858 40974
rect 20806 40898 20858 40910
rect 22374 40962 22426 40974
rect 23426 40966 23438 41018
rect 23490 40966 23502 41018
rect 27134 41010 27186 41022
rect 27638 41074 27690 41086
rect 28130 41078 28142 41130
rect 28194 41078 28206 41130
rect 28354 41078 28366 41130
rect 28418 41078 28430 41130
rect 29038 41122 29090 41134
rect 29262 41186 29314 41198
rect 29262 41122 29314 41134
rect 29822 41186 29874 41198
rect 29822 41122 29874 41134
rect 30046 41186 30098 41198
rect 31614 41186 31666 41198
rect 30930 41134 30942 41186
rect 30994 41134 31006 41186
rect 31266 41134 31278 41186
rect 31330 41134 31342 41186
rect 30046 41122 30098 41134
rect 31614 41122 31666 41134
rect 31838 41186 31890 41198
rect 31838 41122 31890 41134
rect 33294 41186 33346 41198
rect 33294 41122 33346 41134
rect 35982 41186 36034 41198
rect 40126 41186 40178 41198
rect 49310 41186 49362 41198
rect 37650 41134 37662 41186
rect 37714 41134 37726 41186
rect 35982 41122 36034 41134
rect 39890 41106 39902 41158
rect 39954 41106 39966 41158
rect 40126 41122 40178 41134
rect 42254 41151 42306 41163
rect 44370 41134 44382 41186
rect 44434 41134 44446 41186
rect 44930 41134 44942 41186
rect 44994 41134 45006 41186
rect 45154 41134 45166 41186
rect 45218 41134 45230 41186
rect 45714 41134 45726 41186
rect 45778 41134 45790 41186
rect 45938 41134 45950 41186
rect 46002 41134 46014 41186
rect 48514 41134 48526 41186
rect 48578 41134 48590 41186
rect 42254 41087 42306 41099
rect 42354 41078 42366 41130
rect 42418 41078 42430 41130
rect 42578 41078 42590 41130
rect 42642 41078 42654 41130
rect 42802 41078 42814 41130
rect 42866 41078 42878 41130
rect 49310 41122 49362 41134
rect 28478 41066 28530 41078
rect 46622 41074 46674 41086
rect 30314 41022 30326 41074
rect 30378 41022 30390 41074
rect 32106 41022 32118 41074
rect 32170 41022 32182 41074
rect 27638 41010 27690 41022
rect 46622 41010 46674 41022
rect 22374 40898 22426 40910
rect 24110 40962 24162 40974
rect 24110 40898 24162 40910
rect 36486 40962 36538 40974
rect 36486 40898 36538 40910
rect 37158 40962 37210 40974
rect 37158 40898 37210 40910
rect 41078 40962 41130 40974
rect 41078 40898 41130 40910
rect 41526 40962 41578 40974
rect 41526 40898 41578 40910
rect 41974 40962 42026 40974
rect 41974 40898 42026 40910
rect 43878 40962 43930 40974
rect 43878 40898 43930 40910
rect 44214 40962 44266 40974
rect 44214 40898 44266 40910
rect 1344 40794 49616 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 49616 40794
rect 1344 40708 49616 40742
rect 34470 40626 34522 40638
rect 25790 40570 25842 40582
rect 20750 40514 20802 40526
rect 24098 40518 24110 40570
rect 24162 40518 24174 40570
rect 25790 40506 25842 40518
rect 26630 40570 26682 40582
rect 26630 40506 26682 40518
rect 28142 40514 28194 40526
rect 30258 40518 30270 40570
rect 30322 40518 30334 40570
rect 34470 40562 34522 40574
rect 41526 40626 41578 40638
rect 41526 40562 41578 40574
rect 41974 40626 42026 40638
rect 41974 40562 42026 40574
rect 46454 40626 46506 40638
rect 46454 40562 46506 40574
rect 33910 40514 33962 40526
rect 5394 40350 5406 40402
rect 5458 40350 5470 40402
rect 6626 40377 6638 40429
rect 6690 40377 6702 40429
rect 8318 40402 8370 40414
rect 11442 40406 11454 40458
rect 11506 40406 11518 40458
rect 11790 40402 11842 40414
rect 13234 40406 13246 40458
rect 13298 40406 13310 40458
rect 16382 40441 16434 40453
rect 20750 40450 20802 40462
rect 28970 40462 28982 40514
rect 29034 40462 29046 40514
rect 13582 40402 13634 40414
rect 9538 40350 9550 40402
rect 9602 40350 9614 40402
rect 9874 40350 9886 40402
rect 9938 40350 9950 40402
rect 10434 40350 10446 40402
rect 10498 40350 10510 40402
rect 10658 40350 10670 40402
rect 10722 40350 10734 40402
rect 11106 40350 11118 40402
rect 11170 40350 11182 40402
rect 12898 40350 12910 40402
rect 12962 40350 12974 40402
rect 8318 40338 8370 40350
rect 11790 40338 11842 40350
rect 13582 40338 13634 40350
rect 13918 40402 13970 40414
rect 15822 40402 15874 40414
rect 14466 40350 14478 40402
rect 14530 40350 14542 40402
rect 14802 40350 14814 40402
rect 14866 40350 14878 40402
rect 13918 40338 13970 40350
rect 15822 40338 15874 40350
rect 16158 40402 16210 40414
rect 25678 40441 25730 40453
rect 28142 40450 28194 40462
rect 33070 40458 33122 40470
rect 37270 40514 37322 40526
rect 17726 40402 17778 40414
rect 20414 40402 20466 40414
rect 16382 40377 16434 40389
rect 16818 40350 16830 40402
rect 16882 40350 16894 40402
rect 19618 40350 19630 40402
rect 19682 40350 19694 40402
rect 16158 40338 16210 40350
rect 17726 40338 17778 40350
rect 20414 40338 20466 40350
rect 23438 40402 23490 40414
rect 23438 40338 23490 40350
rect 23998 40402 24050 40414
rect 24322 40377 24334 40429
rect 24386 40377 24398 40429
rect 25454 40402 25506 40414
rect 24546 40350 24558 40402
rect 24610 40350 24622 40402
rect 27022 40402 27074 40414
rect 28478 40402 28530 40414
rect 25678 40377 25730 40389
rect 26114 40350 26126 40402
rect 26178 40350 26190 40402
rect 26786 40350 26798 40402
rect 26850 40350 26862 40402
rect 27886 40350 27898 40402
rect 27950 40350 27962 40402
rect 23998 40338 24050 40350
rect 25454 40338 25506 40350
rect 27022 40338 27074 40350
rect 28478 40338 28530 40350
rect 28702 40402 28754 40414
rect 28702 40338 28754 40350
rect 29710 40402 29762 40414
rect 29922 40406 29934 40458
rect 29986 40406 29998 40458
rect 31210 40406 31222 40458
rect 31274 40406 31286 40458
rect 31614 40402 31666 40414
rect 30370 40350 30382 40402
rect 30434 40350 30446 40402
rect 31042 40350 31054 40402
rect 31106 40350 31118 40402
rect 29710 40338 29762 40350
rect 31614 40338 31666 40350
rect 31950 40402 32002 40414
rect 33070 40394 33122 40406
rect 33182 40430 33234 40442
rect 33182 40366 33234 40378
rect 33406 40430 33458 40442
rect 33618 40406 33630 40458
rect 33682 40406 33694 40458
rect 33910 40450 33962 40462
rect 36430 40458 36482 40470
rect 33406 40366 33458 40378
rect 34862 40402 34914 40414
rect 31950 40338 32002 40350
rect 34862 40338 34914 40350
rect 35198 40402 35250 40414
rect 35198 40338 35250 40350
rect 35310 40402 35362 40414
rect 37270 40450 37322 40462
rect 40238 40514 40290 40526
rect 48078 40514 48130 40526
rect 40238 40450 40290 40462
rect 42926 40458 42978 40470
rect 36430 40394 36482 40406
rect 36542 40430 36594 40442
rect 36542 40366 36594 40378
rect 36766 40430 36818 40442
rect 36766 40366 36818 40378
rect 36990 40430 37042 40442
rect 36990 40366 37042 40378
rect 37550 40402 37602 40414
rect 44214 40458 44266 40470
rect 35310 40338 35362 40350
rect 38322 40350 38334 40402
rect 38386 40350 38398 40402
rect 41346 40350 41358 40402
rect 41410 40350 41422 40402
rect 41794 40350 41806 40402
rect 41858 40350 41870 40402
rect 42578 40350 42590 40402
rect 42642 40350 42654 40402
rect 42926 40394 42978 40406
rect 43654 40402 43706 40414
rect 37550 40338 37602 40350
rect 10110 40290 10162 40302
rect 10110 40226 10162 40238
rect 11454 40290 11506 40302
rect 16494 40290 16546 40302
rect 31278 40290 31330 40302
rect 42802 40294 42814 40346
rect 42866 40294 42878 40346
rect 43654 40338 43706 40350
rect 43990 40402 44042 40414
rect 45091 40458 45143 40470
rect 45782 40458 45834 40470
rect 44214 40394 44266 40406
rect 44494 40430 44546 40442
rect 44494 40366 44546 40378
rect 44718 40430 44770 40442
rect 44718 40366 44770 40378
rect 44874 40366 44886 40418
rect 44938 40366 44950 40418
rect 45091 40394 45143 40406
rect 45278 40430 45330 40442
rect 45490 40406 45502 40458
rect 45554 40406 45566 40458
rect 45782 40394 45834 40406
rect 46958 40402 47010 40414
rect 47822 40406 47834 40458
rect 47886 40406 47898 40458
rect 48078 40450 48130 40462
rect 45278 40366 45330 40378
rect 46274 40350 46286 40402
rect 46338 40350 46350 40402
rect 48850 40365 48862 40417
rect 48914 40365 48926 40417
rect 49074 40350 49086 40402
rect 49138 40350 49150 40402
rect 43990 40338 44042 40350
rect 46958 40338 47010 40350
rect 13122 40238 13134 40290
rect 13186 40238 13198 40290
rect 22642 40238 22654 40290
rect 22706 40238 22718 40290
rect 11454 40226 11506 40238
rect 14802 40182 14814 40234
rect 14866 40182 14878 40234
rect 16494 40226 16546 40238
rect 31278 40226 31330 40238
rect 43486 40290 43538 40302
rect 48738 40238 48750 40290
rect 48802 40238 48814 40290
rect 43486 40226 43538 40238
rect 42422 40178 42474 40190
rect 42422 40114 42474 40126
rect 46006 40178 46058 40190
rect 46006 40114 46058 40126
rect 1344 40010 49616 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 49616 40010
rect 1344 39924 49616 39958
rect 17278 39842 17330 39854
rect 8822 39786 8874 39798
rect 17278 39778 17330 39790
rect 19686 39842 19738 39854
rect 25454 39842 25506 39854
rect 24938 39790 24950 39842
rect 25002 39790 25014 39842
rect 19686 39778 19738 39790
rect 25454 39778 25506 39790
rect 29486 39842 29538 39854
rect 37830 39842 37882 39854
rect 29486 39778 29538 39790
rect 31278 39786 31330 39798
rect 5618 39678 5630 39730
rect 5682 39678 5694 39730
rect 8822 39722 8874 39734
rect 11454 39730 11506 39742
rect 11454 39666 11506 39678
rect 16158 39730 16210 39742
rect 16158 39666 16210 39678
rect 24278 39730 24330 39742
rect 24278 39666 24330 39678
rect 26406 39730 26458 39742
rect 30594 39734 30606 39786
rect 30658 39734 30670 39786
rect 37830 39778 37882 39790
rect 44886 39842 44938 39854
rect 44886 39778 44938 39790
rect 31278 39722 31330 39734
rect 32174 39730 32226 39742
rect 47630 39730 47682 39742
rect 26406 39666 26458 39678
rect 27862 39674 27914 39686
rect 6638 39618 6690 39630
rect 8486 39618 8538 39630
rect 10782 39618 10834 39630
rect 14254 39618 14306 39630
rect 15486 39618 15538 39630
rect 15764 39618 15816 39630
rect 5730 39522 5742 39574
rect 5794 39522 5806 39574
rect 5954 39566 5966 39618
rect 6018 39566 6030 39618
rect 6638 39554 6690 39566
rect 6862 39579 6914 39591
rect 7298 39566 7310 39618
rect 7362 39566 7374 39618
rect 7758 39580 7810 39592
rect 6862 39515 6914 39527
rect 7646 39562 7698 39574
rect 8642 39566 8654 39618
rect 8706 39566 8718 39618
rect 9214 39583 9266 39595
rect 8486 39554 8538 39566
rect 7758 39516 7810 39528
rect 9214 39519 9266 39531
rect 9382 39583 9434 39595
rect 9774 39590 9826 39602
rect 9382 39519 9434 39531
rect 7646 39498 7698 39510
rect 8318 39506 8370 39518
rect 9538 39510 9550 39562
rect 9602 39510 9614 39562
rect 10882 39566 10894 39618
rect 10946 39566 10958 39618
rect 12014 39583 12066 39595
rect 10782 39554 10834 39566
rect 9774 39526 9826 39538
rect 6514 39398 6526 39450
rect 6578 39398 6590 39450
rect 8318 39442 8370 39454
rect 10054 39506 10106 39518
rect 11048 39510 11060 39562
rect 11112 39510 11124 39562
rect 12574 39590 12626 39602
rect 12406 39562 12458 39574
rect 12014 39519 12066 39531
rect 12114 39510 12126 39562
rect 12178 39510 12190 39562
rect 14914 39566 14926 39618
rect 14978 39566 14990 39618
rect 15586 39566 15598 39618
rect 15650 39566 15662 39618
rect 14254 39554 14306 39566
rect 12574 39526 12626 39538
rect 12406 39498 12458 39510
rect 12854 39506 12906 39518
rect 14634 39510 14646 39562
rect 14698 39510 14710 39562
rect 15486 39554 15538 39566
rect 15764 39554 15816 39566
rect 16606 39618 16658 39630
rect 18174 39618 18226 39630
rect 16706 39566 16718 39618
rect 16770 39566 16782 39618
rect 16606 39554 16658 39566
rect 16872 39510 16884 39562
rect 16936 39510 16948 39562
rect 18174 39554 18226 39566
rect 19406 39618 19458 39630
rect 23326 39618 23378 39630
rect 19406 39554 19458 39566
rect 19966 39590 20018 39602
rect 20526 39562 20578 39574
rect 19966 39526 20018 39538
rect 10054 39442 10106 39454
rect 12854 39442 12906 39454
rect 19070 39506 19122 39518
rect 20178 39510 20190 39562
rect 20242 39510 20254 39562
rect 20402 39510 20414 39562
rect 20466 39510 20478 39562
rect 21634 39538 21646 39590
rect 21698 39538 21710 39590
rect 23326 39554 23378 39566
rect 24446 39618 24498 39630
rect 24446 39554 24498 39566
rect 24670 39618 24722 39630
rect 24670 39554 24722 39566
rect 25790 39618 25842 39630
rect 25790 39554 25842 39566
rect 27694 39618 27746 39630
rect 35074 39678 35086 39730
rect 35138 39678 35150 39730
rect 38882 39678 38894 39730
rect 38946 39678 38958 39730
rect 40786 39678 40798 39730
rect 40850 39678 40862 39730
rect 46386 39678 46398 39730
rect 46450 39678 46462 39730
rect 32174 39666 32226 39678
rect 47630 39666 47682 39678
rect 48750 39730 48802 39742
rect 48750 39666 48802 39678
rect 48918 39674 48970 39686
rect 27862 39610 27914 39622
rect 28142 39618 28194 39630
rect 27694 39554 27746 39566
rect 28142 39554 28194 39566
rect 28422 39618 28474 39630
rect 28422 39554 28474 39566
rect 29878 39618 29930 39630
rect 30158 39618 30210 39630
rect 32846 39618 32898 39630
rect 35422 39618 35474 39630
rect 30034 39566 30046 39618
rect 30098 39566 30110 39618
rect 30482 39566 30494 39618
rect 30546 39566 30558 39618
rect 30818 39566 30830 39618
rect 30882 39566 30894 39618
rect 31378 39566 31390 39618
rect 31442 39566 31454 39618
rect 31602 39566 31614 39618
rect 31666 39566 31678 39618
rect 32722 39566 32734 39618
rect 32786 39566 32798 39618
rect 34626 39566 34638 39618
rect 34690 39566 34702 39618
rect 29878 39554 29930 39566
rect 30158 39554 30210 39566
rect 20526 39498 20578 39510
rect 28030 39506 28082 39518
rect 32556 39510 32568 39562
rect 32620 39510 32632 39562
rect 32846 39554 32898 39566
rect 34962 39551 34974 39603
rect 35026 39551 35038 39603
rect 38110 39618 38162 39630
rect 43486 39618 43538 39630
rect 45614 39618 45666 39630
rect 35422 39554 35474 39566
rect 36990 39583 37042 39595
rect 37326 39590 37378 39602
rect 36990 39519 37042 39531
rect 37090 39510 37102 39562
rect 37154 39510 37166 39562
rect 42802 39566 42814 39618
rect 42866 39566 42878 39618
rect 45042 39566 45054 39618
rect 45106 39566 45118 39618
rect 37326 39526 37378 39538
rect 37538 39510 37550 39562
rect 37602 39510 37614 39562
rect 38110 39554 38162 39566
rect 43250 39510 43262 39562
rect 43314 39510 43326 39562
rect 43486 39554 43538 39566
rect 45614 39554 45666 39566
rect 45950 39618 46002 39630
rect 46958 39618 47010 39630
rect 46498 39566 46510 39618
rect 46562 39566 46574 39618
rect 47058 39566 47070 39618
rect 47122 39566 47134 39618
rect 48190 39580 48242 39592
rect 45950 39554 46002 39566
rect 46162 39510 46174 39562
rect 46226 39510 46238 39562
rect 46958 39554 47010 39566
rect 47224 39510 47236 39562
rect 47288 39510 47300 39562
rect 48514 39566 48526 39618
rect 48578 39566 48590 39618
rect 48918 39610 48970 39622
rect 48190 39516 48242 39528
rect 14130 39398 14142 39450
rect 14194 39398 14206 39450
rect 19070 39442 19122 39454
rect 28030 39442 28082 39454
rect 18510 39394 18562 39406
rect 18510 39330 18562 39342
rect 33350 39394 33402 39406
rect 33350 39330 33402 39342
rect 33798 39394 33850 39406
rect 33798 39330 33850 39342
rect 34358 39394 34410 39406
rect 34358 39330 34410 39342
rect 35758 39394 35810 39406
rect 35758 39330 35810 39342
rect 36486 39394 36538 39406
rect 36486 39330 36538 39342
rect 41638 39394 41690 39406
rect 41638 39330 41690 39342
rect 42086 39394 42138 39406
rect 42086 39330 42138 39342
rect 42534 39394 42586 39406
rect 43026 39398 43038 39450
rect 43090 39398 43102 39450
rect 42534 39330 42586 39342
rect 44326 39394 44378 39406
rect 44326 39330 44378 39342
rect 1344 39226 49616 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 49616 39226
rect 1344 39140 49616 39174
rect 11790 39058 11842 39070
rect 25454 39058 25506 39070
rect 11790 38994 11842 39006
rect 14646 39002 14698 39014
rect 6526 38946 6578 38958
rect 10446 38946 10498 38958
rect 12562 38950 12574 39002
rect 12626 38950 12638 39002
rect 25454 38994 25506 39006
rect 26126 39058 26178 39070
rect 26126 38994 26178 39006
rect 29262 39058 29314 39070
rect 29262 38994 29314 39006
rect 29934 39058 29986 39070
rect 48974 39058 49026 39070
rect 29934 38994 29986 39006
rect 44606 39002 44658 39014
rect 6526 38882 6578 38894
rect 9494 38890 9546 38902
rect 14646 38938 14698 38950
rect 15710 38946 15762 38958
rect 48974 38994 49026 39006
rect 6190 38834 6242 38846
rect 6757 38838 6769 38890
rect 6821 38838 6833 38890
rect 5394 38782 5406 38834
rect 5458 38782 5470 38834
rect 6190 38770 6242 38782
rect 7646 38834 7698 38846
rect 8878 38834 8930 38846
rect 8586 38782 8598 38834
rect 8650 38782 8662 38834
rect 7646 38770 7698 38782
rect 8878 38770 8930 38782
rect 9102 38834 9154 38846
rect 9650 38838 9662 38890
rect 9714 38838 9726 38890
rect 10446 38882 10498 38894
rect 9494 38826 9546 38838
rect 9874 38821 9886 38873
rect 9938 38821 9950 38873
rect 12126 38834 12178 38846
rect 12898 38838 12910 38890
rect 12962 38838 12974 38890
rect 15710 38882 15762 38894
rect 15878 38890 15930 38902
rect 16426 38894 16438 38946
rect 16490 38894 16502 38946
rect 44606 38938 44658 38950
rect 31222 38890 31274 38902
rect 13134 38834 13186 38846
rect 10994 38782 11006 38834
rect 11058 38782 11070 38834
rect 11330 38782 11342 38834
rect 11394 38782 11406 38834
rect 12450 38782 12462 38834
rect 12514 38782 12526 38834
rect 14802 38782 14814 38834
rect 14866 38782 14878 38834
rect 15250 38810 15262 38862
rect 15314 38810 15326 38862
rect 15474 38782 15486 38834
rect 15538 38782 15550 38834
rect 15878 38826 15930 38838
rect 16718 38834 16770 38846
rect 9102 38770 9154 38782
rect 12126 38770 12178 38782
rect 13134 38770 13186 38782
rect 16718 38770 16770 38782
rect 16942 38834 16994 38846
rect 16942 38770 16994 38782
rect 20638 38834 20690 38846
rect 20962 38826 20974 38878
rect 21026 38826 21038 38878
rect 21298 38782 21310 38834
rect 21362 38782 21374 38834
rect 22082 38782 22094 38834
rect 22146 38782 22158 38834
rect 22306 38797 22318 38849
rect 22370 38797 22382 38849
rect 22922 38838 22934 38890
rect 22986 38838 22998 38890
rect 23090 38782 23102 38834
rect 23154 38782 23166 38834
rect 23874 38797 23886 38849
rect 23938 38797 23950 38849
rect 25118 38834 25170 38846
rect 24210 38782 24222 38834
rect 24274 38782 24286 38834
rect 20638 38770 20690 38782
rect 25118 38770 25170 38782
rect 25790 38834 25842 38846
rect 25790 38770 25842 38782
rect 26462 38834 26514 38846
rect 26462 38770 26514 38782
rect 26686 38834 26738 38846
rect 27246 38834 27298 38846
rect 26954 38782 26966 38834
rect 27018 38782 27030 38834
rect 26686 38770 26738 38782
rect 27246 38770 27298 38782
rect 28814 38834 28866 38846
rect 28814 38770 28866 38782
rect 28926 38834 28978 38846
rect 28926 38770 28978 38782
rect 29598 38834 29650 38846
rect 30650 38838 30662 38890
rect 30714 38838 30726 38890
rect 30818 38782 30830 38834
rect 30882 38782 30894 38834
rect 31222 38826 31274 38838
rect 31614 38890 31666 38902
rect 31714 38838 31726 38890
rect 31778 38838 31790 38890
rect 31938 38838 31950 38890
rect 32002 38838 32014 38890
rect 32174 38862 32226 38874
rect 31614 38826 31666 38838
rect 36766 38869 36818 38881
rect 32174 38798 32226 38810
rect 33182 38834 33234 38846
rect 29598 38770 29650 38782
rect 33182 38770 33234 38782
rect 35870 38834 35922 38846
rect 35870 38770 35922 38782
rect 35982 38834 36034 38846
rect 36866 38838 36878 38890
rect 36930 38838 36942 38890
rect 37090 38838 37102 38890
rect 37154 38838 37166 38890
rect 45576 38871 45628 38883
rect 36766 38805 36818 38817
rect 37352 38798 37364 38850
rect 37416 38798 37428 38850
rect 37606 38834 37658 38846
rect 35982 38770 36034 38782
rect 37606 38770 37658 38782
rect 37998 38834 38050 38846
rect 37998 38770 38050 38782
rect 40798 38834 40850 38846
rect 40798 38770 40850 38782
rect 44270 38834 44322 38846
rect 44594 38809 44606 38861
rect 44658 38809 44670 38861
rect 45278 38834 45330 38846
rect 44818 38782 44830 38834
rect 44882 38782 44894 38834
rect 45378 38782 45390 38834
rect 45442 38782 45454 38834
rect 47070 38869 47122 38881
rect 45576 38807 45628 38819
rect 46846 38834 46898 38846
rect 47070 38805 47122 38817
rect 47238 38869 47290 38881
rect 47238 38805 47290 38817
rect 47406 38862 47458 38874
rect 47406 38798 47458 38810
rect 47680 38862 47732 38874
rect 47680 38798 47732 38810
rect 48638 38834 48690 38846
rect 44270 38770 44322 38782
rect 45278 38770 45330 38782
rect 46846 38770 46898 38782
rect 48638 38770 48690 38782
rect 8262 38722 8314 38734
rect 3490 38670 3502 38722
rect 3554 38670 3566 38722
rect 8262 38658 8314 38670
rect 17558 38722 17610 38734
rect 24726 38722 24778 38734
rect 17938 38670 17950 38722
rect 18002 38670 18014 38722
rect 19842 38670 19854 38722
rect 19906 38670 19918 38722
rect 20850 38670 20862 38722
rect 20914 38670 20926 38722
rect 22418 38670 22430 38722
rect 22482 38670 22494 38722
rect 22754 38670 22766 38722
rect 22818 38670 22830 38722
rect 23762 38670 23774 38722
rect 23826 38670 23838 38722
rect 11106 38614 11118 38666
rect 11170 38614 11182 38666
rect 17558 38658 17610 38670
rect 24726 38658 24778 38670
rect 27582 38722 27634 38734
rect 27582 38658 27634 38670
rect 28478 38722 28530 38734
rect 28478 38658 28530 38670
rect 31054 38722 31106 38734
rect 31054 38658 31106 38670
rect 32454 38722 32506 38734
rect 38950 38722 39002 38734
rect 45950 38722 46002 38734
rect 35074 38670 35086 38722
rect 35138 38670 35150 38722
rect 41570 38670 41582 38722
rect 41634 38670 41646 38722
rect 43474 38670 43486 38722
rect 43538 38670 43550 38722
rect 32454 38658 32506 38670
rect 38950 38658 39002 38670
rect 45950 38658 46002 38670
rect 46510 38722 46562 38734
rect 46510 38658 46562 38670
rect 36318 38610 36370 38622
rect 36318 38546 36370 38558
rect 38334 38610 38386 38622
rect 38334 38546 38386 38558
rect 47910 38610 47962 38622
rect 47910 38546 47962 38558
rect 1344 38442 49616 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 49616 38442
rect 1344 38356 49616 38390
rect 11678 38274 11730 38286
rect 10602 38222 10614 38274
rect 10666 38222 10678 38274
rect 11678 38210 11730 38222
rect 16550 38274 16602 38286
rect 30102 38274 30154 38286
rect 31782 38274 31834 38286
rect 16550 38210 16602 38222
rect 23214 38218 23266 38230
rect 9214 38162 9266 38174
rect 30874 38222 30886 38274
rect 30938 38222 30950 38274
rect 30102 38210 30154 38222
rect 31782 38210 31834 38222
rect 33294 38274 33346 38286
rect 45950 38274 46002 38286
rect 34794 38222 34806 38274
rect 34858 38222 34870 38274
rect 33294 38210 33346 38222
rect 45950 38210 46002 38222
rect 8194 38110 8206 38162
rect 8258 38110 8270 38162
rect 18722 38110 18734 38162
rect 18786 38110 18798 38162
rect 21410 38110 21422 38162
rect 21474 38110 21486 38162
rect 23214 38154 23266 38166
rect 24098 38110 24110 38162
rect 24162 38110 24174 38162
rect 26562 38110 26574 38162
rect 26626 38110 26638 38162
rect 28466 38110 28478 38162
rect 28530 38110 28542 38162
rect 38546 38110 38558 38162
rect 38610 38110 38622 38162
rect 40450 38110 40462 38162
rect 40514 38110 40526 38162
rect 41682 38110 41694 38162
rect 41746 38110 41758 38162
rect 43698 38110 43710 38162
rect 43762 38110 43774 38162
rect 46610 38110 46622 38162
rect 46674 38110 46686 38162
rect 48514 38110 48526 38162
rect 48578 38110 48590 38162
rect 9214 38098 9266 38110
rect 5518 38050 5570 38062
rect 10110 38050 10162 38062
rect 6290 37998 6302 38050
rect 6354 37998 6366 38050
rect 8642 37998 8654 38050
rect 8706 37998 8718 38050
rect 8978 37998 8990 38050
rect 9042 37998 9054 38050
rect 9538 37998 9550 38050
rect 9602 37998 9614 38050
rect 9762 37998 9774 38050
rect 9826 37998 9838 38050
rect 5518 37986 5570 37998
rect 10110 37986 10162 37998
rect 10334 38050 10386 38062
rect 10334 37986 10386 37998
rect 12014 38050 12066 38062
rect 12014 37986 12066 37998
rect 12350 38050 12402 38062
rect 12350 37986 12402 37998
rect 12574 38050 12626 38062
rect 12574 37986 12626 37998
rect 13358 38050 13410 38062
rect 16046 38050 16098 38062
rect 18958 38050 19010 38062
rect 14130 37998 14142 38050
rect 14194 37998 14206 38050
rect 13358 37986 13410 37998
rect 16046 37986 16098 37998
rect 16830 38022 16882 38034
rect 16830 37958 16882 37970
rect 16998 38015 17050 38027
rect 17390 38015 17442 38027
rect 16998 37951 17050 37963
rect 17266 37942 17278 37994
rect 17330 37942 17342 37994
rect 17602 37998 17614 38050
rect 17666 37998 17678 38050
rect 18386 37998 18398 38050
rect 18450 37998 18462 38050
rect 17390 37951 17442 37963
rect 18610 37954 18622 38006
rect 18674 37954 18686 38006
rect 18958 37986 19010 37998
rect 19294 38050 19346 38062
rect 19294 37986 19346 37998
rect 20302 38050 20354 38062
rect 20302 37986 20354 37998
rect 20582 38050 20634 38062
rect 20582 37986 20634 37998
rect 20750 38050 20802 38062
rect 21982 38050 22034 38062
rect 21298 37998 21310 38050
rect 21362 37998 21374 38050
rect 20750 37986 20802 37998
rect 20022 37938 20074 37950
rect 12842 37886 12854 37938
rect 12906 37886 12918 37938
rect 20022 37874 20074 37886
rect 20414 37938 20466 37950
rect 21634 37942 21646 37994
rect 21698 37942 21710 37994
rect 21982 37986 22034 37998
rect 22318 38050 22370 38062
rect 24670 38050 24722 38062
rect 23314 37998 23326 38050
rect 23378 37998 23390 38050
rect 23650 37998 23662 38050
rect 23714 37998 23726 38050
rect 23986 37998 23998 38050
rect 24050 37998 24062 38050
rect 24446 38011 24498 38023
rect 22318 37986 22370 37998
rect 24670 37986 24722 37998
rect 25006 38050 25058 38062
rect 25006 37986 25058 37998
rect 25790 38050 25842 38062
rect 30382 38050 30434 38062
rect 25790 37986 25842 37998
rect 29262 38015 29314 38027
rect 24446 37947 24498 37959
rect 29598 38022 29650 38034
rect 29262 37951 29314 37963
rect 29362 37942 29374 37994
rect 29426 37942 29438 37994
rect 29598 37958 29650 37970
rect 29810 37942 29822 37994
rect 29874 37942 29886 37994
rect 30382 37986 30434 37998
rect 30606 38050 30658 38062
rect 32958 38050 33010 38062
rect 30606 37986 30658 37998
rect 31502 37994 31554 38006
rect 31602 37998 31614 38050
rect 31666 37998 31678 38050
rect 32958 37986 33010 37998
rect 35086 38050 35138 38062
rect 35086 37986 35138 37998
rect 35310 38050 35362 38062
rect 36374 38050 36426 38062
rect 35646 38022 35698 38034
rect 35310 37986 35362 37998
rect 35534 37994 35586 38006
rect 31502 37930 31554 37942
rect 35646 37958 35698 37970
rect 35926 38015 35978 38027
rect 35926 37951 35978 37963
rect 36082 37942 36094 37994
rect 36146 37942 36158 37994
rect 36374 37986 36426 37998
rect 36878 38050 36930 38062
rect 36878 37986 36930 37998
rect 37774 38050 37826 38062
rect 42254 38050 42306 38062
rect 43374 38050 43426 38062
rect 44718 38050 44770 38062
rect 41234 37998 41246 38050
rect 41298 37998 41310 38050
rect 37774 37986 37826 37998
rect 41570 37983 41582 38035
rect 41634 37983 41646 38035
rect 42485 37998 42497 38050
rect 42549 37998 42561 38050
rect 42254 37986 42306 37998
rect 43374 37986 43426 37998
rect 43810 37954 43822 38006
rect 43874 37954 43886 38006
rect 44146 37998 44158 38050
rect 44210 37998 44222 38050
rect 44718 37986 44770 37998
rect 44942 38050 44994 38062
rect 44942 37986 44994 37998
rect 46286 38050 46338 38062
rect 46286 37986 46338 37998
rect 49310 38050 49362 38062
rect 49310 37986 49362 37998
rect 35534 37930 35586 37942
rect 20414 37874 20466 37886
rect 31334 37882 31386 37894
rect 45210 37886 45222 37938
rect 45274 37886 45286 37938
rect 17782 37826 17834 37838
rect 31334 37818 31386 37830
rect 32790 37826 32842 37838
rect 17782 37762 17834 37774
rect 32790 37762 32842 37774
rect 33910 37826 33962 37838
rect 33910 37762 33962 37774
rect 34470 37826 34522 37838
rect 34470 37762 34522 37774
rect 37214 37826 37266 37838
rect 37214 37762 37266 37774
rect 1344 37658 49616 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 49616 37658
rect 1344 37572 49616 37606
rect 8598 37490 8650 37502
rect 8598 37426 8650 37438
rect 9606 37490 9658 37502
rect 9606 37426 9658 37438
rect 13582 37490 13634 37502
rect 13582 37426 13634 37438
rect 15822 37490 15874 37502
rect 15822 37426 15874 37438
rect 16774 37490 16826 37502
rect 16774 37426 16826 37438
rect 19126 37490 19178 37502
rect 19126 37426 19178 37438
rect 21086 37490 21138 37502
rect 21086 37426 21138 37438
rect 25734 37490 25786 37502
rect 25734 37426 25786 37438
rect 28310 37490 28362 37502
rect 28310 37426 28362 37438
rect 30998 37490 31050 37502
rect 30998 37426 31050 37438
rect 45110 37490 45162 37502
rect 12910 37378 12962 37390
rect 6234 37270 6246 37322
rect 6298 37270 6310 37322
rect 12910 37314 12962 37326
rect 17502 37378 17554 37390
rect 17502 37314 17554 37326
rect 24222 37378 24274 37390
rect 10222 37266 10274 37278
rect 5954 37214 5966 37266
rect 6018 37214 6030 37266
rect 8418 37214 8430 37266
rect 8482 37214 8494 37266
rect 9762 37214 9774 37266
rect 9826 37214 9838 37266
rect 10222 37202 10274 37214
rect 13246 37266 13298 37278
rect 13246 37202 13298 37214
rect 16158 37266 16210 37278
rect 17733 37270 17745 37322
rect 17797 37270 17809 37322
rect 24222 37314 24274 37326
rect 27134 37378 27186 37390
rect 27134 37314 27186 37326
rect 31894 37378 31946 37390
rect 31894 37314 31946 37326
rect 32398 37378 32450 37390
rect 32398 37314 32450 37326
rect 34414 37378 34466 37390
rect 18622 37266 18674 37278
rect 16930 37214 16942 37266
rect 16994 37214 17006 37266
rect 16158 37202 16210 37214
rect 18622 37202 18674 37214
rect 19854 37266 19906 37278
rect 21422 37266 21474 37278
rect 20178 37214 20190 37266
rect 20242 37214 20254 37266
rect 20514 37214 20526 37266
rect 20578 37214 20590 37266
rect 19854 37202 19906 37214
rect 21422 37202 21474 37214
rect 21534 37266 21586 37278
rect 26014 37266 26066 37278
rect 22306 37214 22318 37266
rect 22370 37214 22382 37266
rect 26878 37214 26890 37266
rect 26942 37214 26954 37266
rect 28578 37214 28590 37266
rect 28642 37214 28654 37266
rect 28914 37229 28926 37281
rect 28978 37229 28990 37281
rect 29262 37266 29314 37278
rect 21534 37202 21586 37214
rect 26014 37202 26066 37214
rect 29262 37202 29314 37214
rect 30158 37266 30210 37278
rect 32062 37266 32114 37278
rect 30818 37214 30830 37266
rect 30882 37214 30894 37266
rect 30158 37202 30210 37214
rect 32062 37202 32114 37214
rect 33294 37266 33346 37278
rect 34158 37270 34170 37322
rect 34222 37270 34234 37322
rect 34414 37314 34466 37326
rect 39118 37378 39170 37390
rect 39118 37314 39170 37326
rect 40406 37378 40458 37390
rect 41682 37382 41694 37434
rect 41746 37382 41758 37434
rect 45110 37426 45162 37438
rect 45950 37490 46002 37502
rect 45950 37426 46002 37438
rect 47058 37382 47070 37434
rect 47122 37382 47134 37434
rect 40406 37314 40458 37326
rect 36430 37266 36482 37278
rect 35746 37214 35758 37266
rect 35810 37214 35822 37266
rect 37202 37214 37214 37266
rect 37266 37214 37278 37266
rect 41010 37214 41022 37266
rect 41074 37214 41086 37266
rect 41234 37241 41246 37293
rect 41298 37241 41310 37293
rect 41582 37266 41634 37278
rect 42354 37214 42366 37266
rect 42418 37214 42430 37266
rect 44258 37241 44270 37293
rect 44322 37241 44334 37293
rect 46286 37266 46338 37278
rect 46778 37270 46790 37322
rect 46842 37270 46854 37322
rect 47182 37266 47234 37278
rect 49310 37266 49362 37278
rect 44930 37214 44942 37266
rect 44994 37214 45006 37266
rect 46610 37214 46622 37266
rect 46674 37214 46686 37266
rect 47730 37214 47742 37266
rect 47794 37214 47806 37266
rect 48066 37214 48078 37266
rect 48130 37214 48142 37266
rect 33294 37202 33346 37214
rect 36430 37202 36482 37214
rect 41582 37202 41634 37214
rect 46286 37202 46338 37214
rect 47182 37202 47234 37214
rect 49310 37202 49362 37214
rect 27750 37154 27802 37166
rect 36150 37154 36202 37166
rect 6402 37102 6414 37154
rect 6466 37102 6478 37154
rect 10994 37102 11006 37154
rect 11058 37102 11070 37154
rect 20078 37098 20130 37110
rect 19518 37042 19570 37054
rect 29026 37102 29038 37154
rect 29090 37102 29102 37154
rect 27750 37090 27802 37102
rect 36150 37090 36202 37102
rect 39734 37154 39786 37166
rect 39734 37090 39786 37102
rect 48190 37098 48242 37110
rect 20078 37034 20130 37046
rect 29598 37042 29650 37054
rect 19518 36978 19570 36990
rect 29598 36978 29650 36990
rect 30494 37042 30546 37054
rect 48190 37034 48242 37046
rect 48974 37042 49026 37054
rect 30494 36978 30546 36990
rect 48974 36978 49026 36990
rect 1344 36874 49616 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 49616 36874
rect 1344 36788 49616 36822
rect 11454 36706 11506 36718
rect 11454 36642 11506 36654
rect 14926 36706 14978 36718
rect 23382 36706 23434 36718
rect 14926 36642 14978 36654
rect 22542 36650 22594 36662
rect 20806 36594 20858 36606
rect 9986 36542 9998 36594
rect 10050 36542 10062 36594
rect 17714 36542 17726 36594
rect 17778 36542 17790 36594
rect 20806 36530 20858 36542
rect 21702 36594 21754 36606
rect 21702 36530 21754 36542
rect 22150 36594 22202 36606
rect 23382 36642 23434 36654
rect 37102 36706 37154 36718
rect 37102 36642 37154 36654
rect 44930 36598 44942 36650
rect 44994 36598 45006 36650
rect 22542 36586 22594 36598
rect 22150 36530 22202 36542
rect 23942 36538 23994 36550
rect 27010 36542 27022 36594
rect 27074 36542 27086 36594
rect 29810 36542 29822 36594
rect 29874 36542 29886 36594
rect 31714 36542 31726 36594
rect 31778 36542 31790 36594
rect 35746 36542 35758 36594
rect 35810 36542 35822 36594
rect 43698 36542 43710 36594
rect 43762 36542 43774 36594
rect 6638 36482 6690 36494
rect 6638 36418 6690 36430
rect 7310 36482 7362 36494
rect 11790 36482 11842 36494
rect 8082 36430 8094 36482
rect 8146 36430 8158 36482
rect 7310 36418 7362 36430
rect 11790 36418 11842 36430
rect 12070 36482 12122 36494
rect 14590 36482 14642 36494
rect 20414 36482 20466 36494
rect 23662 36482 23714 36494
rect 12070 36418 12122 36430
rect 12294 36447 12346 36459
rect 12294 36383 12346 36395
rect 12574 36454 12626 36466
rect 12574 36390 12626 36402
rect 12786 36374 12798 36426
rect 12850 36374 12862 36426
rect 12954 36414 12966 36466
rect 13018 36414 13030 36466
rect 16718 36454 16770 36466
rect 14590 36418 14642 36430
rect 16382 36426 16434 36438
rect 16482 36374 16494 36426
rect 16546 36374 16558 36426
rect 16718 36390 16770 36402
rect 16942 36454 16994 36466
rect 19618 36430 19630 36482
rect 19682 36430 19694 36482
rect 22642 36430 22654 36482
rect 22706 36430 22718 36482
rect 22866 36430 22878 36482
rect 22930 36430 22942 36482
rect 23942 36474 23994 36486
rect 24110 36482 24162 36494
rect 20414 36418 20466 36430
rect 23662 36418 23714 36430
rect 24110 36418 24162 36430
rect 24334 36482 24386 36494
rect 32510 36482 32562 36494
rect 25106 36430 25118 36482
rect 25170 36430 25182 36482
rect 27750 36447 27802 36459
rect 24334 36418 24386 36430
rect 16942 36390 16994 36402
rect 27750 36383 27802 36395
rect 28030 36454 28082 36466
rect 28366 36426 28418 36438
rect 28030 36390 28082 36402
rect 16382 36362 16434 36374
rect 17222 36370 17274 36382
rect 17222 36306 17274 36318
rect 23774 36370 23826 36382
rect 23774 36306 23826 36318
rect 27526 36370 27578 36382
rect 28242 36374 28254 36426
rect 28306 36374 28318 36426
rect 32510 36418 32562 36430
rect 33182 36482 33234 36494
rect 33182 36418 33234 36430
rect 36542 36482 36594 36494
rect 36542 36418 36594 36430
rect 37438 36482 37490 36494
rect 37438 36418 37490 36430
rect 38278 36482 38330 36494
rect 38278 36418 38330 36430
rect 39342 36482 39394 36494
rect 42366 36482 42418 36494
rect 45614 36482 45666 36494
rect 41570 36430 41582 36482
rect 41634 36430 41646 36482
rect 39342 36418 39394 36430
rect 42366 36418 42418 36430
rect 42478 36461 42530 36473
rect 43810 36415 43822 36467
rect 43874 36415 43886 36467
rect 44034 36430 44046 36482
rect 44098 36430 44110 36482
rect 44818 36430 44830 36482
rect 44882 36430 44894 36482
rect 45154 36430 45166 36482
rect 45218 36430 45230 36482
rect 45614 36418 45666 36430
rect 45838 36482 45890 36494
rect 49310 36482 49362 36494
rect 48514 36430 48526 36482
rect 48578 36430 48590 36482
rect 45838 36418 45890 36430
rect 49310 36418 49362 36430
rect 42478 36397 42530 36409
rect 28366 36362 28418 36374
rect 29318 36370 29370 36382
rect 27526 36306 27578 36318
rect 29318 36306 29370 36318
rect 33854 36370 33906 36382
rect 33854 36306 33906 36318
rect 39678 36370 39730 36382
rect 46622 36370 46674 36382
rect 46106 36318 46118 36370
rect 46170 36318 46182 36370
rect 39678 36306 39730 36318
rect 46622 36306 46674 36318
rect 6302 36258 6354 36270
rect 6302 36194 6354 36206
rect 13638 36258 13690 36270
rect 13638 36194 13690 36206
rect 16102 36258 16154 36270
rect 16102 36194 16154 36206
rect 32846 36258 32898 36270
rect 32846 36194 32898 36206
rect 37830 36258 37882 36270
rect 37830 36194 37882 36206
rect 39006 36258 39058 36270
rect 39006 36194 39058 36206
rect 1344 36090 49616 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 49616 36090
rect 1344 36004 49616 36038
rect 8766 35922 8818 35934
rect 8766 35858 8818 35870
rect 18398 35922 18450 35934
rect 18398 35858 18450 35870
rect 19182 35922 19234 35934
rect 19182 35858 19234 35870
rect 24166 35922 24218 35934
rect 24166 35858 24218 35870
rect 25790 35922 25842 35934
rect 25790 35858 25842 35870
rect 31222 35922 31274 35934
rect 31222 35858 31274 35870
rect 31614 35922 31666 35934
rect 31614 35858 31666 35870
rect 35422 35922 35474 35934
rect 35422 35858 35474 35870
rect 39622 35922 39674 35934
rect 42366 35922 42418 35934
rect 39622 35858 39674 35870
rect 40238 35866 40290 35878
rect 7870 35810 7922 35822
rect 7870 35746 7922 35758
rect 16158 35810 16210 35822
rect 5182 35698 5234 35710
rect 9102 35698 9154 35710
rect 5954 35646 5966 35698
rect 6018 35646 6030 35698
rect 5182 35634 5234 35646
rect 9102 35634 9154 35646
rect 9606 35698 9658 35710
rect 9874 35702 9886 35754
rect 9938 35702 9950 35754
rect 10110 35726 10162 35738
rect 10110 35662 10162 35674
rect 10334 35726 10386 35738
rect 10334 35662 10386 35674
rect 10490 35662 10502 35714
rect 10554 35662 10566 35714
rect 12226 35702 12238 35754
rect 12290 35702 12302 35754
rect 12450 35702 12462 35754
rect 12514 35702 12526 35754
rect 12674 35702 12686 35754
rect 12738 35702 12750 35754
rect 16158 35746 16210 35758
rect 21198 35810 21250 35822
rect 30102 35810 30154 35822
rect 21198 35746 21250 35758
rect 27694 35754 27746 35766
rect 41010 35814 41022 35866
rect 41074 35814 41086 35866
rect 42366 35858 42418 35870
rect 40238 35802 40290 35814
rect 12798 35733 12850 35745
rect 27134 35726 27186 35738
rect 12798 35669 12850 35681
rect 13470 35698 13522 35710
rect 18734 35698 18786 35710
rect 9606 35634 9658 35646
rect 14242 35646 14254 35698
rect 14306 35646 14318 35698
rect 17490 35646 17502 35698
rect 17554 35646 17566 35698
rect 17714 35646 17726 35698
rect 17778 35646 17790 35698
rect 13470 35634 13522 35646
rect 18734 35634 18786 35646
rect 18846 35698 18898 35710
rect 20806 35698 20858 35710
rect 20066 35646 20078 35698
rect 20130 35646 20142 35698
rect 20290 35646 20302 35698
rect 20354 35646 20366 35698
rect 18846 35634 18898 35646
rect 20806 35634 20858 35646
rect 21086 35698 21138 35710
rect 21534 35698 21586 35710
rect 21086 35634 21138 35646
rect 21366 35642 21418 35654
rect 10950 35586 11002 35598
rect 10950 35522 11002 35534
rect 16886 35586 16938 35598
rect 21534 35634 21586 35646
rect 22766 35698 22818 35710
rect 25398 35698 25450 35710
rect 23426 35646 23438 35698
rect 23490 35646 23502 35698
rect 22766 35634 22818 35646
rect 25398 35634 25450 35646
rect 26126 35698 26178 35710
rect 27346 35702 27358 35754
rect 27410 35702 27422 35754
rect 27582 35726 27634 35738
rect 27134 35662 27186 35674
rect 29262 35733 29314 35745
rect 27694 35690 27746 35702
rect 29038 35698 29090 35710
rect 27582 35662 27634 35674
rect 26126 35634 26178 35646
rect 29262 35669 29314 35681
rect 29374 35726 29426 35738
rect 29586 35702 29598 35754
rect 29650 35702 29662 35754
rect 29810 35702 29822 35754
rect 29874 35702 29886 35754
rect 30102 35746 30154 35758
rect 29374 35662 29426 35674
rect 31950 35698 32002 35710
rect 29038 35634 29090 35646
rect 31950 35634 32002 35646
rect 32062 35698 32114 35710
rect 34414 35698 34466 35710
rect 33170 35646 33182 35698
rect 33234 35646 33246 35698
rect 33506 35646 33518 35698
rect 33570 35646 33582 35698
rect 37090 35673 37102 35725
rect 37154 35673 37166 35725
rect 37326 35698 37378 35710
rect 32062 35634 32114 35646
rect 34414 35634 34466 35646
rect 37326 35634 37378 35646
rect 38558 35698 38610 35710
rect 38558 35634 38610 35646
rect 39230 35698 39282 35710
rect 39890 35646 39902 35698
rect 39954 35646 39966 35698
rect 40226 35661 40238 35713
rect 40290 35661 40302 35713
rect 41010 35646 41022 35698
rect 41074 35646 41086 35698
rect 41234 35673 41246 35725
rect 41298 35673 41310 35725
rect 42030 35698 42082 35710
rect 39230 35634 39282 35646
rect 21366 35578 21418 35590
rect 22374 35586 22426 35598
rect 16886 35522 16938 35534
rect 17838 35530 17890 35542
rect 11958 35474 12010 35486
rect 20178 35478 20190 35530
rect 20242 35478 20254 35530
rect 22374 35522 22426 35534
rect 23102 35586 23154 35598
rect 23102 35522 23154 35534
rect 24614 35586 24666 35598
rect 24614 35522 24666 35534
rect 26518 35586 26570 35598
rect 26518 35522 26570 35534
rect 28198 35586 28250 35598
rect 28198 35522 28250 35534
rect 30662 35586 30714 35598
rect 30662 35522 30714 35534
rect 37662 35586 37714 35598
rect 41570 35590 41582 35642
rect 41634 35590 41646 35642
rect 42030 35634 42082 35646
rect 42702 35698 42754 35710
rect 43474 35646 43486 35698
rect 43538 35646 43550 35698
rect 45826 35646 45838 35698
rect 45890 35646 45902 35698
rect 46162 35673 46174 35725
rect 46226 35673 46238 35725
rect 46510 35698 46562 35710
rect 42702 35634 42754 35646
rect 46510 35634 46562 35646
rect 46846 35698 46898 35710
rect 47506 35661 47518 35713
rect 47570 35661 47582 35713
rect 47730 35646 47742 35698
rect 47794 35646 47806 35698
rect 48850 35690 48862 35742
rect 48914 35690 48926 35742
rect 49074 35646 49086 35698
rect 49138 35646 49150 35698
rect 46846 35634 46898 35646
rect 45378 35534 45390 35586
rect 45442 35534 45454 35586
rect 45938 35534 45950 35586
rect 46002 35534 46014 35586
rect 47394 35534 47406 35586
rect 47458 35534 47470 35586
rect 48738 35534 48750 35586
rect 48802 35534 48814 35586
rect 17838 35466 17890 35478
rect 26854 35474 26906 35486
rect 11958 35410 12010 35422
rect 26854 35410 26906 35422
rect 28702 35474 28754 35486
rect 28702 35410 28754 35422
rect 32398 35474 32450 35486
rect 33282 35478 33294 35530
rect 33346 35478 33358 35530
rect 37662 35522 37714 35534
rect 32398 35410 32450 35422
rect 34078 35474 34130 35486
rect 34078 35410 34130 35422
rect 38222 35474 38274 35486
rect 38222 35410 38274 35422
rect 38894 35474 38946 35486
rect 38894 35410 38946 35422
rect 1344 35306 49616 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 49616 35306
rect 1344 35220 49616 35254
rect 14422 35138 14474 35150
rect 43598 35138 43650 35150
rect 14422 35074 14474 35086
rect 35646 35082 35698 35094
rect 34078 35026 34130 35038
rect 7410 34974 7422 35026
rect 7474 34974 7486 35026
rect 23426 34974 23438 35026
rect 23490 34974 23502 35026
rect 28466 34974 28478 35026
rect 28530 34974 28542 35026
rect 35646 35018 35698 35030
rect 37774 35082 37826 35094
rect 43598 35074 43650 35086
rect 44886 35138 44938 35150
rect 44886 35074 44938 35086
rect 35970 34974 35982 35026
rect 36034 34974 36046 35026
rect 37774 35018 37826 35030
rect 38770 34974 38782 35026
rect 38834 34974 38846 35026
rect 47170 34974 47182 35026
rect 47234 34974 47246 35026
rect 6190 34914 6242 34926
rect 4834 34862 4846 34914
rect 4898 34862 4910 34914
rect 10110 34914 10162 34926
rect 20862 34914 20914 34926
rect 6190 34850 6242 34862
rect 6626 34834 6638 34886
rect 6690 34834 6702 34886
rect 10882 34862 10894 34914
rect 10946 34862 10958 34914
rect 14646 34879 14698 34891
rect 10110 34850 10162 34862
rect 14646 34815 14698 34827
rect 14926 34886 14978 34898
rect 14926 34822 14978 34834
rect 15150 34886 15202 34898
rect 15150 34822 15202 34834
rect 15262 34858 15314 34870
rect 15810 34862 15822 34914
rect 15874 34862 15886 34914
rect 17490 34862 17502 34914
rect 17554 34862 17566 34914
rect 20066 34862 20078 34914
rect 20130 34862 20142 34914
rect 12798 34802 12850 34814
rect 20862 34850 20914 34862
rect 24222 34914 24274 34926
rect 25790 34914 25842 34926
rect 29038 34914 29090 34926
rect 32734 34914 32786 34926
rect 24222 34850 24274 34862
rect 24446 34858 24498 34870
rect 26562 34862 26574 34914
rect 26626 34862 26638 34914
rect 29810 34862 29822 34914
rect 29874 34862 29886 34914
rect 15262 34794 15314 34806
rect 18174 34802 18226 34814
rect 12798 34738 12850 34750
rect 18174 34738 18226 34750
rect 21534 34802 21586 34814
rect 24546 34806 24558 34858
rect 24610 34806 24622 34858
rect 24770 34806 24782 34858
rect 24834 34806 24846 34858
rect 24994 34806 25006 34858
rect 25058 34806 25070 34858
rect 25790 34850 25842 34862
rect 29038 34850 29090 34862
rect 32734 34850 32786 34862
rect 32958 34914 33010 34926
rect 32958 34850 33010 34862
rect 33406 34914 33458 34926
rect 33730 34918 33742 34970
rect 33794 34918 33806 34970
rect 34078 34962 34130 34974
rect 34918 34914 34970 34926
rect 37998 34914 38050 34926
rect 34290 34862 34302 34914
rect 34354 34862 34366 34914
rect 35186 34862 35198 34914
rect 35250 34862 35262 34914
rect 35522 34862 35534 34914
rect 35586 34862 35598 34914
rect 33406 34850 33458 34862
rect 24446 34794 24498 34806
rect 25286 34802 25338 34814
rect 21534 34738 21586 34750
rect 25286 34738 25338 34750
rect 31726 34802 31778 34814
rect 34066 34806 34078 34858
rect 34130 34806 34142 34858
rect 34918 34850 34970 34862
rect 36082 34847 36094 34899
rect 36146 34847 36158 34899
rect 36418 34862 36430 34914
rect 36482 34862 36494 34914
rect 36922 34815 36934 34867
rect 36986 34815 36998 34867
rect 37650 34862 37662 34914
rect 37714 34862 37726 34914
rect 37998 34850 38050 34862
rect 40686 34914 40738 34926
rect 40686 34850 40738 34862
rect 41694 34914 41746 34926
rect 43262 34914 43314 34926
rect 42242 34862 42254 34914
rect 42306 34862 42318 34914
rect 42578 34862 42590 34914
rect 42642 34862 42654 34914
rect 41694 34850 41746 34862
rect 42018 34806 42030 34858
rect 42082 34806 42094 34858
rect 43262 34850 43314 34862
rect 45166 34914 45218 34926
rect 45614 34914 45666 34926
rect 45266 34862 45278 34914
rect 45330 34862 45342 34914
rect 46398 34914 46450 34926
rect 45166 34850 45218 34862
rect 45434 34806 45446 34858
rect 45498 34806 45510 34858
rect 45614 34850 45666 34862
rect 46286 34858 46338 34870
rect 46398 34850 46450 34862
rect 32442 34750 32454 34802
rect 32506 34750 32518 34802
rect 46286 34794 46338 34806
rect 49086 34802 49138 34814
rect 31726 34738 31778 34750
rect 42758 34746 42810 34758
rect 5854 34690 5906 34702
rect 5854 34626 5906 34638
rect 9382 34690 9434 34702
rect 9382 34626 9434 34638
rect 9942 34690 9994 34702
rect 9942 34626 9994 34638
rect 15654 34690 15706 34702
rect 15654 34626 15706 34638
rect 16214 34690 16266 34702
rect 16214 34626 16266 34638
rect 16774 34690 16826 34702
rect 16774 34626 16826 34638
rect 17334 34690 17386 34702
rect 17334 34626 17386 34638
rect 17670 34690 17722 34702
rect 42130 34694 42142 34746
rect 42194 34694 42206 34746
rect 49086 34738 49138 34750
rect 42758 34682 42810 34694
rect 44326 34690 44378 34702
rect 17670 34626 17722 34638
rect 44326 34626 44378 34638
rect 46118 34690 46170 34702
rect 46118 34626 46170 34638
rect 1344 34522 49616 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 49616 34522
rect 1344 34436 49616 34470
rect 12238 34354 12290 34366
rect 12238 34290 12290 34302
rect 12854 34354 12906 34366
rect 12854 34290 12906 34302
rect 27246 34354 27298 34366
rect 9606 34242 9658 34254
rect 17502 34242 17554 34254
rect 19842 34246 19854 34298
rect 19906 34246 19918 34298
rect 27246 34290 27298 34302
rect 30270 34354 30322 34366
rect 30270 34290 30322 34302
rect 31670 34354 31722 34366
rect 31670 34290 31722 34302
rect 34974 34354 35026 34366
rect 34974 34290 35026 34302
rect 43094 34354 43146 34366
rect 43094 34290 43146 34302
rect 44158 34354 44210 34366
rect 44158 34290 44210 34302
rect 47966 34354 48018 34366
rect 47966 34290 48018 34302
rect 9606 34178 9658 34190
rect 10446 34186 10498 34198
rect 33742 34242 33794 34254
rect 5518 34130 5570 34142
rect 8206 34130 8258 34142
rect 6290 34078 6302 34130
rect 6354 34078 6366 34130
rect 5518 34066 5570 34078
rect 8206 34066 8258 34078
rect 9102 34130 9154 34142
rect 9874 34134 9886 34186
rect 9938 34134 9950 34186
rect 10110 34158 10162 34170
rect 10110 34094 10162 34106
rect 10334 34158 10386 34170
rect 10446 34122 10498 34134
rect 10838 34130 10890 34142
rect 11106 34134 11118 34186
rect 11170 34134 11182 34186
rect 17502 34178 17554 34190
rect 28814 34186 28866 34198
rect 11286 34165 11338 34177
rect 10334 34094 10386 34106
rect 9102 34066 9154 34078
rect 11286 34101 11338 34113
rect 11566 34158 11618 34170
rect 11566 34094 11618 34106
rect 11678 34165 11730 34177
rect 11678 34101 11730 34113
rect 11902 34130 11954 34142
rect 10838 34066 10890 34078
rect 11902 34066 11954 34078
rect 13022 34130 13074 34142
rect 16370 34078 16382 34130
rect 16434 34078 16446 34130
rect 16706 34122 16718 34174
rect 16770 34122 16782 34174
rect 18622 34130 18674 34142
rect 19294 34130 19346 34142
rect 17733 34078 17745 34130
rect 17797 34078 17809 34130
rect 19002 34078 19014 34130
rect 19066 34078 19078 34130
rect 13022 34066 13074 34078
rect 18622 34066 18674 34078
rect 19294 34066 19346 34078
rect 19518 34130 19570 34142
rect 19730 34078 19742 34130
rect 19794 34078 19806 34130
rect 20066 34122 20078 34174
rect 20130 34122 20142 34174
rect 21086 34169 21138 34181
rect 20626 34078 20638 34130
rect 20690 34078 20702 34130
rect 21086 34105 21138 34117
rect 21310 34130 21362 34142
rect 19518 34066 19570 34078
rect 21310 34066 21362 34078
rect 21646 34130 21698 34142
rect 22194 34105 22206 34157
rect 22258 34105 22270 34157
rect 25118 34130 25170 34142
rect 21646 34066 21698 34078
rect 25118 34066 25170 34078
rect 26518 34130 26570 34142
rect 26518 34066 26570 34078
rect 26910 34130 26962 34142
rect 28914 34134 28926 34186
rect 28978 34134 28990 34186
rect 29138 34134 29150 34186
rect 29202 34134 29214 34186
rect 29362 34134 29374 34186
rect 29426 34134 29438 34186
rect 28814 34122 28866 34134
rect 29654 34130 29706 34142
rect 26910 34066 26962 34078
rect 29654 34066 29706 34078
rect 29934 34130 29986 34142
rect 29934 34066 29986 34078
rect 31278 34130 31330 34142
rect 31278 34066 31330 34078
rect 33406 34130 33458 34142
rect 33562 34134 33574 34186
rect 33626 34134 33638 34186
rect 33742 34178 33794 34190
rect 37998 34242 38050 34254
rect 45502 34242 45554 34254
rect 37998 34178 38050 34190
rect 39062 34186 39114 34198
rect 41066 34190 41078 34242
rect 41130 34190 41142 34242
rect 33406 34066 33458 34078
rect 33854 34130 33906 34142
rect 33854 34066 33906 34078
rect 34638 34130 34690 34142
rect 34638 34066 34690 34078
rect 35310 34130 35362 34142
rect 36082 34078 36094 34130
rect 36146 34078 36158 34130
rect 38546 34108 38558 34160
rect 38610 34108 38622 34160
rect 38882 34134 38894 34186
rect 38946 34134 38958 34186
rect 45222 34186 45274 34198
rect 39062 34122 39114 34134
rect 40238 34130 40290 34142
rect 35310 34066 35362 34078
rect 40238 34066 40290 34078
rect 41358 34130 41410 34142
rect 41358 34066 41410 34078
rect 41582 34130 41634 34142
rect 41906 34122 41918 34174
rect 41970 34122 41982 34174
rect 43654 34130 43706 34142
rect 42130 34078 42142 34130
rect 42194 34078 42206 34130
rect 42466 34078 42478 34130
rect 42530 34078 42542 34130
rect 42914 34078 42926 34130
rect 42978 34078 42990 34130
rect 41582 34066 41634 34078
rect 43654 34066 43706 34078
rect 43822 34130 43874 34142
rect 44706 34108 44718 34160
rect 44770 34108 44782 34160
rect 44930 34117 44942 34169
rect 44994 34117 45006 34169
rect 45502 34178 45554 34190
rect 47294 34242 47346 34254
rect 45222 34122 45274 34134
rect 46174 34130 46226 34142
rect 47038 34134 47050 34186
rect 47102 34134 47114 34186
rect 47294 34178 47346 34190
rect 43822 34066 43874 34078
rect 46174 34066 46226 34078
rect 47630 34130 47682 34142
rect 47630 34066 47682 34078
rect 49310 34130 49362 34142
rect 49310 34066 49362 34078
rect 20974 34018 21026 34030
rect 13794 33966 13806 34018
rect 13858 33966 13870 34018
rect 15698 33966 15710 34018
rect 15762 33966 15774 34018
rect 16818 33966 16830 34018
rect 16882 33966 16894 34018
rect 20974 33954 21026 33966
rect 26070 34018 26122 34030
rect 48974 34018 49026 34030
rect 41794 33966 41806 34018
rect 41858 33966 41870 34018
rect 26070 33954 26122 33966
rect 48974 33954 49026 33966
rect 8766 33906 8818 33918
rect 8766 33842 8818 33854
rect 23214 33906 23266 33918
rect 23214 33842 23266 33854
rect 25454 33906 25506 33918
rect 25454 33842 25506 33854
rect 30942 33906 30994 33918
rect 30942 33842 30994 33854
rect 34134 33906 34186 33918
rect 34134 33842 34186 33854
rect 39342 33906 39394 33918
rect 39342 33842 39394 33854
rect 39902 33906 39954 33918
rect 39902 33842 39954 33854
rect 42646 33906 42698 33918
rect 42646 33842 42698 33854
rect 1344 33738 49616 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 49616 33738
rect 1344 33652 49616 33686
rect 10166 33570 10218 33582
rect 22374 33570 22426 33582
rect 10166 33506 10218 33518
rect 15038 33514 15090 33526
rect 22374 33506 22426 33518
rect 38110 33570 38162 33582
rect 38110 33506 38162 33518
rect 41974 33570 42026 33582
rect 41974 33506 42026 33518
rect 7746 33406 7758 33458
rect 7810 33406 7822 33458
rect 11442 33406 11454 33458
rect 11506 33406 11518 33458
rect 12898 33406 12910 33458
rect 12962 33406 12974 33458
rect 15038 33450 15090 33462
rect 16594 33406 16606 33458
rect 16658 33406 16670 33458
rect 18498 33406 18510 33458
rect 18562 33406 18574 33458
rect 23762 33406 23774 33458
rect 23826 33406 23838 33458
rect 25666 33406 25678 33458
rect 25730 33406 25742 33458
rect 30482 33406 30494 33458
rect 30546 33406 30558 33458
rect 32386 33406 32398 33458
rect 32450 33406 32462 33458
rect 33842 33406 33854 33458
rect 33906 33406 33918 33458
rect 35746 33406 35758 33458
rect 35810 33406 35822 33458
rect 46610 33406 46622 33458
rect 46674 33406 46686 33458
rect 6974 33346 7026 33358
rect 6974 33282 7026 33294
rect 9662 33346 9714 33358
rect 13582 33346 13634 33358
rect 9662 33282 9714 33294
rect 10446 33318 10498 33330
rect 11510 33316 11562 33328
rect 11006 33290 11058 33302
rect 10446 33254 10498 33266
rect 10658 33238 10670 33290
rect 10722 33238 10734 33290
rect 10882 33238 10894 33290
rect 10946 33238 10958 33290
rect 11890 33294 11902 33346
rect 11954 33294 11966 33346
rect 12450 33294 12462 33346
rect 12514 33294 12526 33346
rect 12786 33279 12798 33331
rect 12850 33279 12862 33331
rect 13582 33282 13634 33294
rect 14702 33346 14754 33358
rect 15822 33346 15874 33358
rect 22094 33346 22146 33358
rect 15138 33294 15150 33346
rect 15202 33294 15214 33346
rect 15474 33294 15486 33346
rect 15538 33294 15550 33346
rect 19394 33294 19406 33346
rect 19458 33294 19470 33346
rect 19742 33318 19794 33330
rect 11510 33252 11562 33264
rect 13813 33238 13825 33290
rect 13877 33238 13889 33290
rect 14702 33282 14754 33294
rect 15822 33282 15874 33294
rect 19630 33290 19682 33302
rect 20190 33318 20242 33330
rect 19742 33254 19794 33266
rect 19954 33238 19966 33290
rect 20018 33238 20030 33290
rect 26462 33346 26514 33358
rect 22094 33282 22146 33294
rect 22654 33318 22706 33330
rect 20190 33254 20242 33266
rect 22654 33254 22706 33266
rect 22878 33318 22930 33330
rect 23214 33311 23266 33323
rect 22878 33254 22930 33266
rect 11006 33226 11058 33238
rect 19630 33226 19682 33238
rect 20470 33234 20522 33246
rect 23090 33238 23102 33290
rect 23154 33238 23166 33290
rect 26462 33282 26514 33294
rect 29710 33346 29762 33358
rect 29710 33282 29762 33294
rect 33070 33346 33122 33358
rect 39678 33346 39730 33358
rect 49310 33346 49362 33358
rect 33070 33282 33122 33294
rect 39442 33266 39454 33318
rect 39506 33266 39518 33318
rect 39678 33282 39730 33294
rect 40518 33290 40570 33302
rect 23214 33247 23266 33259
rect 19238 33178 19290 33190
rect 20470 33170 20522 33182
rect 26854 33234 26906 33246
rect 40674 33238 40686 33290
rect 40738 33238 40750 33290
rect 40898 33255 40910 33307
rect 40962 33255 40974 33307
rect 41794 33294 41806 33346
rect 41858 33294 41870 33346
rect 42590 33311 42642 33323
rect 42590 33247 42642 33259
rect 42758 33311 42810 33323
rect 43150 33318 43202 33330
rect 42758 33247 42810 33259
rect 40518 33226 40570 33238
rect 41470 33234 41522 33246
rect 42914 33238 42926 33290
rect 42978 33238 42990 33290
rect 44034 33294 44046 33346
rect 44098 33294 44110 33346
rect 45726 33290 45778 33302
rect 45938 33294 45950 33346
rect 46002 33294 46014 33346
rect 48514 33294 48526 33346
rect 48578 33294 48590 33346
rect 43150 33254 43202 33266
rect 26854 33170 26906 33182
rect 41470 33170 41522 33182
rect 43430 33234 43482 33246
rect 44886 33234 44938 33246
rect 45154 33238 45166 33290
rect 45218 33238 45230 33290
rect 45378 33238 45390 33290
rect 45442 33238 45454 33290
rect 45602 33238 45614 33290
rect 45666 33238 45678 33290
rect 49310 33282 49362 33294
rect 43430 33170 43482 33182
rect 43878 33178 43930 33190
rect 19238 33114 19290 33126
rect 21758 33122 21810 33134
rect 21758 33058 21810 33070
rect 36374 33122 36426 33134
rect 36374 33058 36426 33070
rect 40014 33122 40066 33134
rect 45726 33226 45778 33238
rect 44886 33170 44938 33182
rect 46118 33178 46170 33190
rect 43878 33114 43930 33126
rect 46118 33114 46170 33126
rect 40014 33058 40066 33070
rect 1344 32954 49616 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 49616 32954
rect 1344 32868 49616 32902
rect 8766 32786 8818 32798
rect 8766 32722 8818 32734
rect 25342 32786 25394 32798
rect 25342 32722 25394 32734
rect 32566 32674 32618 32686
rect 19406 32601 19458 32613
rect 32566 32610 32618 32622
rect 33126 32674 33178 32686
rect 35142 32674 35194 32686
rect 33126 32610 33178 32622
rect 33350 32618 33402 32630
rect 33966 32618 34018 32630
rect 5070 32562 5122 32574
rect 7074 32510 7086 32562
rect 7138 32510 7150 32562
rect 7410 32525 7422 32577
rect 7474 32525 7486 32577
rect 9102 32562 9154 32574
rect 5070 32498 5122 32510
rect 9102 32498 9154 32510
rect 9998 32562 10050 32574
rect 10770 32510 10782 32562
rect 10834 32510 10846 32562
rect 13234 32525 13246 32577
rect 13298 32525 13310 32577
rect 13570 32510 13582 32562
rect 13634 32510 13646 32562
rect 14354 32537 14366 32589
rect 14418 32537 14430 32589
rect 19182 32562 19234 32574
rect 16258 32510 16270 32562
rect 16322 32510 16334 32562
rect 17378 32510 17390 32562
rect 17442 32510 17454 32562
rect 17714 32510 17726 32562
rect 17778 32510 17790 32562
rect 18274 32510 18286 32562
rect 18338 32510 18350 32562
rect 18498 32510 18510 32562
rect 18562 32510 18574 32562
rect 20190 32562 20242 32574
rect 19406 32537 19458 32549
rect 19842 32510 19854 32562
rect 19906 32510 19918 32562
rect 9998 32498 10050 32510
rect 19182 32498 19234 32510
rect 20190 32498 20242 32510
rect 20302 32562 20354 32574
rect 20302 32498 20354 32510
rect 20862 32562 20914 32574
rect 20862 32498 20914 32510
rect 21758 32562 21810 32574
rect 25678 32562 25730 32574
rect 22530 32510 22542 32562
rect 22594 32510 22606 32562
rect 21758 32498 21810 32510
rect 25678 32498 25730 32510
rect 28702 32562 28754 32574
rect 29138 32510 29150 32562
rect 29202 32510 29214 32562
rect 31042 32537 31054 32589
rect 31106 32537 31118 32589
rect 31614 32562 31666 32574
rect 33350 32554 33402 32566
rect 33630 32590 33682 32602
rect 33842 32566 33854 32618
rect 33906 32566 33918 32618
rect 33966 32554 34018 32566
rect 34302 32597 34354 32609
rect 33630 32526 33682 32538
rect 34402 32566 34414 32618
rect 34466 32566 34478 32618
rect 34638 32590 34690 32602
rect 34302 32533 34354 32545
rect 34850 32566 34862 32618
rect 34914 32566 34926 32618
rect 35142 32610 35194 32622
rect 39006 32674 39058 32686
rect 39006 32610 39058 32622
rect 39454 32597 39506 32609
rect 36318 32562 36370 32574
rect 34638 32526 34690 32538
rect 35522 32510 35534 32562
rect 35586 32510 35598 32562
rect 37090 32510 37102 32562
rect 37154 32510 37166 32562
rect 39454 32533 39506 32545
rect 39566 32590 39618 32602
rect 39566 32526 39618 32538
rect 39846 32597 39898 32609
rect 40002 32566 40014 32618
rect 40066 32566 40078 32618
rect 43000 32600 43052 32612
rect 39846 32533 39898 32545
rect 40294 32562 40346 32574
rect 28702 32498 28754 32510
rect 31614 32498 31666 32510
rect 36318 32498 36370 32510
rect 40294 32498 40346 32510
rect 40798 32562 40850 32574
rect 42702 32562 42754 32574
rect 42018 32510 42030 32562
rect 42082 32510 42094 32562
rect 42242 32510 42254 32562
rect 42306 32510 42318 32562
rect 42802 32510 42814 32562
rect 42866 32510 42878 32562
rect 43000 32536 43052 32548
rect 44258 32510 44270 32562
rect 44322 32510 44334 32562
rect 44594 32510 44606 32562
rect 44658 32510 44670 32562
rect 45042 32510 45054 32562
rect 45106 32510 45118 32562
rect 45266 32510 45278 32562
rect 45330 32510 45342 32562
rect 45826 32537 45838 32589
rect 45890 32537 45902 32589
rect 47954 32510 47966 32562
rect 48018 32510 48030 32562
rect 48626 32510 48638 32562
rect 48690 32510 48702 32562
rect 40798 32498 40850 32510
rect 42702 32498 42754 32510
rect 9718 32450 9770 32462
rect 17278 32450 17330 32462
rect 2370 32398 2382 32450
rect 2434 32398 2446 32450
rect 4274 32398 4286 32450
rect 4338 32398 4350 32450
rect 7522 32398 7534 32450
rect 7586 32398 7598 32450
rect 12674 32398 12686 32450
rect 12738 32398 12750 32450
rect 13122 32398 13134 32450
rect 13186 32398 13198 32450
rect 9718 32386 9770 32398
rect 17278 32386 17330 32398
rect 19518 32450 19570 32462
rect 43374 32450 43426 32462
rect 24434 32398 24446 32450
rect 24498 32398 24510 32450
rect 26002 32398 26014 32450
rect 26066 32398 26078 32450
rect 27906 32398 27918 32450
rect 27970 32398 27982 32450
rect 45154 32398 45166 32450
rect 45218 32398 45230 32450
rect 19518 32386 19570 32398
rect 21198 32338 21250 32350
rect 20570 32286 20582 32338
rect 20634 32286 20646 32338
rect 21198 32274 21250 32286
rect 31950 32338 32002 32350
rect 31950 32274 32002 32286
rect 41134 32338 41186 32350
rect 42242 32342 42254 32394
rect 42306 32342 42318 32394
rect 43374 32386 43426 32398
rect 41134 32274 41186 32286
rect 1344 32170 49616 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 49616 32170
rect 1344 32084 49616 32118
rect 11006 32002 11058 32014
rect 4622 31946 4674 31958
rect 11006 31938 11058 31950
rect 22934 32002 22986 32014
rect 38670 32002 38722 32014
rect 22934 31938 22986 31950
rect 36262 31946 36314 31958
rect 3602 31838 3614 31890
rect 3666 31838 3678 31890
rect 4622 31882 4674 31894
rect 21422 31890 21474 31902
rect 26574 31890 26626 31902
rect 48862 32002 48914 32014
rect 38670 31938 38722 31950
rect 45222 31946 45274 31958
rect 8530 31838 8542 31890
rect 8594 31838 8606 31890
rect 9650 31838 9662 31890
rect 9714 31838 9726 31890
rect 16594 31838 16606 31890
rect 16658 31838 16670 31890
rect 20514 31838 20526 31890
rect 20578 31838 20590 31890
rect 24322 31838 24334 31890
rect 24386 31838 24398 31890
rect 27066 31838 27078 31890
rect 27130 31838 27142 31890
rect 27850 31838 27862 31890
rect 27914 31838 27926 31890
rect 29810 31838 29822 31890
rect 29874 31838 29886 31890
rect 31714 31838 31726 31890
rect 31778 31838 31790 31890
rect 32162 31838 32174 31890
rect 32226 31838 32238 31890
rect 33842 31838 33854 31890
rect 33906 31838 33918 31890
rect 36262 31882 36314 31894
rect 48862 31938 48914 31950
rect 40674 31838 40686 31890
rect 40738 31838 40750 31890
rect 42578 31838 42590 31890
rect 42642 31838 42654 31890
rect 45222 31882 45274 31894
rect 21422 31826 21474 31838
rect 26574 31826 26626 31838
rect 5518 31778 5570 31790
rect 3154 31726 3166 31778
rect 3218 31726 3230 31778
rect 3490 31682 3502 31734
rect 3554 31682 3566 31734
rect 4722 31726 4734 31778
rect 4786 31726 4798 31778
rect 4946 31726 4958 31778
rect 5010 31726 5022 31778
rect 5518 31714 5570 31726
rect 5742 31778 5794 31790
rect 5742 31714 5794 31726
rect 9326 31778 9378 31790
rect 12126 31778 12178 31790
rect 9326 31714 9378 31726
rect 9762 31711 9774 31763
rect 9826 31711 9838 31763
rect 10098 31726 10110 31778
rect 10162 31726 10174 31778
rect 11237 31726 11249 31778
rect 11301 31726 11313 31778
rect 12126 31714 12178 31726
rect 12798 31778 12850 31790
rect 12798 31714 12850 31726
rect 13022 31778 13074 31790
rect 17838 31778 17890 31790
rect 22094 31778 22146 31790
rect 25958 31778 26010 31790
rect 13346 31726 13358 31778
rect 13410 31726 13422 31778
rect 14254 31750 14306 31762
rect 13022 31714 13074 31726
rect 13918 31722 13970 31734
rect 6638 31666 6690 31678
rect 14018 31670 14030 31722
rect 14082 31670 14094 31722
rect 14254 31686 14306 31698
rect 14478 31750 14530 31762
rect 17602 31698 17614 31750
rect 17666 31698 17678 31750
rect 18610 31726 18622 31778
rect 18674 31726 18686 31778
rect 21970 31726 21982 31778
rect 22034 31726 22046 31778
rect 22642 31726 22654 31778
rect 22706 31726 22718 31778
rect 23214 31750 23266 31762
rect 17838 31714 17890 31726
rect 14478 31686 14530 31698
rect 6010 31614 6022 31666
rect 6074 31614 6086 31666
rect 12506 31614 12518 31666
rect 12570 31614 12582 31666
rect 13918 31658 13970 31670
rect 14758 31666 14810 31678
rect 21802 31670 21814 31722
rect 21866 31670 21878 31722
rect 22094 31714 22146 31726
rect 23214 31686 23266 31698
rect 23438 31750 23490 31762
rect 23438 31686 23490 31698
rect 23662 31750 23714 31762
rect 23662 31686 23714 31698
rect 23774 31743 23826 31755
rect 23774 31679 23826 31691
rect 24434 31682 24446 31734
rect 24498 31682 24510 31734
rect 24770 31726 24782 31778
rect 24834 31726 24846 31778
rect 25118 31743 25170 31755
rect 25118 31679 25170 31691
rect 25286 31743 25338 31755
rect 25286 31679 25338 31691
rect 25454 31750 25506 31762
rect 25454 31686 25506 31698
rect 25678 31750 25730 31762
rect 25958 31714 26010 31726
rect 26238 31778 26290 31790
rect 26238 31714 26290 31726
rect 27358 31778 27410 31790
rect 27358 31714 27410 31726
rect 27582 31778 27634 31790
rect 27582 31714 27634 31726
rect 28142 31778 28194 31790
rect 28142 31714 28194 31726
rect 28366 31778 28418 31790
rect 28366 31714 28418 31726
rect 29038 31778 29090 31790
rect 33070 31778 33122 31790
rect 39902 31778 39954 31790
rect 29038 31714 29090 31726
rect 25678 31686 25730 31698
rect 32274 31682 32286 31734
rect 32338 31682 32350 31734
rect 32610 31726 32622 31778
rect 32674 31726 32686 31778
rect 36082 31726 36094 31778
rect 36146 31726 36158 31778
rect 33070 31714 33122 31726
rect 37314 31698 37326 31750
rect 37378 31698 37390 31750
rect 39902 31714 39954 31726
rect 42926 31778 42978 31790
rect 42926 31714 42978 31726
rect 44158 31778 44210 31790
rect 48526 31778 48578 31790
rect 45378 31726 45390 31778
rect 45442 31726 45454 31778
rect 47730 31726 47742 31778
rect 47794 31726 47806 31778
rect 44158 31714 44210 31726
rect 48526 31714 48578 31726
rect 49198 31778 49250 31790
rect 49198 31714 49250 31726
rect 35758 31666 35810 31678
rect 6638 31602 6690 31614
rect 14758 31602 14810 31614
rect 22486 31610 22538 31622
rect 10614 31554 10666 31566
rect 10614 31490 10666 31502
rect 13526 31554 13578 31566
rect 35758 31602 35810 31614
rect 45838 31666 45890 31678
rect 45838 31602 45890 31614
rect 22486 31546 22538 31558
rect 43262 31554 43314 31566
rect 13526 31490 13578 31502
rect 43262 31490 43314 31502
rect 43822 31554 43874 31566
rect 43822 31490 43874 31502
rect 1344 31386 49616 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 49616 31386
rect 1344 31300 49616 31334
rect 10390 31218 10442 31230
rect 10390 31154 10442 31166
rect 11902 31218 11954 31230
rect 11902 31154 11954 31166
rect 16606 31218 16658 31230
rect 30382 31218 30434 31230
rect 16606 31154 16658 31166
rect 19126 31162 19178 31174
rect 5686 31106 5738 31118
rect 5686 31042 5738 31054
rect 7310 31106 7362 31118
rect 7310 31042 7362 31054
rect 12518 31106 12570 31118
rect 30382 31154 30434 31166
rect 40294 31218 40346 31230
rect 40294 31154 40346 31166
rect 46174 31218 46226 31230
rect 46174 31154 46226 31166
rect 46790 31218 46842 31230
rect 46790 31154 46842 31166
rect 47910 31218 47962 31230
rect 47910 31154 47962 31166
rect 48974 31218 49026 31230
rect 48974 31154 49026 31166
rect 19126 31098 19178 31110
rect 31558 31106 31610 31118
rect 12518 31042 12570 31054
rect 12742 31050 12794 31062
rect 20302 31050 20354 31062
rect 26126 31050 26178 31062
rect 28634 31054 28646 31106
rect 28698 31054 28710 31106
rect 34470 31106 34522 31118
rect 1598 30994 1650 31006
rect 1598 30930 1650 30942
rect 4958 30994 5010 31006
rect 5406 30994 5458 31006
rect 4958 30930 5010 30942
rect 5126 30938 5178 30950
rect 5282 30942 5294 30994
rect 5346 30942 5358 30994
rect 5406 30930 5458 30942
rect 6190 30994 6242 31006
rect 11006 30994 11058 31006
rect 7054 30942 7066 30994
rect 7118 30942 7130 30994
rect 6190 30930 6242 30942
rect 11006 30930 11058 30942
rect 12238 30994 12290 31006
rect 12742 30986 12794 30998
rect 13022 31022 13074 31034
rect 13022 30958 13074 30970
rect 13246 31022 13298 31034
rect 13246 30958 13298 30970
rect 13358 31029 13410 31041
rect 15586 30998 15598 31050
rect 15650 30998 15662 31050
rect 15810 30998 15822 31050
rect 15874 30998 15886 31050
rect 16034 30998 16046 31050
rect 16098 30998 16110 31050
rect 16158 31029 16210 31041
rect 13358 30965 13410 30977
rect 13682 30942 13694 30994
rect 13746 30942 13758 30994
rect 14018 30942 14030 30994
rect 14082 30942 14094 30994
rect 14578 30942 14590 30994
rect 14642 30942 14654 30994
rect 14802 30942 14814 30994
rect 14866 30942 14878 30994
rect 16158 30965 16210 30977
rect 16942 30994 16994 31006
rect 12238 30930 12290 30942
rect 16942 30930 16994 30942
rect 17390 30994 17442 31006
rect 18254 30998 18266 31050
rect 18318 30998 18330 31050
rect 19406 30994 19458 31006
rect 18946 30942 18958 30994
rect 19010 30942 19022 30994
rect 17390 30930 17442 30942
rect 19406 30930 19458 30942
rect 19630 30994 19682 31006
rect 20402 30998 20414 31050
rect 20466 30998 20478 31050
rect 20638 31022 20690 31034
rect 20302 30986 20354 30998
rect 20850 30998 20862 31050
rect 20914 30998 20926 31050
rect 22284 31031 22336 31043
rect 20638 30958 20690 30970
rect 21142 30994 21194 31006
rect 19630 30930 19682 30942
rect 25510 31029 25562 31041
rect 22542 30994 22594 31006
rect 22284 30967 22336 30979
rect 22418 30942 22430 30994
rect 22482 30942 22494 30994
rect 21142 30930 21194 30942
rect 22542 30930 22594 30942
rect 22766 30994 22818 31006
rect 22766 30930 22818 30942
rect 22990 30994 23042 31006
rect 22990 30930 23042 30942
rect 24110 30994 24162 31006
rect 24110 30930 24162 30942
rect 24222 30994 24274 31006
rect 24222 30930 24274 30942
rect 24558 30994 24610 31006
rect 25510 30965 25562 30977
rect 25790 31022 25842 31034
rect 25790 30958 25842 30970
rect 25958 31029 26010 31041
rect 31558 31042 31610 31054
rect 32398 31050 32450 31062
rect 26126 30986 26178 30998
rect 26798 30994 26850 31006
rect 25958 30965 26010 30977
rect 24558 30930 24610 30942
rect 26798 30930 26850 30942
rect 28926 30994 28978 31006
rect 28926 30930 28978 30942
rect 29038 30994 29090 31006
rect 29038 30930 29090 30942
rect 30718 30994 30770 31006
rect 30718 30930 30770 30942
rect 31110 30994 31162 31006
rect 31826 30998 31838 31050
rect 31890 30998 31902 31050
rect 32050 30998 32062 31050
rect 32114 30998 32126 31050
rect 32286 31022 32338 31034
rect 32398 30986 32450 30998
rect 33630 31050 33682 31062
rect 34022 31050 34074 31062
rect 33630 30986 33682 30998
rect 33742 31022 33794 31034
rect 32286 30958 32338 30970
rect 34178 30998 34190 31050
rect 34242 30998 34254 31050
rect 34470 31042 34522 31054
rect 38446 31106 38498 31118
rect 39734 31106 39786 31118
rect 38446 31042 38498 31054
rect 38819 31050 38871 31062
rect 34022 30986 34074 30998
rect 34974 30994 35026 31006
rect 33742 30958 33794 30970
rect 31110 30930 31162 30942
rect 34974 30930 35026 30942
rect 35198 30994 35250 31006
rect 35198 30930 35250 30942
rect 35758 30994 35810 31006
rect 36530 30942 36542 30994
rect 36594 30942 36606 30994
rect 38819 30986 38871 30998
rect 39006 31022 39058 31034
rect 39006 30958 39058 30970
rect 39230 31022 39282 31034
rect 39442 30998 39454 31050
rect 39506 30998 39518 31050
rect 39734 31042 39786 31054
rect 42254 31106 42306 31118
rect 42254 31042 42306 31054
rect 40910 31029 40962 31041
rect 39230 30958 39282 30970
rect 40450 30942 40462 30994
rect 40514 30942 40526 30994
rect 40910 30965 40962 30977
rect 41022 31022 41074 31034
rect 41022 30958 41074 30970
rect 41246 31022 41298 31034
rect 41246 30958 41298 30970
rect 41496 30958 41508 31010
rect 41560 30958 41572 31010
rect 42590 30994 42642 31006
rect 35758 30930 35810 30942
rect 42590 30930 42642 30942
rect 42814 30994 42866 31006
rect 45838 30994 45890 31006
rect 48638 30994 48690 31006
rect 43586 30942 43598 30994
rect 43650 30942 43662 30994
rect 47170 30942 47182 30994
rect 47234 30942 47246 30994
rect 47394 30942 47406 30994
rect 47458 30942 47470 30994
rect 47730 30942 47742 30994
rect 47794 30942 47806 30994
rect 42814 30930 42866 30942
rect 45838 30930 45890 30942
rect 48638 30930 48690 30942
rect 2370 30830 2382 30882
rect 2434 30830 2446 30882
rect 4274 30830 4286 30882
rect 4338 30830 4350 30882
rect 5126 30874 5178 30886
rect 15038 30882 15090 30894
rect 15038 30818 15090 30830
rect 26630 30882 26682 30894
rect 26630 30818 26682 30830
rect 27750 30882 27802 30894
rect 27750 30818 27802 30830
rect 33238 30882 33290 30894
rect 45490 30830 45502 30882
rect 45554 30830 45566 30882
rect 33238 30818 33290 30830
rect 47518 30826 47570 30838
rect 11342 30770 11394 30782
rect 11342 30706 11394 30718
rect 15318 30770 15370 30782
rect 15318 30706 15370 30718
rect 18510 30770 18562 30782
rect 21870 30770 21922 30782
rect 23774 30770 23826 30782
rect 19898 30718 19910 30770
rect 19962 30718 19974 30770
rect 23258 30718 23270 30770
rect 23322 30718 23334 30770
rect 18510 30706 18562 30718
rect 21870 30706 21922 30718
rect 23774 30706 23826 30718
rect 25286 30770 25338 30782
rect 25286 30706 25338 30718
rect 27134 30770 27186 30782
rect 41750 30770 41802 30782
rect 35466 30718 35478 30770
rect 35530 30718 35542 30770
rect 47518 30762 47570 30774
rect 27134 30706 27186 30718
rect 41750 30706 41802 30718
rect 1344 30602 49616 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 49616 30602
rect 1344 30516 49616 30550
rect 2494 30434 2546 30446
rect 2494 30370 2546 30382
rect 12406 30434 12458 30446
rect 22150 30434 22202 30446
rect 32734 30434 32786 30446
rect 12406 30370 12458 30382
rect 20302 30378 20354 30390
rect 16382 30322 16434 30334
rect 32106 30382 32118 30434
rect 32170 30382 32182 30434
rect 22150 30370 22202 30382
rect 32734 30370 32786 30382
rect 44102 30434 44154 30446
rect 44102 30370 44154 30382
rect 45670 30434 45722 30446
rect 45670 30370 45722 30382
rect 4946 30270 4958 30322
rect 5010 30270 5022 30322
rect 18162 30270 18174 30322
rect 18226 30270 18238 30322
rect 20302 30314 20354 30326
rect 38166 30322 38218 30334
rect 27906 30270 27918 30322
rect 27970 30270 27982 30322
rect 41906 30270 41918 30322
rect 41970 30270 41982 30322
rect 16382 30258 16434 30270
rect 38166 30258 38218 30270
rect 2830 30210 2882 30222
rect 2830 30146 2882 30158
rect 4062 30210 4114 30222
rect 4062 30146 4114 30158
rect 4398 30210 4450 30222
rect 6302 30210 6354 30222
rect 7534 30210 7586 30222
rect 5058 30158 5070 30210
rect 5122 30158 5134 30210
rect 5618 30158 5630 30210
rect 5682 30158 5694 30210
rect 6850 30158 6862 30210
rect 6914 30158 6926 30210
rect 4398 30146 4450 30158
rect 4722 30102 4734 30154
rect 4786 30102 4798 30154
rect 5898 30102 5910 30154
rect 5962 30102 5974 30154
rect 6302 30146 6354 30158
rect 7186 30114 7198 30166
rect 7250 30114 7262 30166
rect 7534 30146 7586 30158
rect 8318 30210 8370 30222
rect 11006 30210 11058 30222
rect 9090 30158 9102 30210
rect 9154 30158 9166 30210
rect 8318 30146 8370 30158
rect 11006 30146 11058 30158
rect 11454 30210 11506 30222
rect 11454 30146 11506 30158
rect 11678 30210 11730 30222
rect 15710 30210 15762 30222
rect 15988 30210 16040 30222
rect 17614 30210 17666 30222
rect 18846 30210 18898 30222
rect 12226 30158 12238 30210
rect 12290 30158 12302 30210
rect 13906 30158 13918 30210
rect 13970 30158 13982 30210
rect 14758 30175 14810 30187
rect 11678 30146 11730 30158
rect 14758 30111 14810 30123
rect 15038 30182 15090 30194
rect 15374 30154 15426 30166
rect 15038 30118 15090 30130
rect 14534 30098 14586 30110
rect 15250 30102 15262 30154
rect 15314 30102 15326 30154
rect 15810 30158 15822 30210
rect 15874 30158 15886 30210
rect 16930 30158 16942 30210
rect 16994 30158 17006 30210
rect 15710 30146 15762 30158
rect 15988 30146 16040 30158
rect 17266 30131 17278 30183
rect 17330 30131 17342 30183
rect 17614 30146 17666 30158
rect 18274 30114 18286 30166
rect 18338 30114 18350 30166
rect 18610 30158 18622 30210
rect 18674 30158 18686 30210
rect 18846 30146 18898 30158
rect 19070 30210 19122 30222
rect 19910 30210 19962 30222
rect 22766 30210 22818 30222
rect 26014 30210 26066 30222
rect 19338 30158 19350 30210
rect 19402 30158 19414 30210
rect 20402 30158 20414 30210
rect 20466 30158 20478 30210
rect 20738 30158 20750 30210
rect 20802 30158 20814 30210
rect 21422 30182 21474 30194
rect 19070 30146 19122 30158
rect 19910 30146 19962 30158
rect 21310 30154 21362 30166
rect 11946 30046 11958 30098
rect 12010 30046 12022 30098
rect 14086 30042 14138 30054
rect 5730 29990 5742 30042
rect 5794 29990 5806 30042
rect 7074 29990 7086 30042
rect 7138 29990 7150 30042
rect 7870 29986 7922 29998
rect 15374 30090 15426 30102
rect 21422 30118 21474 30130
rect 21702 30175 21754 30187
rect 21702 30111 21754 30123
rect 21926 30175 21978 30187
rect 23538 30158 23550 30210
rect 23602 30158 23614 30210
rect 22766 30146 22818 30158
rect 26014 30146 26066 30158
rect 28702 30210 28754 30222
rect 28702 30146 28754 30158
rect 31726 30210 31778 30222
rect 31726 30146 31778 30158
rect 31838 30210 31890 30222
rect 31838 30146 31890 30158
rect 32398 30210 32450 30222
rect 32398 30146 32450 30158
rect 33070 30210 33122 30222
rect 33070 30146 33122 30158
rect 33294 30210 33346 30222
rect 34638 30210 34690 30222
rect 35870 30210 35922 30222
rect 33562 30158 33574 30210
rect 33626 30158 33638 30210
rect 33954 30158 33966 30210
rect 34018 30158 34030 30210
rect 35186 30158 35198 30210
rect 35250 30158 35262 30210
rect 38670 30210 38722 30222
rect 33294 30146 33346 30158
rect 21926 30111 21978 30123
rect 21310 30090 21362 30102
rect 25454 30098 25506 30110
rect 34290 30102 34302 30154
rect 34354 30102 34366 30154
rect 34638 30146 34690 30158
rect 35522 30102 35534 30154
rect 35586 30102 35598 30154
rect 35870 30146 35922 30158
rect 37326 30175 37378 30187
rect 37326 30111 37378 30123
rect 37438 30182 37490 30194
rect 37886 30182 37938 30194
rect 37438 30118 37490 30130
rect 37650 30102 37662 30154
rect 37714 30102 37726 30154
rect 38670 30146 38722 30158
rect 39006 30210 39058 30222
rect 39006 30146 39058 30158
rect 39230 30210 39282 30222
rect 42254 30210 42306 30222
rect 40002 30158 40014 30210
rect 40066 30158 40078 30210
rect 46398 30210 46450 30222
rect 43598 30182 43650 30194
rect 39230 30146 39282 30158
rect 42254 30146 42306 30158
rect 43262 30154 43314 30166
rect 37886 30118 37938 30130
rect 43362 30102 43374 30154
rect 43426 30102 43438 30154
rect 43598 30118 43650 30130
rect 43822 30182 43874 30194
rect 45166 30182 45218 30194
rect 43822 30118 43874 30130
rect 44830 30154 44882 30166
rect 44930 30102 44942 30154
rect 44994 30102 45006 30154
rect 45166 30118 45218 30130
rect 45390 30182 45442 30194
rect 47170 30158 47182 30210
rect 47234 30158 47246 30210
rect 46398 30146 46450 30158
rect 45390 30118 45442 30130
rect 14534 30034 14586 30046
rect 43262 30090 43314 30102
rect 44830 30090 44882 30102
rect 49086 30098 49138 30110
rect 17714 29990 17726 30042
rect 17778 29990 17790 30042
rect 25454 30034 25506 30046
rect 34178 29990 34190 30042
rect 34242 29990 34254 30042
rect 35298 29990 35310 30042
rect 35362 29990 35374 30042
rect 49086 30034 49138 30046
rect 14086 29978 14138 29990
rect 42590 29986 42642 29998
rect 7870 29922 7922 29934
rect 42590 29922 42642 29934
rect 46230 29986 46282 29998
rect 46230 29922 46282 29934
rect 1344 29818 49616 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 49616 29818
rect 1344 29732 49616 29766
rect 9046 29650 9098 29662
rect 9046 29586 9098 29598
rect 14982 29650 15034 29662
rect 4622 29538 4674 29550
rect 4622 29474 4674 29486
rect 10446 29538 10498 29550
rect 12674 29542 12686 29594
rect 12738 29542 12750 29594
rect 14982 29586 15034 29598
rect 15654 29650 15706 29662
rect 15654 29586 15706 29598
rect 24446 29650 24498 29662
rect 22530 29542 22542 29594
rect 22594 29542 22606 29594
rect 24446 29586 24498 29598
rect 33574 29650 33626 29662
rect 33574 29586 33626 29598
rect 35366 29650 35418 29662
rect 10446 29474 10498 29486
rect 24054 29538 24106 29550
rect 26966 29538 27018 29550
rect 34066 29542 34078 29594
rect 34130 29542 34142 29594
rect 35366 29586 35418 29598
rect 40126 29650 40178 29662
rect 40126 29586 40178 29598
rect 47014 29650 47066 29662
rect 47014 29586 47066 29598
rect 1934 29426 1986 29438
rect 5282 29374 5294 29426
rect 5346 29374 5358 29426
rect 7522 29401 7534 29453
rect 7586 29401 7598 29453
rect 8194 29389 8206 29441
rect 8258 29389 8270 29441
rect 8530 29374 8542 29426
rect 8594 29374 8606 29426
rect 9650 29418 9662 29470
rect 9714 29418 9726 29470
rect 10677 29430 10689 29482
rect 10741 29430 10753 29482
rect 12350 29465 12402 29477
rect 11566 29426 11618 29438
rect 9986 29374 9998 29426
rect 10050 29374 10062 29426
rect 1934 29362 1986 29374
rect 11566 29362 11618 29374
rect 12126 29426 12178 29438
rect 17278 29426 17330 29438
rect 12350 29401 12402 29413
rect 12786 29374 12798 29426
rect 12850 29374 12862 29426
rect 15138 29374 15150 29426
rect 15202 29374 15214 29426
rect 15754 29374 15766 29426
rect 15818 29374 15830 29426
rect 15922 29374 15934 29426
rect 15986 29374 15998 29426
rect 12126 29362 12178 29374
rect 17278 29362 17330 29374
rect 19966 29426 20018 29438
rect 21074 29418 21086 29470
rect 21138 29418 21150 29470
rect 22206 29465 22258 29477
rect 24054 29474 24106 29486
rect 26126 29482 26178 29494
rect 46454 29538 46506 29550
rect 47842 29542 47854 29594
rect 47906 29542 47918 29594
rect 21982 29426 22034 29438
rect 21298 29374 21310 29426
rect 21362 29374 21374 29426
rect 22878 29426 22930 29438
rect 22206 29401 22258 29413
rect 22642 29374 22654 29426
rect 22706 29374 22718 29426
rect 19966 29362 20018 29374
rect 21982 29362 22034 29374
rect 22878 29362 22930 29374
rect 23102 29426 23154 29438
rect 23102 29362 23154 29374
rect 24782 29426 24834 29438
rect 24782 29362 24834 29374
rect 25342 29426 25394 29438
rect 26126 29418 26178 29430
rect 26238 29454 26290 29466
rect 26450 29430 26462 29482
rect 26514 29430 26526 29482
rect 26674 29430 26686 29482
rect 26738 29430 26750 29482
rect 26966 29474 27018 29486
rect 44382 29482 44434 29494
rect 44998 29482 45050 29494
rect 27806 29426 27858 29438
rect 26238 29390 26290 29402
rect 27514 29374 27526 29426
rect 27578 29374 27590 29426
rect 25342 29362 25394 29374
rect 27806 29362 27858 29374
rect 28030 29426 28082 29438
rect 28030 29362 28082 29374
rect 28142 29426 28194 29438
rect 28142 29362 28194 29374
rect 31278 29426 31330 29438
rect 31278 29362 31330 29374
rect 31390 29426 31442 29438
rect 33394 29374 33406 29426
rect 33458 29374 33470 29426
rect 33954 29374 33966 29426
rect 34018 29374 34030 29426
rect 34290 29401 34302 29453
rect 34354 29401 34366 29453
rect 34638 29426 34690 29438
rect 35970 29401 35982 29453
rect 36034 29401 36046 29453
rect 40462 29426 40514 29438
rect 38546 29374 38558 29426
rect 38610 29374 38622 29426
rect 38770 29374 38782 29426
rect 38834 29374 38846 29426
rect 39442 29374 39454 29426
rect 39506 29374 39518 29426
rect 31390 29362 31442 29374
rect 34638 29362 34690 29374
rect 40462 29362 40514 29374
rect 41078 29426 41130 29438
rect 41458 29401 41470 29453
rect 41522 29401 41534 29453
rect 44482 29430 44494 29482
rect 44546 29430 44558 29482
rect 44706 29430 44718 29482
rect 44770 29430 44782 29482
rect 46454 29474 46506 29486
rect 44382 29418 44434 29430
rect 44998 29418 45050 29430
rect 45222 29426 45274 29438
rect 41078 29362 41130 29374
rect 45222 29362 45274 29374
rect 45502 29426 45554 29438
rect 47406 29426 47458 29438
rect 47170 29374 47182 29426
rect 47234 29374 47246 29426
rect 48066 29374 48078 29426
rect 48130 29374 48142 29426
rect 45502 29362 45554 29374
rect 47406 29362 47458 29374
rect 2706 29262 2718 29314
rect 2770 29262 2782 29314
rect 8082 29262 8094 29314
rect 8146 29262 8158 29314
rect 9538 29262 9550 29314
rect 9602 29262 9614 29314
rect 18050 29262 18062 29314
rect 18114 29262 18126 29314
rect 20962 29262 20974 29314
rect 21026 29262 21038 29314
rect 28914 29262 28926 29314
rect 28978 29262 28990 29314
rect 30818 29262 30830 29314
rect 30882 29262 30894 29314
rect 38446 29258 38498 29270
rect 25678 29202 25730 29214
rect 23370 29150 23382 29202
rect 23434 29150 23446 29202
rect 31658 29150 31670 29202
rect 31722 29150 31734 29202
rect 38446 29194 38498 29206
rect 39286 29202 39338 29214
rect 25678 29138 25730 29150
rect 39286 29138 39338 29150
rect 42814 29202 42866 29214
rect 42814 29138 42866 29150
rect 45838 29202 45890 29214
rect 45838 29138 45890 29150
rect 1344 29034 49616 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 49616 29034
rect 1344 28948 49616 28982
rect 16942 28866 16994 28878
rect 11386 28814 11398 28866
rect 11450 28814 11462 28866
rect 16942 28802 16994 28814
rect 18398 28866 18450 28878
rect 18398 28802 18450 28814
rect 19294 28866 19346 28878
rect 19294 28802 19346 28814
rect 22598 28866 22650 28878
rect 22598 28802 22650 28814
rect 24950 28866 25002 28878
rect 35366 28866 35418 28878
rect 30314 28814 30326 28866
rect 30378 28814 30390 28866
rect 33338 28814 33350 28866
rect 33402 28814 33414 28866
rect 24950 28802 25002 28814
rect 5742 28754 5794 28766
rect 25734 28754 25786 28766
rect 3602 28702 3614 28754
rect 3666 28702 3678 28754
rect 7746 28702 7758 28754
rect 7810 28702 7822 28754
rect 12114 28702 12126 28754
rect 12178 28702 12190 28754
rect 5742 28690 5794 28702
rect 25734 28690 25786 28702
rect 28534 28754 28586 28766
rect 31826 28758 31838 28810
rect 31890 28758 31902 28810
rect 35366 28802 35418 28814
rect 43934 28866 43986 28878
rect 43934 28802 43986 28814
rect 36038 28754 36090 28766
rect 32610 28702 32622 28754
rect 32674 28702 32686 28754
rect 28534 28690 28586 28702
rect 36038 28690 36090 28702
rect 37886 28754 37938 28766
rect 42242 28702 42254 28754
rect 42306 28702 42318 28754
rect 44930 28702 44942 28754
rect 44994 28702 45006 28754
rect 46834 28702 46846 28754
rect 46898 28702 46910 28754
rect 37886 28690 37938 28702
rect 4286 28642 4338 28654
rect 6974 28642 7026 28654
rect 2930 28590 2942 28642
rect 2994 28590 3006 28642
rect 3110 28612 3162 28624
rect 3714 28575 3726 28627
rect 3778 28575 3790 28627
rect 3938 28590 3950 28642
rect 4002 28590 4014 28642
rect 4286 28578 4338 28590
rect 5574 28586 5626 28598
rect 5954 28590 5966 28642
rect 6018 28590 6030 28642
rect 3110 28548 3162 28560
rect 5574 28522 5626 28534
rect 6302 28586 6354 28598
rect 6974 28578 7026 28590
rect 11678 28642 11730 28654
rect 11678 28578 11730 28590
rect 11902 28642 11954 28654
rect 13358 28642 13410 28654
rect 11902 28578 11954 28590
rect 12226 28575 12238 28627
rect 12290 28575 12302 28627
rect 12450 28590 12462 28642
rect 12514 28590 12526 28642
rect 13358 28578 13410 28590
rect 13694 28642 13746 28654
rect 13694 28578 13746 28590
rect 14814 28642 14866 28654
rect 14814 28578 14866 28590
rect 15262 28642 15314 28654
rect 17278 28642 17330 28654
rect 15922 28590 15934 28642
rect 15986 28590 15998 28642
rect 6302 28522 6354 28534
rect 9662 28530 9714 28542
rect 14970 28534 14982 28586
rect 15034 28534 15046 28586
rect 15262 28578 15314 28590
rect 16258 28575 16270 28627
rect 16322 28575 16334 28627
rect 17278 28578 17330 28590
rect 17390 28642 17442 28654
rect 17390 28578 17442 28590
rect 18062 28642 18114 28654
rect 18062 28578 18114 28590
rect 19630 28642 19682 28654
rect 26798 28642 26850 28654
rect 19630 28578 19682 28590
rect 21646 28614 21698 28626
rect 2930 28422 2942 28474
rect 2994 28422 3006 28474
rect 9662 28466 9714 28478
rect 15150 28530 15202 28542
rect 15150 28466 15202 28478
rect 15542 28530 15594 28542
rect 21242 28534 21254 28586
rect 21306 28534 21318 28586
rect 21410 28534 21422 28586
rect 21474 28534 21486 28586
rect 21646 28550 21698 28562
rect 21870 28614 21922 28626
rect 22418 28590 22430 28642
rect 22482 28590 22494 28642
rect 25106 28590 25118 28642
rect 25170 28590 25182 28642
rect 26462 28614 26514 28626
rect 21870 28550 21922 28562
rect 15542 28466 15594 28478
rect 22150 28530 22202 28542
rect 26002 28534 26014 28586
rect 26066 28534 26078 28586
rect 26226 28534 26238 28586
rect 26290 28534 26302 28586
rect 26462 28550 26514 28562
rect 26574 28607 26626 28619
rect 26798 28578 26850 28590
rect 27134 28642 27186 28654
rect 27918 28642 27970 28654
rect 27626 28590 27638 28642
rect 27690 28590 27702 28642
rect 27134 28578 27186 28590
rect 27918 28578 27970 28590
rect 28142 28642 28194 28654
rect 28142 28578 28194 28590
rect 29486 28642 29538 28654
rect 29486 28578 29538 28590
rect 29710 28642 29762 28654
rect 29710 28578 29762 28590
rect 30606 28642 30658 28654
rect 30606 28578 30658 28590
rect 30830 28642 30882 28654
rect 30830 28578 30882 28590
rect 31054 28642 31106 28654
rect 32846 28642 32898 28654
rect 31714 28590 31726 28642
rect 31778 28590 31790 28642
rect 32162 28590 32174 28642
rect 32226 28590 32238 28642
rect 31054 28578 31106 28590
rect 26574 28543 26626 28555
rect 32498 28546 32510 28598
rect 32562 28546 32574 28598
rect 32846 28578 32898 28590
rect 33070 28642 33122 28654
rect 33070 28578 33122 28590
rect 34302 28642 34354 28654
rect 36486 28642 36538 28654
rect 34302 28578 34354 28590
rect 34526 28603 34578 28615
rect 34962 28590 34974 28642
rect 35026 28590 35038 28642
rect 35186 28590 35198 28642
rect 35250 28590 35262 28642
rect 36486 28578 36538 28590
rect 37214 28642 37266 28654
rect 37214 28578 37266 28590
rect 37550 28642 37602 28654
rect 38894 28642 38946 28654
rect 41582 28642 41634 28654
rect 44270 28642 44322 28654
rect 37550 28578 37602 28590
rect 37774 28603 37826 28615
rect 34526 28539 34578 28551
rect 38210 28590 38222 28642
rect 38274 28590 38286 28642
rect 40786 28590 40798 28642
rect 40850 28590 40862 28642
rect 41906 28590 41918 28642
rect 41970 28590 41982 28642
rect 38894 28578 38946 28590
rect 41582 28578 41634 28590
rect 42130 28575 42142 28627
rect 42194 28575 42206 28627
rect 42522 28574 42534 28626
rect 42586 28574 42598 28626
rect 42702 28614 42754 28626
rect 37774 28539 37826 28551
rect 42702 28550 42754 28562
rect 42926 28614 42978 28626
rect 42926 28550 42978 28562
rect 43150 28614 43202 28626
rect 44270 28578 44322 28590
rect 47630 28642 47682 28654
rect 47630 28578 47682 28590
rect 43150 28550 43202 28562
rect 43430 28530 43482 28542
rect 29194 28478 29206 28530
rect 29258 28478 29270 28530
rect 16146 28422 16158 28474
rect 16210 28422 16222 28474
rect 22150 28466 22202 28478
rect 17726 28418 17778 28430
rect 34178 28422 34190 28474
rect 34242 28422 34254 28474
rect 43430 28466 43482 28478
rect 17726 28354 17778 28366
rect 49254 28418 49306 28430
rect 49254 28354 49306 28366
rect 1344 28250 49616 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 49616 28250
rect 1344 28164 49616 28198
rect 7254 28082 7306 28094
rect 7254 28018 7306 28030
rect 16886 28082 16938 28094
rect 16886 28018 16938 28030
rect 29374 28082 29426 28094
rect 7870 27970 7922 27982
rect 17602 27974 17614 28026
rect 17666 27974 17678 28026
rect 20402 27974 20414 28026
rect 20466 27974 20478 28026
rect 29374 28018 29426 28030
rect 30046 28082 30098 28094
rect 30046 28018 30098 28030
rect 32398 28082 32450 28094
rect 22766 27970 22818 27982
rect 31042 27974 31054 28026
rect 31106 27974 31118 28026
rect 32398 28018 32450 28030
rect 36150 28082 36202 28094
rect 36150 28018 36202 28030
rect 36598 28082 36650 28094
rect 36598 28018 36650 28030
rect 40238 28082 40290 28094
rect 37762 27974 37774 28026
rect 37826 27974 37838 28026
rect 40238 28018 40290 28030
rect 41078 28082 41130 28094
rect 41078 28018 41130 28030
rect 42646 28082 42698 28094
rect 42646 28018 42698 28030
rect 48974 28082 49026 28094
rect 48974 28018 49026 28030
rect 45502 27970 45554 27982
rect 7870 27906 7922 27918
rect 9494 27914 9546 27926
rect 1922 27806 1934 27858
rect 1986 27806 1998 27858
rect 2146 27850 2158 27902
rect 2210 27850 2222 27902
rect 2718 27858 2770 27870
rect 3838 27858 3890 27870
rect 2949 27806 2961 27858
rect 3013 27806 3025 27858
rect 2718 27794 2770 27806
rect 3838 27794 3890 27806
rect 4062 27858 4114 27870
rect 6750 27858 6802 27870
rect 8101 27862 8113 27914
rect 8165 27862 8177 27914
rect 8990 27858 9042 27870
rect 4834 27806 4846 27858
rect 4898 27806 4910 27858
rect 7074 27806 7086 27858
rect 7138 27806 7150 27858
rect 9494 27850 9546 27862
rect 10222 27914 10274 27926
rect 34234 27918 34246 27970
rect 34298 27918 34310 27970
rect 15072 27896 15124 27908
rect 9874 27806 9886 27858
rect 9938 27806 9950 27858
rect 10222 27850 10274 27862
rect 14030 27858 14082 27870
rect 13234 27806 13246 27858
rect 13298 27806 13310 27858
rect 4062 27794 4114 27806
rect 6750 27794 6802 27806
rect 8990 27794 9042 27806
rect 14030 27794 14082 27806
rect 14814 27858 14866 27870
rect 14914 27806 14926 27858
rect 14978 27806 14990 27858
rect 15072 27832 15124 27844
rect 15822 27858 15874 27870
rect 14814 27794 14866 27806
rect 15822 27794 15874 27806
rect 16046 27858 16098 27870
rect 17826 27862 17838 27914
rect 17890 27862 17902 27914
rect 22766 27906 22818 27918
rect 18902 27887 18954 27899
rect 18062 27858 18114 27870
rect 17490 27806 17502 27858
rect 17554 27806 17566 27858
rect 18902 27823 18954 27835
rect 19170 27806 19182 27858
rect 19234 27806 19246 27858
rect 19618 27850 19630 27902
rect 19682 27850 19694 27902
rect 20526 27858 20578 27870
rect 19954 27806 19966 27858
rect 20018 27806 20030 27858
rect 20850 27833 20862 27885
rect 20914 27833 20926 27885
rect 21186 27806 21198 27858
rect 21250 27806 21262 27858
rect 21634 27839 21646 27891
rect 21698 27839 21710 27891
rect 21970 27842 21982 27894
rect 22034 27842 22046 27894
rect 22418 27842 22430 27894
rect 22482 27842 22494 27894
rect 22574 27846 22586 27898
rect 22638 27846 22650 27898
rect 38110 27897 38162 27909
rect 23202 27806 23214 27858
rect 23266 27806 23278 27858
rect 23426 27806 23438 27858
rect 23490 27806 23502 27858
rect 25666 27833 25678 27885
rect 25730 27833 25742 27885
rect 28814 27858 28866 27870
rect 27906 27806 27918 27858
rect 27970 27806 27982 27858
rect 16046 27794 16098 27806
rect 18062 27794 18114 27806
rect 20526 27794 20578 27806
rect 28814 27794 28866 27806
rect 28926 27858 28978 27870
rect 28926 27794 28978 27806
rect 29710 27858 29762 27870
rect 29710 27794 29762 27806
rect 30382 27858 30434 27870
rect 31838 27858 31890 27870
rect 31154 27806 31166 27858
rect 31218 27806 31230 27858
rect 30382 27794 30434 27806
rect 31838 27794 31890 27806
rect 32062 27858 32114 27870
rect 32062 27794 32114 27806
rect 33406 27858 33458 27870
rect 33406 27794 33458 27806
rect 33630 27858 33682 27870
rect 33630 27794 33682 27806
rect 33742 27858 33794 27870
rect 33742 27794 33794 27806
rect 33966 27858 34018 27870
rect 33966 27794 34018 27806
rect 35086 27858 35138 27870
rect 35086 27794 35138 27806
rect 36766 27858 36818 27870
rect 36766 27794 36818 27806
rect 36990 27858 37042 27870
rect 36990 27794 37042 27806
rect 37886 27858 37938 27870
rect 39152 27896 39204 27908
rect 45502 27906 45554 27918
rect 38894 27858 38946 27870
rect 38110 27833 38162 27845
rect 38434 27806 38446 27858
rect 38498 27806 38510 27858
rect 38994 27806 39006 27858
rect 39058 27806 39070 27858
rect 39152 27832 39204 27844
rect 39902 27858 39954 27870
rect 37886 27794 37938 27806
rect 38894 27794 38946 27806
rect 39902 27794 39954 27806
rect 41358 27858 41410 27870
rect 41358 27794 41410 27806
rect 42814 27858 42866 27870
rect 42814 27794 42866 27806
rect 49310 27858 49362 27870
rect 49310 27794 49362 27806
rect 9662 27746 9714 27758
rect 25398 27746 25450 27758
rect 48246 27746 48298 27758
rect 2258 27694 2270 27746
rect 2322 27694 2334 27746
rect 11330 27694 11342 27746
rect 11394 27694 11406 27746
rect 18722 27694 18734 27746
rect 18786 27694 18798 27746
rect 19506 27694 19518 27746
rect 19570 27694 19582 27746
rect 43586 27694 43598 27746
rect 43650 27694 43662 27746
rect 9662 27682 9714 27694
rect 15486 27634 15538 27646
rect 23314 27638 23326 27690
rect 23378 27638 23390 27690
rect 25398 27682 25450 27694
rect 48246 27682 48298 27694
rect 34750 27634 34802 27646
rect 39566 27634 39618 27646
rect 16314 27582 16326 27634
rect 16378 27582 16390 27634
rect 28522 27582 28534 27634
rect 28586 27582 28598 27634
rect 33114 27582 33126 27634
rect 33178 27582 33190 27634
rect 37258 27582 37270 27634
rect 37322 27582 37334 27634
rect 15486 27570 15538 27582
rect 34750 27570 34802 27582
rect 39566 27570 39618 27582
rect 1344 27466 49616 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 49616 27466
rect 1344 27380 49616 27414
rect 14310 27298 14362 27310
rect 21366 27298 21418 27310
rect 4790 27242 4842 27254
rect 2370 27134 2382 27186
rect 2434 27134 2446 27186
rect 4274 27134 4286 27186
rect 4338 27134 4350 27186
rect 4790 27178 4842 27190
rect 10278 27242 10330 27254
rect 12842 27246 12854 27298
rect 12906 27246 12918 27298
rect 14858 27246 14870 27298
rect 14922 27246 14934 27298
rect 14310 27234 14362 27246
rect 21366 27234 21418 27246
rect 22990 27298 23042 27310
rect 48974 27298 49026 27310
rect 30762 27246 30774 27298
rect 30826 27246 30838 27298
rect 38378 27246 38390 27298
rect 38442 27246 38454 27298
rect 39386 27246 39398 27298
rect 39450 27246 39462 27298
rect 22990 27234 23042 27246
rect 48974 27234 49026 27246
rect 9762 27134 9774 27186
rect 9826 27134 9838 27186
rect 10278 27178 10330 27190
rect 16270 27186 16322 27198
rect 11666 27134 11678 27186
rect 11730 27134 11742 27186
rect 16270 27122 16322 27134
rect 17166 27186 17218 27198
rect 17166 27122 17218 27134
rect 18342 27186 18394 27198
rect 40798 27186 40850 27198
rect 24210 27134 24222 27186
rect 24274 27134 24286 27186
rect 26114 27134 26126 27186
rect 26178 27134 26190 27186
rect 32330 27134 32342 27186
rect 32394 27134 32406 27186
rect 41906 27134 41918 27186
rect 41970 27134 41982 27186
rect 18342 27122 18394 27134
rect 40798 27122 40850 27134
rect 1598 27074 1650 27086
rect 6302 27074 6354 27086
rect 4610 27022 4622 27074
rect 4674 27022 4686 27074
rect 5618 27022 5630 27074
rect 5682 27022 5694 27074
rect 6078 27035 6130 27047
rect 1598 27010 1650 27022
rect 6302 27010 6354 27022
rect 7086 27074 7138 27086
rect 11454 27074 11506 27086
rect 12462 27074 12514 27086
rect 7858 27022 7870 27074
rect 7922 27022 7934 27074
rect 10098 27022 10110 27074
rect 10162 27022 10174 27074
rect 10658 27022 10670 27074
rect 10722 27022 10734 27074
rect 11106 27022 11118 27074
rect 11170 27022 11182 27074
rect 11778 27022 11790 27074
rect 11842 27022 11854 27074
rect 7086 27010 7138 27022
rect 11454 27010 11506 27022
rect 12462 27010 12514 27022
rect 12574 27074 12626 27086
rect 15150 27074 15202 27086
rect 12574 27010 12626 27022
rect 13470 27039 13522 27051
rect 6078 26971 6130 26983
rect 13806 27046 13858 27058
rect 13470 26975 13522 26987
rect 13570 26966 13582 27018
rect 13634 26966 13646 27018
rect 13806 26982 13858 26994
rect 14030 27046 14082 27058
rect 15150 27010 15202 27022
rect 15374 27074 15426 27086
rect 15374 27010 15426 27022
rect 15598 27074 15650 27086
rect 15878 27074 15930 27086
rect 17838 27074 17890 27086
rect 19294 27074 19346 27086
rect 20414 27074 20466 27086
rect 15698 27022 15710 27074
rect 15762 27022 15774 27074
rect 17714 27022 17726 27074
rect 17778 27022 17790 27074
rect 18610 27022 18622 27074
rect 18674 27022 18686 27074
rect 15598 27010 15650 27022
rect 15878 27010 15930 27022
rect 14030 26982 14082 26994
rect 17546 26966 17558 27018
rect 17610 26966 17622 27018
rect 17838 27010 17890 27022
rect 18946 26995 18958 27047
rect 19010 26995 19022 27047
rect 20122 27022 20134 27074
rect 20186 27022 20198 27074
rect 19294 27010 19346 27022
rect 20414 27010 20466 27022
rect 20638 27074 20690 27086
rect 21870 27074 21922 27086
rect 26910 27074 26962 27086
rect 21522 27022 21534 27074
rect 21586 27022 21598 27074
rect 22734 27022 22746 27074
rect 22798 27022 22810 27074
rect 20638 27010 20690 27022
rect 21870 27010 21922 27022
rect 26910 27010 26962 27022
rect 27022 27074 27074 27086
rect 27022 27010 27074 27022
rect 27358 27074 27410 27086
rect 28366 27074 28418 27086
rect 28074 27022 28086 27074
rect 28138 27022 28150 27074
rect 27358 27010 27410 27022
rect 28366 27010 28418 27022
rect 28590 27074 28642 27086
rect 28590 27010 28642 27022
rect 29038 27074 29090 27086
rect 29038 27010 29090 27022
rect 29710 27074 29762 27086
rect 29710 27010 29762 27022
rect 31054 27074 31106 27086
rect 31054 27010 31106 27022
rect 31278 27074 31330 27086
rect 31838 27074 31890 27086
rect 31546 27022 31558 27074
rect 31610 27022 31622 27074
rect 31278 27010 31330 27022
rect 31838 27010 31890 27022
rect 31950 27074 32002 27086
rect 31950 27010 32002 27022
rect 32622 27074 32674 27086
rect 32622 27010 32674 27022
rect 32734 27074 32786 27086
rect 32734 27010 32786 27022
rect 33518 27074 33570 27086
rect 33518 27010 33570 27022
rect 33854 27074 33906 27086
rect 33854 27010 33906 27022
rect 34078 27074 34130 27086
rect 34078 27010 34130 27022
rect 34190 27074 34242 27086
rect 34750 27074 34802 27086
rect 34458 27022 34470 27074
rect 34522 27022 34534 27074
rect 34190 27010 34242 27022
rect 34750 27010 34802 27022
rect 34974 27074 35026 27086
rect 35534 27074 35586 27086
rect 35242 27022 35254 27074
rect 35306 27022 35318 27074
rect 34974 27010 35026 27022
rect 35534 27010 35586 27022
rect 37158 27074 37210 27086
rect 37158 27010 37210 27022
rect 37886 27074 37938 27086
rect 37886 27010 37938 27022
rect 38110 27074 38162 27086
rect 38110 27010 38162 27022
rect 39006 27074 39058 27086
rect 39006 27010 39058 27022
rect 39118 27074 39170 27086
rect 39118 27010 39170 27022
rect 39678 27074 39730 27086
rect 39678 27010 39730 27022
rect 40462 27074 40514 27086
rect 40462 27010 40514 27022
rect 41134 27074 41186 27086
rect 41134 27010 41186 27022
rect 44718 27074 44770 27086
rect 47742 27074 47794 27086
rect 45490 27022 45502 27074
rect 45554 27022 45566 27074
rect 44718 27010 44770 27022
rect 47742 27010 47794 27022
rect 47966 27074 48018 27086
rect 47966 27010 48018 27022
rect 49310 27074 49362 27086
rect 49310 27010 49362 27022
rect 29374 26962 29426 26974
rect 6402 26854 6414 26906
rect 6466 26854 6478 26906
rect 19394 26854 19406 26906
rect 19458 26854 19470 26906
rect 29374 26898 29426 26910
rect 36486 26962 36538 26974
rect 36486 26898 36538 26910
rect 43822 26962 43874 26974
rect 43822 26898 43874 26910
rect 47406 26962 47458 26974
rect 48234 26910 48246 26962
rect 48298 26910 48310 26962
rect 47406 26898 47458 26910
rect 30046 26850 30098 26862
rect 30046 26786 30098 26798
rect 35870 26850 35922 26862
rect 35870 26786 35922 26798
rect 37606 26850 37658 26862
rect 37606 26786 37658 26798
rect 40014 26850 40066 26862
rect 40014 26786 40066 26798
rect 1344 26682 49616 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 49616 26682
rect 1344 26596 49616 26630
rect 10278 26514 10330 26526
rect 10278 26450 10330 26462
rect 11958 26514 12010 26526
rect 11958 26450 12010 26462
rect 13302 26514 13354 26526
rect 13302 26450 13354 26462
rect 17614 26514 17666 26526
rect 17614 26450 17666 26462
rect 27190 26514 27242 26526
rect 27190 26450 27242 26462
rect 38390 26514 38442 26526
rect 38390 26450 38442 26462
rect 42086 26514 42138 26526
rect 42086 26450 42138 26462
rect 43598 26514 43650 26526
rect 43598 26450 43650 26462
rect 44214 26514 44266 26526
rect 44214 26450 44266 26462
rect 46118 26458 46170 26470
rect 21758 26402 21810 26414
rect 5674 26350 5686 26402
rect 5738 26350 5750 26402
rect 13694 26346 13746 26358
rect 2706 26238 2718 26290
rect 2770 26238 2782 26290
rect 3042 26253 3054 26305
rect 3106 26253 3118 26305
rect 5014 26290 5066 26302
rect 5014 26226 5066 26238
rect 5182 26290 5234 26302
rect 5182 26226 5234 26238
rect 5406 26290 5458 26302
rect 5406 26226 5458 26238
rect 5966 26290 6018 26302
rect 6962 26282 6974 26334
rect 7026 26282 7038 26334
rect 7186 26238 7198 26290
rect 7250 26238 7262 26290
rect 8306 26282 8318 26334
rect 8370 26282 8382 26334
rect 9998 26290 10050 26302
rect 8642 26238 8654 26290
rect 8706 26238 8718 26290
rect 10098 26238 10110 26290
rect 10162 26238 10174 26290
rect 10882 26238 10894 26290
rect 10946 26238 10958 26290
rect 11106 26282 11118 26334
rect 11170 26282 11182 26334
rect 12238 26290 12290 26302
rect 21758 26338 21810 26350
rect 26070 26402 26122 26414
rect 11778 26238 11790 26290
rect 11842 26238 11854 26290
rect 13458 26238 13470 26290
rect 13522 26238 13534 26290
rect 13694 26282 13746 26294
rect 13806 26318 13858 26330
rect 13806 26254 13858 26266
rect 14086 26325 14138 26337
rect 14086 26261 14138 26273
rect 14254 26318 14306 26330
rect 14254 26254 14306 26266
rect 14534 26290 14586 26302
rect 5966 26226 6018 26238
rect 9998 26226 10050 26238
rect 12238 26226 12290 26238
rect 14534 26226 14586 26238
rect 14814 26290 14866 26302
rect 14814 26226 14866 26238
rect 17278 26290 17330 26302
rect 17278 26226 17330 26238
rect 17950 26290 18002 26302
rect 17950 26226 18002 26238
rect 19070 26290 19122 26302
rect 22306 26238 22318 26290
rect 22370 26238 22382 26290
rect 23046 26276 23058 26328
rect 23110 26276 23122 26328
rect 25230 26325 25282 26337
rect 24726 26290 24778 26302
rect 25330 26294 25342 26346
rect 25394 26294 25406 26346
rect 25622 26325 25674 26337
rect 25230 26261 25282 26273
rect 25778 26294 25790 26346
rect 25842 26294 25854 26346
rect 26070 26338 26122 26350
rect 30270 26402 30322 26414
rect 30270 26338 30322 26350
rect 32286 26402 32338 26414
rect 31726 26328 31778 26340
rect 32286 26338 32338 26350
rect 34638 26402 34690 26414
rect 25622 26261 25674 26273
rect 26910 26290 26962 26302
rect 27582 26290 27634 26302
rect 19070 26226 19122 26238
rect 24726 26226 24778 26238
rect 27010 26238 27022 26290
rect 27074 26238 27086 26290
rect 28354 26238 28366 26290
rect 28418 26238 28430 26290
rect 31378 26238 31390 26290
rect 31442 26238 31454 26290
rect 34078 26328 34130 26340
rect 34638 26338 34690 26350
rect 35310 26402 35362 26414
rect 40182 26402 40234 26414
rect 35310 26338 35362 26350
rect 39118 26346 39170 26358
rect 31726 26264 31778 26276
rect 33182 26290 33234 26302
rect 26910 26226 26962 26238
rect 27582 26226 27634 26238
rect 32454 26234 32506 26246
rect 15766 26178 15818 26190
rect 3154 26126 3166 26178
rect 3218 26126 3230 26178
rect 6850 26126 6862 26178
rect 6914 26126 6926 26178
rect 8194 26126 8206 26178
rect 8258 26126 8270 26178
rect 11218 26126 11230 26178
rect 11282 26126 11294 26178
rect 15766 26114 15818 26126
rect 16662 26178 16714 26190
rect 24278 26178 24330 26190
rect 19842 26126 19854 26178
rect 19906 26126 19918 26178
rect 16662 26114 16714 26126
rect 6302 26066 6354 26078
rect 6302 26002 6354 26014
rect 9662 26066 9714 26078
rect 9662 26002 9714 26014
rect 12574 26066 12626 26078
rect 12574 26002 12626 26014
rect 15150 26066 15202 26078
rect 15150 26002 15202 26014
rect 18286 26066 18338 26078
rect 22530 26070 22542 26122
rect 22594 26070 22606 26122
rect 24278 26114 24330 26126
rect 30886 26178 30938 26190
rect 31602 26182 31614 26234
rect 31666 26182 31678 26234
rect 33182 26226 33234 26238
rect 33294 26290 33346 26302
rect 37998 26290 38050 26302
rect 34078 26264 34130 26276
rect 33294 26226 33346 26238
rect 34806 26234 34858 26246
rect 37202 26238 37214 26290
rect 37266 26238 37278 26290
rect 39118 26282 39170 26294
rect 39342 26346 39394 26358
rect 46118 26394 46170 26406
rect 39342 26282 39394 26294
rect 39454 26318 39506 26330
rect 39454 26254 39506 26266
rect 39734 26325 39786 26337
rect 39890 26294 39902 26346
rect 39954 26294 39966 26346
rect 40182 26338 40234 26350
rect 39734 26261 39786 26273
rect 41134 26290 41186 26302
rect 33954 26182 33966 26234
rect 34018 26182 34030 26234
rect 37998 26226 38050 26238
rect 41134 26226 41186 26238
rect 43262 26290 43314 26302
rect 43262 26226 43314 26238
rect 44942 26290 44994 26302
rect 45098 26294 45110 26346
rect 45162 26294 45174 26346
rect 47966 26328 48018 26340
rect 45390 26290 45442 26302
rect 45266 26238 45278 26290
rect 45330 26238 45342 26290
rect 46274 26238 46286 26290
rect 46338 26238 46350 26290
rect 44942 26226 44994 26238
rect 45390 26226 45442 26238
rect 47238 26234 47290 26246
rect 47618 26238 47630 26290
rect 47682 26238 47694 26290
rect 47966 26264 48018 26276
rect 49198 26290 49250 26302
rect 32454 26170 32506 26182
rect 34806 26170 34858 26182
rect 42534 26178 42586 26190
rect 30886 26114 30938 26126
rect 49198 26226 49250 26238
rect 47238 26170 47290 26182
rect 47406 26178 47458 26190
rect 42534 26114 42586 26126
rect 47406 26114 47458 26126
rect 18286 26002 18338 26014
rect 26574 26066 26626 26078
rect 26574 26002 26626 26014
rect 31222 26066 31274 26078
rect 38782 26066 38834 26078
rect 33562 26014 33574 26066
rect 33626 26014 33638 26066
rect 31222 26002 31274 26014
rect 38782 26002 38834 26014
rect 41470 26066 41522 26078
rect 41470 26002 41522 26014
rect 45670 26066 45722 26078
rect 45670 26002 45722 26014
rect 48862 26066 48914 26078
rect 48862 26002 48914 26014
rect 1344 25898 49616 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 49616 25898
rect 1344 25812 49616 25846
rect 11510 25730 11562 25742
rect 11510 25666 11562 25678
rect 20302 25730 20354 25742
rect 20302 25666 20354 25678
rect 21702 25730 21754 25742
rect 21702 25666 21754 25678
rect 37438 25730 37490 25742
rect 37438 25666 37490 25678
rect 38950 25730 39002 25742
rect 38950 25666 39002 25678
rect 44886 25730 44938 25742
rect 44886 25666 44938 25678
rect 28254 25618 28306 25630
rect 32790 25618 32842 25630
rect 44326 25618 44378 25630
rect 3714 25566 3726 25618
rect 3778 25566 3790 25618
rect 9090 25566 9102 25618
rect 9154 25566 9166 25618
rect 10994 25566 11006 25618
rect 11058 25566 11070 25618
rect 13906 25566 13918 25618
rect 13970 25566 13982 25618
rect 15810 25566 15822 25618
rect 15874 25566 15886 25618
rect 17714 25566 17726 25618
rect 17778 25566 17790 25618
rect 19618 25566 19630 25618
rect 19682 25566 19694 25618
rect 23426 25566 23438 25618
rect 23490 25566 23502 25618
rect 25330 25566 25342 25618
rect 25394 25566 25406 25618
rect 29810 25566 29822 25618
rect 29874 25566 29886 25618
rect 40002 25566 40014 25618
rect 40066 25566 40078 25618
rect 28254 25554 28306 25566
rect 32790 25554 32842 25566
rect 44326 25554 44378 25566
rect 46062 25618 46114 25630
rect 46610 25566 46622 25618
rect 46674 25566 46686 25618
rect 48514 25566 48526 25618
rect 48578 25566 48590 25618
rect 46062 25554 46114 25566
rect 4510 25506 4562 25518
rect 4510 25442 4562 25454
rect 5854 25506 5906 25518
rect 7982 25506 8034 25518
rect 5854 25442 5906 25454
rect 6178 25427 6190 25479
rect 6242 25427 6254 25479
rect 6402 25454 6414 25506
rect 6466 25454 6478 25506
rect 7982 25442 8034 25454
rect 8318 25506 8370 25518
rect 16606 25506 16658 25518
rect 8318 25442 8370 25454
rect 11790 25478 11842 25490
rect 12238 25478 12290 25490
rect 11790 25414 11842 25426
rect 1822 25394 1874 25406
rect 12002 25398 12014 25450
rect 12066 25398 12078 25450
rect 12238 25414 12290 25426
rect 12350 25450 12402 25462
rect 16606 25442 16658 25454
rect 16942 25506 16994 25518
rect 16942 25442 16994 25454
rect 19966 25506 20018 25518
rect 23102 25506 23154 25518
rect 21858 25454 21870 25506
rect 21922 25454 21934 25506
rect 19966 25442 20018 25454
rect 23102 25442 23154 25454
rect 26126 25506 26178 25518
rect 29038 25506 29090 25518
rect 34750 25506 34802 25518
rect 26338 25454 26350 25506
rect 26402 25454 26414 25506
rect 26126 25442 26178 25454
rect 27794 25426 27806 25478
rect 27858 25426 27870 25478
rect 28018 25454 28030 25506
rect 28082 25454 28094 25506
rect 28422 25450 28474 25462
rect 12350 25386 12402 25398
rect 33842 25454 33854 25506
rect 33906 25454 33918 25506
rect 34190 25468 34242 25480
rect 29038 25442 29090 25454
rect 34514 25454 34526 25506
rect 34578 25454 34590 25506
rect 35086 25506 35138 25518
rect 34750 25442 34802 25454
rect 34918 25450 34970 25462
rect 28422 25386 28474 25398
rect 31726 25394 31778 25406
rect 34190 25404 34242 25416
rect 1822 25330 1874 25342
rect 35086 25442 35138 25454
rect 35310 25506 35362 25518
rect 35870 25506 35922 25518
rect 35578 25454 35590 25506
rect 35642 25454 35654 25506
rect 35310 25442 35362 25454
rect 35870 25442 35922 25454
rect 37774 25506 37826 25518
rect 39230 25506 39282 25518
rect 37774 25442 37826 25454
rect 38110 25471 38162 25483
rect 38502 25471 38554 25483
rect 38110 25407 38162 25419
rect 38210 25398 38222 25450
rect 38274 25398 38286 25450
rect 38502 25407 38554 25419
rect 38670 25478 38722 25490
rect 39230 25442 39282 25454
rect 41918 25506 41970 25518
rect 41918 25442 41970 25454
rect 42590 25506 42642 25518
rect 49310 25506 49362 25518
rect 43454 25454 43466 25506
rect 43518 25454 43530 25506
rect 44706 25454 44718 25506
rect 44770 25454 44782 25506
rect 45826 25454 45838 25506
rect 45890 25454 45902 25506
rect 42590 25442 42642 25454
rect 46230 25450 46282 25462
rect 38670 25414 38722 25426
rect 34918 25386 34970 25398
rect 43710 25394 43762 25406
rect 45602 25398 45614 25450
rect 45666 25398 45678 25450
rect 49310 25442 49362 25454
rect 5954 25286 5966 25338
rect 6018 25286 6030 25338
rect 31726 25330 31778 25342
rect 46230 25386 46282 25398
rect 43710 25330 43762 25342
rect 12854 25282 12906 25294
rect 12854 25218 12906 25230
rect 22766 25282 22818 25294
rect 22766 25218 22818 25230
rect 32342 25282 32394 25294
rect 32342 25218 32394 25230
rect 33350 25282 33402 25294
rect 33350 25218 33402 25230
rect 33686 25282 33738 25294
rect 33686 25218 33738 25230
rect 36206 25282 36258 25294
rect 36206 25218 36258 25230
rect 1344 25114 49616 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 49616 25114
rect 1344 25028 49616 25062
rect 15262 24946 15314 24958
rect 15262 24882 15314 24894
rect 29038 24946 29090 24958
rect 29038 24882 29090 24894
rect 33182 24946 33234 24958
rect 33182 24882 33234 24894
rect 34246 24946 34298 24958
rect 34246 24882 34298 24894
rect 3950 24834 4002 24846
rect 5406 24834 5458 24846
rect 4554 24782 4566 24834
rect 4618 24782 4630 24834
rect 35310 24834 35362 24846
rect 3950 24770 4002 24782
rect 5406 24770 5458 24782
rect 11006 24778 11058 24790
rect 40294 24834 40346 24846
rect 2830 24722 2882 24734
rect 4846 24722 4898 24734
rect 3694 24670 3706 24722
rect 3758 24670 3770 24722
rect 2830 24658 2882 24670
rect 4846 24658 4898 24670
rect 5070 24722 5122 24734
rect 8094 24722 8146 24734
rect 7298 24670 7310 24722
rect 7362 24670 7374 24722
rect 5070 24658 5122 24670
rect 8094 24658 8146 24670
rect 9102 24722 9154 24734
rect 9102 24658 9154 24670
rect 10166 24722 10218 24734
rect 10434 24726 10446 24778
rect 10498 24726 10510 24778
rect 10658 24726 10670 24778
rect 10722 24726 10734 24778
rect 10882 24726 10894 24778
rect 10946 24726 10958 24778
rect 11006 24714 11058 24726
rect 11230 24722 11282 24734
rect 10166 24658 10218 24670
rect 12002 24670 12014 24722
rect 12066 24670 12078 24722
rect 14466 24714 14478 24766
rect 14530 24714 14542 24766
rect 15598 24722 15650 24734
rect 14690 24670 14702 24722
rect 14754 24670 14766 24722
rect 11230 24658 11282 24670
rect 15598 24658 15650 24670
rect 16494 24722 16546 24734
rect 18174 24722 18226 24734
rect 16594 24670 16606 24722
rect 16658 24670 16670 24722
rect 17378 24670 17390 24722
rect 17442 24670 17454 24722
rect 17714 24670 17726 24722
rect 17778 24670 17790 24722
rect 16494 24658 16546 24670
rect 18174 24658 18226 24670
rect 18286 24722 18338 24734
rect 21074 24697 21086 24749
rect 21138 24697 21150 24749
rect 21758 24722 21810 24734
rect 25118 24722 25170 24734
rect 18286 24658 18338 24670
rect 22530 24670 22542 24722
rect 22594 24670 22606 24722
rect 25890 24670 25902 24722
rect 25954 24670 25966 24722
rect 30706 24697 30718 24749
rect 30770 24697 30782 24749
rect 31397 24726 31409 24778
rect 31461 24726 31473 24778
rect 35310 24770 35362 24782
rect 39454 24778 39506 24790
rect 32286 24722 32338 24734
rect 21758 24658 21810 24670
rect 25118 24658 25170 24670
rect 32286 24658 32338 24670
rect 33518 24722 33570 24734
rect 37998 24722 38050 24734
rect 38490 24726 38502 24778
rect 38554 24726 38566 24778
rect 34066 24670 34078 24722
rect 34130 24670 34142 24722
rect 37202 24670 37214 24722
rect 37266 24670 37278 24722
rect 38210 24670 38222 24722
rect 38274 24670 38286 24722
rect 39454 24714 39506 24726
rect 39566 24750 39618 24762
rect 39566 24686 39618 24698
rect 39846 24757 39898 24769
rect 40002 24726 40014 24778
rect 40066 24726 40078 24778
rect 40294 24770 40346 24782
rect 43822 24834 43874 24846
rect 49130 24782 49142 24834
rect 49194 24782 49206 24834
rect 43822 24770 43874 24782
rect 44568 24760 44620 24772
rect 39846 24693 39898 24705
rect 41134 24722 41186 24734
rect 44270 24722 44322 24734
rect 41906 24670 41918 24722
rect 41970 24670 41982 24722
rect 44370 24670 44382 24722
rect 44434 24670 44446 24722
rect 44568 24696 44620 24708
rect 45838 24722 45890 24734
rect 33518 24658 33570 24670
rect 37998 24658 38050 24670
rect 41134 24658 41186 24670
rect 44270 24658 44322 24670
rect 45838 24658 45890 24670
rect 45950 24722 46002 24734
rect 46946 24670 46958 24722
rect 47010 24670 47022 24722
rect 47282 24697 47294 24749
rect 47346 24697 47358 24749
rect 47630 24722 47682 24734
rect 45950 24658 46002 24670
rect 47630 24658 47682 24670
rect 47966 24722 48018 24734
rect 47966 24658 48018 24670
rect 48638 24722 48690 24734
rect 48638 24658 48690 24670
rect 48862 24722 48914 24734
rect 48862 24658 48914 24670
rect 33910 24610 33962 24622
rect 13906 24558 13918 24610
rect 13970 24558 13982 24610
rect 14354 24558 14366 24610
rect 14418 24558 14430 24610
rect 24434 24558 24446 24610
rect 24498 24558 24510 24610
rect 27794 24558 27806 24610
rect 27858 24558 27870 24610
rect 8766 24498 8818 24510
rect 8766 24434 8818 24446
rect 16158 24498 16210 24510
rect 17602 24502 17614 24554
rect 17666 24502 17678 24554
rect 33910 24546 33962 24558
rect 34918 24610 34970 24622
rect 39174 24610 39226 24622
rect 38658 24558 38670 24610
rect 38722 24558 38734 24610
rect 34918 24546 34970 24558
rect 39174 24546 39226 24558
rect 45558 24610 45610 24622
rect 47058 24558 47070 24610
rect 47122 24558 47134 24610
rect 45558 24546 45610 24558
rect 20414 24498 20466 24510
rect 18554 24446 18566 24498
rect 18618 24446 18630 24498
rect 16158 24434 16210 24446
rect 20414 24434 20466 24446
rect 31166 24498 31218 24510
rect 31166 24434 31218 24446
rect 44942 24498 44994 24510
rect 46218 24446 46230 24498
rect 46282 24446 46294 24498
rect 44942 24434 44994 24446
rect 1344 24330 49616 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 49616 24330
rect 1344 24244 49616 24278
rect 12070 24162 12122 24174
rect 12070 24098 12122 24110
rect 16998 24162 17050 24174
rect 26854 24162 26906 24174
rect 34974 24162 35026 24174
rect 23930 24110 23942 24162
rect 23994 24110 24006 24162
rect 28522 24110 28534 24162
rect 28586 24110 28598 24162
rect 16998 24098 17050 24110
rect 26854 24098 26906 24110
rect 34974 24098 35026 24110
rect 35758 24162 35810 24174
rect 35758 24098 35810 24110
rect 37102 24162 37154 24174
rect 37102 24098 37154 24110
rect 37774 24162 37826 24174
rect 37774 24098 37826 24110
rect 5966 24050 6018 24062
rect 13582 24050 13634 24062
rect 8642 23998 8654 24050
rect 8706 23998 8718 24050
rect 10546 23998 10558 24050
rect 10610 23998 10622 24050
rect 5966 23986 6018 23998
rect 13582 23986 13634 23998
rect 14646 24050 14698 24062
rect 14646 23986 14698 23998
rect 15094 24050 15146 24062
rect 15094 23986 15146 23998
rect 15542 24050 15594 24062
rect 15542 23986 15594 23998
rect 15990 24050 16042 24062
rect 15990 23986 16042 23998
rect 25734 24050 25786 24062
rect 34582 24050 34634 24062
rect 45502 24050 45554 24062
rect 34066 23998 34078 24050
rect 34130 23998 34142 24050
rect 40226 23998 40238 24050
rect 40290 23998 40302 24050
rect 25734 23986 25786 23998
rect 34582 23986 34634 23998
rect 45502 23986 45554 23998
rect 1598 23938 1650 23950
rect 6302 23938 6354 23950
rect 2370 23886 2382 23938
rect 2434 23886 2446 23938
rect 5618 23886 5630 23938
rect 5682 23886 5694 23938
rect 6078 23899 6130 23911
rect 1598 23874 1650 23886
rect 6302 23874 6354 23886
rect 6638 23938 6690 23950
rect 6638 23874 6690 23886
rect 7870 23938 7922 23950
rect 13918 23938 13970 23950
rect 7870 23874 7922 23886
rect 12350 23910 12402 23922
rect 4286 23826 4338 23838
rect 6078 23835 6130 23847
rect 12350 23846 12402 23858
rect 12574 23910 12626 23922
rect 12574 23846 12626 23858
rect 12798 23910 12850 23922
rect 12798 23846 12850 23858
rect 12910 23882 12962 23894
rect 4286 23762 4338 23774
rect 11734 23826 11786 23838
rect 13918 23874 13970 23886
rect 16718 23938 16770 23950
rect 16718 23874 16770 23886
rect 17278 23938 17330 23950
rect 17278 23874 17330 23886
rect 17726 23938 17778 23950
rect 12910 23818 12962 23830
rect 16382 23826 16434 23838
rect 11734 23762 11786 23774
rect 16382 23762 16434 23774
rect 17390 23826 17442 23838
rect 17546 23830 17558 23882
rect 17610 23830 17622 23882
rect 17726 23874 17778 23886
rect 17950 23938 18002 23950
rect 21758 23938 21810 23950
rect 18722 23886 18734 23938
rect 18786 23886 18798 23938
rect 17950 23874 18002 23886
rect 21758 23874 21810 23886
rect 22430 23938 22482 23950
rect 23550 23938 23602 23950
rect 22661 23886 22673 23938
rect 22725 23886 22737 23938
rect 22430 23874 22482 23886
rect 23550 23874 23602 23886
rect 24222 23938 24274 23950
rect 24222 23874 24274 23886
rect 24446 23938 24498 23950
rect 27134 23938 27186 23950
rect 24446 23874 24498 23886
rect 25946 23870 25958 23922
rect 26010 23870 26022 23922
rect 26574 23910 26626 23922
rect 17390 23762 17442 23774
rect 20638 23826 20690 23838
rect 26114 23830 26126 23882
rect 26178 23830 26190 23882
rect 26338 23830 26350 23882
rect 26402 23830 26414 23882
rect 27134 23874 27186 23886
rect 27358 23938 27410 23950
rect 27358 23874 27410 23886
rect 28142 23938 28194 23950
rect 28142 23874 28194 23886
rect 28254 23938 28306 23950
rect 28254 23874 28306 23886
rect 29038 23938 29090 23950
rect 32622 23938 32674 23950
rect 29810 23886 29822 23938
rect 29874 23886 29886 23938
rect 29038 23874 29090 23886
rect 32622 23874 32674 23886
rect 33294 23938 33346 23950
rect 35310 23938 35362 23950
rect 33618 23886 33630 23938
rect 33682 23886 33694 23938
rect 33910 23908 33962 23920
rect 33294 23874 33346 23886
rect 26574 23846 26626 23858
rect 35310 23874 35362 23886
rect 35422 23938 35474 23950
rect 35422 23874 35474 23886
rect 37438 23938 37490 23950
rect 37438 23874 37490 23886
rect 38110 23938 38162 23950
rect 39454 23938 39506 23950
rect 38446 23910 38498 23922
rect 38110 23874 38162 23886
rect 38334 23882 38386 23894
rect 33910 23844 33962 23856
rect 31726 23826 31778 23838
rect 27626 23774 27638 23826
rect 27690 23774 27702 23826
rect 38446 23846 38498 23858
rect 38670 23910 38722 23922
rect 38670 23846 38722 23858
rect 38882 23830 38894 23882
rect 38946 23830 38958 23882
rect 39454 23874 39506 23886
rect 42478 23938 42530 23950
rect 42478 23874 42530 23886
rect 42702 23938 42754 23950
rect 44830 23938 44882 23950
rect 45108 23938 45160 23950
rect 42970 23886 42982 23938
rect 43034 23886 43046 23938
rect 44034 23886 44046 23938
rect 44098 23886 44110 23938
rect 44930 23886 44942 23938
rect 44994 23886 45006 23938
rect 42702 23874 42754 23886
rect 44830 23874 44882 23886
rect 45108 23874 45160 23886
rect 46734 23938 46786 23950
rect 47630 23938 47682 23950
rect 46946 23886 46958 23938
rect 47010 23886 47022 23938
rect 46734 23874 46786 23886
rect 38334 23818 38386 23830
rect 39174 23826 39226 23838
rect 20638 23762 20690 23774
rect 31726 23762 31778 23774
rect 39174 23762 39226 23774
rect 42142 23826 42194 23838
rect 47394 23830 47406 23882
rect 47458 23830 47470 23882
rect 47630 23874 47682 23886
rect 48078 23938 48130 23950
rect 48078 23874 48130 23886
rect 48302 23938 48354 23950
rect 48570 23886 48582 23938
rect 48634 23886 48646 23938
rect 48302 23874 48354 23886
rect 42142 23762 42194 23774
rect 44214 23770 44266 23782
rect 21422 23714 21474 23726
rect 21422 23650 21474 23662
rect 32286 23714 32338 23726
rect 32286 23650 32338 23662
rect 32958 23714 33010 23726
rect 32958 23650 33010 23662
rect 36374 23714 36426 23726
rect 36374 23650 36426 23662
rect 43542 23714 43594 23726
rect 44214 23706 44266 23718
rect 46398 23714 46450 23726
rect 47730 23718 47742 23770
rect 47794 23718 47806 23770
rect 43542 23650 43594 23662
rect 46398 23650 46450 23662
rect 1344 23546 49616 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 49616 23546
rect 1344 23460 49616 23494
rect 2382 23378 2434 23390
rect 2382 23314 2434 23326
rect 7870 23378 7922 23390
rect 3602 23270 3614 23322
rect 3666 23270 3678 23322
rect 7870 23314 7922 23326
rect 9662 23378 9714 23390
rect 9662 23314 9714 23326
rect 13190 23378 13242 23390
rect 13190 23314 13242 23326
rect 18790 23378 18842 23390
rect 18790 23314 18842 23326
rect 19294 23378 19346 23390
rect 25398 23378 25450 23390
rect 19294 23314 19346 23326
rect 20918 23322 20970 23334
rect 11398 23266 11450 23278
rect 5338 23214 5350 23266
rect 5402 23214 5414 23266
rect 18174 23266 18226 23278
rect 11398 23202 11450 23214
rect 12574 23210 12626 23222
rect 11958 23189 12010 23201
rect 2718 23154 2770 23166
rect 3490 23102 3502 23154
rect 3554 23102 3566 23154
rect 3826 23129 3838 23181
rect 3890 23129 3902 23181
rect 4174 23154 4226 23166
rect 2718 23090 2770 23102
rect 4174 23090 4226 23102
rect 4846 23154 4898 23166
rect 4846 23090 4898 23102
rect 5070 23154 5122 23166
rect 5730 23102 5742 23154
rect 5794 23102 5806 23154
rect 6066 23117 6078 23169
rect 6130 23117 6142 23169
rect 6850 23129 6862 23181
rect 6914 23129 6926 23181
rect 9998 23154 10050 23166
rect 5070 23090 5122 23102
rect 9998 23090 10050 23102
rect 10838 23154 10890 23166
rect 11958 23125 12010 23137
rect 12238 23182 12290 23194
rect 12238 23118 12290 23130
rect 12462 23182 12514 23194
rect 17614 23210 17666 23222
rect 12574 23146 12626 23158
rect 13358 23154 13410 23166
rect 12462 23118 12514 23130
rect 10838 23090 10890 23102
rect 13358 23090 13410 23102
rect 14590 23154 14642 23166
rect 14590 23090 14642 23102
rect 15262 23154 15314 23166
rect 15262 23090 15314 23102
rect 16494 23154 16546 23166
rect 25398 23314 25450 23326
rect 34470 23378 34522 23390
rect 34470 23314 34522 23326
rect 34918 23378 34970 23390
rect 34918 23314 34970 23326
rect 38334 23378 38386 23390
rect 38334 23314 38386 23326
rect 40406 23378 40458 23390
rect 40406 23314 40458 23326
rect 20918 23258 20970 23270
rect 44718 23266 44770 23278
rect 18174 23202 18226 23214
rect 18342 23210 18394 23222
rect 26649 23210 26701 23222
rect 30158 23210 30210 23222
rect 32585 23210 32637 23222
rect 17614 23146 17666 23158
rect 26014 23182 26066 23194
rect 18342 23146 18394 23158
rect 18958 23154 19010 23166
rect 16494 23090 16546 23102
rect 10390 23042 10442 23054
rect 6178 22990 6190 23042
rect 6242 22990 6254 23042
rect 10390 22978 10442 22990
rect 15094 23042 15146 23054
rect 15094 22978 15146 22990
rect 16886 23042 16938 23054
rect 17490 23046 17502 23098
rect 17554 23046 17566 23098
rect 18958 23090 19010 23102
rect 19910 23154 19962 23166
rect 24782 23154 24834 23166
rect 21074 23102 21086 23154
rect 21138 23102 21150 23154
rect 19910 23090 19962 23102
rect 24782 23090 24834 23102
rect 25734 23154 25786 23166
rect 26226 23158 26238 23210
rect 26290 23158 26302 23210
rect 26406 23189 26458 23201
rect 26014 23118 26066 23130
rect 26649 23146 26701 23158
rect 26798 23154 26850 23166
rect 26406 23125 26458 23137
rect 25734 23090 25786 23102
rect 26798 23090 26850 23102
rect 27022 23154 27074 23166
rect 27794 23102 27806 23154
rect 27858 23102 27870 23154
rect 28130 23146 28142 23198
rect 28194 23146 28206 23198
rect 28702 23154 28754 23166
rect 27022 23090 27074 23102
rect 28702 23090 28754 23102
rect 29038 23154 29090 23166
rect 29038 23090 29090 23102
rect 29318 23154 29370 23166
rect 29586 23158 29598 23210
rect 29650 23158 29662 23210
rect 29810 23158 29822 23210
rect 29874 23158 29886 23210
rect 30034 23158 30046 23210
rect 30098 23158 30110 23210
rect 31950 23182 32002 23194
rect 30158 23146 30210 23158
rect 31166 23154 31218 23166
rect 29318 23090 29370 23102
rect 31166 23090 31218 23102
rect 31278 23154 31330 23166
rect 31278 23090 31330 23102
rect 31670 23154 31722 23166
rect 32162 23158 32174 23210
rect 32226 23158 32238 23210
rect 32386 23158 32398 23210
rect 32450 23158 32462 23210
rect 32585 23146 32637 23158
rect 32958 23154 33010 23166
rect 31950 23118 32002 23130
rect 31670 23090 31722 23102
rect 32958 23090 33010 23102
rect 33910 23154 33962 23166
rect 33910 23090 33962 23102
rect 37998 23154 38050 23166
rect 37998 23090 38050 23102
rect 38670 23154 38722 23166
rect 38670 23090 38722 23102
rect 39006 23154 39058 23166
rect 41234 23129 41246 23181
rect 41298 23129 41310 23181
rect 44046 23154 44098 23166
rect 44538 23158 44550 23210
rect 44602 23158 44614 23210
rect 44718 23202 44770 23214
rect 48078 23266 48130 23278
rect 48078 23202 48130 23214
rect 45390 23154 45442 23166
rect 39006 23090 39058 23102
rect 44930 23102 44942 23154
rect 44994 23102 45006 23154
rect 44046 23090 44098 23102
rect 45390 23090 45442 23102
rect 48638 23154 48690 23166
rect 48638 23090 48690 23102
rect 16886 22978 16938 22990
rect 21926 23042 21978 23054
rect 39958 23042 40010 23054
rect 48974 23042 49026 23054
rect 28242 22990 28254 23042
rect 28306 22990 28318 23042
rect 35298 22990 35310 23042
rect 35362 22990 35374 23042
rect 37202 22990 37214 23042
rect 37266 22990 37278 23042
rect 46162 22990 46174 23042
rect 46226 22990 46238 23042
rect 21926 22978 21978 22990
rect 39958 22978 40010 22990
rect 48974 22978 49026 22990
rect 11734 22930 11786 22942
rect 11734 22866 11786 22878
rect 13694 22930 13746 22942
rect 13694 22866 13746 22878
rect 14254 22930 14306 22942
rect 14254 22866 14306 22878
rect 15598 22930 15650 22942
rect 15598 22866 15650 22878
rect 16158 22930 16210 22942
rect 16158 22866 16210 22878
rect 24446 22930 24498 22942
rect 33294 22930 33346 22942
rect 27290 22878 27302 22930
rect 27354 22878 27366 22930
rect 30874 22878 30886 22930
rect 30938 22878 30950 22930
rect 24446 22866 24498 22878
rect 33294 22866 33346 22878
rect 39342 22930 39394 22942
rect 39342 22866 39394 22878
rect 41918 22930 41970 22942
rect 41918 22866 41970 22878
rect 43804 22930 43856 22942
rect 43804 22866 43856 22878
rect 45110 22930 45162 22942
rect 45110 22866 45162 22878
rect 1344 22762 49616 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 49616 22762
rect 1344 22676 49616 22710
rect 13526 22594 13578 22606
rect 3434 22542 3446 22594
rect 3498 22542 3510 22594
rect 13526 22530 13578 22542
rect 37214 22594 37266 22606
rect 37214 22530 37266 22542
rect 45950 22594 46002 22606
rect 45950 22530 46002 22542
rect 26854 22482 26906 22494
rect 4274 22430 4286 22482
rect 4338 22430 4350 22482
rect 6626 22430 6638 22482
rect 6690 22430 6702 22482
rect 15698 22430 15710 22482
rect 15762 22430 15774 22482
rect 23986 22430 23998 22482
rect 24050 22430 24062 22482
rect 25890 22430 25902 22482
rect 25954 22430 25966 22482
rect 26854 22418 26906 22430
rect 29318 22482 29370 22494
rect 31154 22430 31166 22482
rect 31218 22430 31230 22482
rect 33058 22430 33070 22482
rect 33122 22430 33134 22482
rect 38994 22430 39006 22482
rect 39058 22430 39070 22482
rect 40898 22430 40910 22482
rect 40962 22430 40974 22482
rect 29318 22418 29370 22430
rect 2270 22370 2322 22382
rect 2270 22306 2322 22318
rect 2382 22370 2434 22382
rect 2382 22306 2434 22318
rect 3054 22370 3106 22382
rect 3054 22306 3106 22318
rect 3166 22370 3218 22382
rect 4958 22370 5010 22382
rect 3938 22318 3950 22370
rect 4002 22318 4014 22370
rect 3166 22306 3218 22318
rect 4162 22274 4174 22326
rect 4226 22274 4238 22326
rect 4958 22306 5010 22318
rect 5182 22370 5234 22382
rect 5182 22306 5234 22318
rect 5854 22370 5906 22382
rect 5854 22306 5906 22318
rect 8878 22370 8930 22382
rect 11566 22370 11618 22382
rect 9650 22318 9662 22370
rect 9714 22318 9726 22370
rect 14926 22370 14978 22382
rect 8878 22306 8930 22318
rect 11566 22306 11618 22318
rect 12350 22342 12402 22354
rect 12798 22342 12850 22354
rect 12350 22278 12402 22290
rect 8542 22258 8594 22270
rect 2650 22206 2662 22258
rect 2714 22206 2726 22258
rect 4666 22206 4678 22258
rect 4730 22206 4742 22258
rect 8542 22194 8594 22206
rect 12070 22258 12122 22270
rect 12562 22262 12574 22314
rect 12626 22262 12638 22314
rect 12798 22278 12850 22290
rect 12910 22335 12962 22347
rect 14254 22342 14306 22354
rect 12910 22271 12962 22283
rect 13794 22262 13806 22314
rect 13858 22262 13870 22314
rect 14018 22262 14030 22314
rect 14082 22262 14094 22314
rect 14254 22278 14306 22290
rect 14366 22314 14418 22326
rect 14926 22306 14978 22318
rect 18510 22370 18562 22382
rect 18510 22306 18562 22318
rect 18734 22370 18786 22382
rect 19294 22370 19346 22382
rect 19002 22318 19014 22370
rect 19066 22318 19078 22370
rect 18734 22306 18786 22318
rect 19294 22306 19346 22318
rect 20862 22370 20914 22382
rect 20862 22306 20914 22318
rect 21422 22370 21474 22382
rect 21422 22306 21474 22318
rect 23214 22370 23266 22382
rect 29486 22370 29538 22382
rect 23214 22306 23266 22318
rect 27918 22342 27970 22354
rect 28478 22335 28530 22347
rect 27918 22278 27970 22290
rect 14366 22250 14418 22262
rect 17614 22258 17666 22270
rect 12070 22194 12122 22206
rect 17614 22194 17666 22206
rect 27638 22258 27690 22270
rect 28130 22262 28142 22314
rect 28194 22262 28206 22314
rect 28354 22262 28366 22314
rect 28418 22262 28430 22314
rect 29486 22306 29538 22318
rect 29710 22370 29762 22382
rect 29710 22306 29762 22318
rect 33854 22370 33906 22382
rect 36150 22370 36202 22382
rect 33854 22306 33906 22318
rect 34638 22342 34690 22354
rect 28478 22271 28530 22283
rect 34134 22258 34186 22270
rect 34402 22262 34414 22314
rect 34466 22262 34478 22314
rect 34638 22278 34690 22290
rect 34862 22342 34914 22354
rect 34862 22278 34914 22290
rect 34974 22335 35026 22347
rect 35242 22302 35254 22354
rect 35306 22302 35318 22354
rect 35422 22342 35474 22354
rect 34974 22271 35026 22283
rect 35422 22278 35474 22290
rect 35646 22342 35698 22354
rect 35646 22278 35698 22290
rect 35858 22262 35870 22314
rect 35922 22262 35934 22314
rect 36150 22306 36202 22318
rect 36878 22370 36930 22382
rect 36878 22306 36930 22318
rect 37550 22370 37602 22382
rect 37550 22306 37602 22318
rect 38222 22370 38274 22382
rect 38222 22306 38274 22318
rect 41470 22370 41522 22382
rect 44830 22370 44882 22382
rect 42242 22318 42254 22370
rect 42306 22318 42318 22370
rect 41470 22306 41522 22318
rect 44830 22306 44882 22318
rect 45694 22287 45706 22339
rect 45758 22287 45770 22339
rect 46722 22290 46734 22342
rect 46786 22290 46798 22342
rect 48962 22318 48974 22370
rect 49026 22318 49038 22370
rect 29978 22206 29990 22258
rect 30042 22206 30054 22258
rect 27638 22194 27690 22206
rect 34134 22194 34186 22206
rect 44158 22258 44210 22270
rect 44158 22194 44210 22206
rect 18230 22146 18282 22158
rect 18230 22082 18282 22094
rect 19630 22146 19682 22158
rect 19630 22082 19682 22094
rect 20526 22146 20578 22158
rect 20526 22082 20578 22094
rect 21758 22146 21810 22158
rect 21758 22082 21810 22094
rect 22486 22146 22538 22158
rect 22486 22082 22538 22094
rect 30550 22146 30602 22158
rect 30550 22082 30602 22094
rect 37886 22146 37938 22158
rect 37886 22082 37938 22094
rect 1344 21978 49616 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 49616 21978
rect 1344 21892 49616 21926
rect 9886 21810 9938 21822
rect 9886 21746 9938 21758
rect 11398 21810 11450 21822
rect 11398 21746 11450 21758
rect 37214 21810 37266 21822
rect 37214 21746 37266 21758
rect 38558 21810 38610 21822
rect 38558 21746 38610 21758
rect 39230 21810 39282 21822
rect 39230 21746 39282 21758
rect 43262 21810 43314 21822
rect 43262 21746 43314 21758
rect 44438 21810 44490 21822
rect 44438 21746 44490 21758
rect 6414 21698 6466 21710
rect 6414 21634 6466 21646
rect 15150 21698 15202 21710
rect 16550 21698 16602 21710
rect 15150 21634 15202 21646
rect 15635 21642 15687 21654
rect 1598 21586 1650 21598
rect 1598 21522 1650 21534
rect 5294 21586 5346 21598
rect 5294 21522 5346 21534
rect 5518 21586 5570 21598
rect 7534 21586 7586 21598
rect 6645 21534 6657 21586
rect 6709 21534 6721 21586
rect 5518 21522 5570 21534
rect 7534 21522 7586 21534
rect 10222 21586 10274 21598
rect 10222 21522 10274 21534
rect 10894 21586 10946 21598
rect 12462 21586 12514 21598
rect 15810 21590 15822 21642
rect 15874 21590 15886 21642
rect 16034 21590 16046 21642
rect 16098 21590 16110 21642
rect 16258 21590 16270 21642
rect 16322 21590 16334 21642
rect 16550 21634 16602 21646
rect 33406 21698 33458 21710
rect 46610 21702 46622 21754
rect 46674 21702 46686 21754
rect 12002 21534 12014 21586
rect 12066 21534 12078 21586
rect 13234 21534 13246 21586
rect 13298 21534 13310 21586
rect 15635 21578 15687 21590
rect 20638 21586 20690 21598
rect 23662 21586 23714 21598
rect 17266 21534 17278 21586
rect 17330 21534 17342 21586
rect 19842 21534 19854 21586
rect 19906 21534 19918 21586
rect 22866 21534 22878 21586
rect 22930 21534 22942 21586
rect 23986 21578 23998 21630
rect 24050 21578 24062 21630
rect 25678 21586 25730 21598
rect 24322 21534 24334 21586
rect 24386 21534 24398 21586
rect 10894 21522 10946 21534
rect 12462 21522 12514 21534
rect 20638 21522 20690 21534
rect 23662 21522 23714 21534
rect 25678 21522 25730 21534
rect 26574 21586 26626 21598
rect 26574 21522 26626 21534
rect 26966 21586 27018 21598
rect 26966 21522 27018 21534
rect 27806 21586 27858 21598
rect 31266 21590 31278 21642
rect 31330 21590 31342 21642
rect 33406 21634 33458 21646
rect 31614 21586 31666 21598
rect 30930 21534 30942 21586
rect 30994 21534 31006 21586
rect 27806 21522 27858 21534
rect 31614 21522 31666 21534
rect 36094 21586 36146 21598
rect 36094 21522 36146 21534
rect 36206 21586 36258 21598
rect 36206 21522 36258 21534
rect 37550 21586 37602 21598
rect 37550 21522 37602 21534
rect 38222 21586 38274 21598
rect 38222 21522 38274 21534
rect 38894 21586 38946 21598
rect 38894 21522 38946 21534
rect 39566 21586 39618 21598
rect 39566 21522 39618 21534
rect 39678 21586 39730 21598
rect 41122 21534 41134 21586
rect 41186 21534 41198 21586
rect 41906 21534 41918 21586
rect 41970 21534 41982 21586
rect 42354 21578 42366 21630
rect 42418 21578 42430 21630
rect 43598 21586 43650 21598
rect 42690 21534 42702 21586
rect 42754 21534 42766 21586
rect 39678 21522 39730 21534
rect 43598 21522 43650 21534
rect 44886 21586 44938 21598
rect 45266 21534 45278 21586
rect 45330 21534 45342 21586
rect 45490 21578 45502 21630
rect 45554 21578 45566 21630
rect 46398 21625 46450 21637
rect 46174 21586 46226 21598
rect 46398 21561 46450 21573
rect 46834 21534 46846 21586
rect 46898 21534 46910 21586
rect 47730 21549 47742 21601
rect 47794 21549 47806 21601
rect 48638 21586 48690 21598
rect 48066 21534 48078 21586
rect 48130 21534 48142 21586
rect 44886 21522 44938 21534
rect 46174 21522 46226 21534
rect 48638 21522 48690 21534
rect 48862 21586 48914 21598
rect 48862 21522 48914 21534
rect 11846 21474 11898 21486
rect 31278 21474 31330 21486
rect 2370 21422 2382 21474
rect 2434 21422 2446 21474
rect 4274 21422 4286 21474
rect 4338 21422 4350 21474
rect 17938 21422 17950 21474
rect 18002 21422 18014 21474
rect 20962 21422 20974 21474
rect 21026 21422 21038 21474
rect 23874 21422 23886 21474
rect 23938 21422 23950 21474
rect 28578 21422 28590 21474
rect 28642 21422 28654 21474
rect 30482 21422 30494 21474
rect 30546 21422 30558 21474
rect 11846 21410 11898 21422
rect 31278 21410 31330 21422
rect 32566 21474 32618 21486
rect 37886 21474 37938 21486
rect 43990 21474 44042 21486
rect 47350 21474 47402 21486
rect 35298 21422 35310 21474
rect 35362 21422 35374 21474
rect 32566 21410 32618 21422
rect 37886 21410 37938 21422
rect 41302 21418 41354 21430
rect 42242 21422 42254 21474
rect 42306 21422 42318 21474
rect 45602 21422 45614 21474
rect 45666 21422 45678 21474
rect 47618 21422 47630 21474
rect 47682 21422 47694 21474
rect 10558 21362 10610 21374
rect 5786 21310 5798 21362
rect 5850 21310 5862 21362
rect 10558 21298 10610 21310
rect 12182 21362 12234 21374
rect 12182 21298 12234 21310
rect 17446 21362 17498 21374
rect 17446 21298 17498 21310
rect 25342 21362 25394 21374
rect 25342 21298 25394 21310
rect 26238 21362 26290 21374
rect 26238 21298 26290 21310
rect 36542 21362 36594 21374
rect 36542 21298 36594 21310
rect 40014 21362 40066 21374
rect 43990 21410 44042 21422
rect 47350 21410 47402 21422
rect 41302 21354 41354 21366
rect 41750 21362 41802 21374
rect 40014 21298 40066 21310
rect 49130 21310 49142 21362
rect 49194 21310 49206 21362
rect 41750 21298 41802 21310
rect 1344 21194 49616 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 49616 21194
rect 1344 21108 49616 21142
rect 2046 21026 2098 21038
rect 2046 20962 2098 20974
rect 7086 21026 7138 21038
rect 7086 20962 7138 20974
rect 7702 21026 7754 21038
rect 7702 20962 7754 20974
rect 19518 21026 19570 21038
rect 14690 20918 14702 20970
rect 14754 20918 14766 20970
rect 19518 20962 19570 20974
rect 21366 21026 21418 21038
rect 21366 20962 21418 20974
rect 22766 21026 22818 21038
rect 22766 20962 22818 20974
rect 24110 21026 24162 21038
rect 24110 20962 24162 20974
rect 24782 21026 24834 21038
rect 24782 20962 24834 20974
rect 28366 21026 28418 21038
rect 34302 21026 34354 21038
rect 28366 20962 28418 20974
rect 32958 20970 33010 20982
rect 20358 20914 20410 20926
rect 30550 20914 30602 20926
rect 2594 20862 2606 20914
rect 2658 20862 2670 20914
rect 6470 20858 6522 20870
rect 10098 20862 10110 20914
rect 10162 20862 10174 20914
rect 25890 20862 25902 20914
rect 25954 20862 25966 20914
rect 27794 20862 27806 20914
rect 27858 20862 27870 20914
rect 34302 20962 34354 20974
rect 32958 20906 33010 20918
rect 43150 20914 43202 20926
rect 34738 20862 34750 20914
rect 34802 20862 34814 20914
rect 38770 20862 38782 20914
rect 38834 20862 38846 20914
rect 45042 20862 45054 20914
rect 45106 20862 45118 20914
rect 2382 20802 2434 20814
rect 4062 20802 4114 20814
rect 2382 20738 2434 20750
rect 2706 20735 2718 20787
rect 2770 20735 2782 20787
rect 3042 20750 3054 20802
rect 3106 20750 3118 20802
rect 3378 20750 3390 20802
rect 3442 20750 3454 20802
rect 3714 20723 3726 20775
rect 3778 20723 3790 20775
rect 4062 20738 4114 20750
rect 4958 20802 5010 20814
rect 4958 20738 5010 20750
rect 5182 20802 5234 20814
rect 5182 20738 5234 20750
rect 6190 20802 6242 20814
rect 20358 20850 20410 20862
rect 30550 20850 30602 20862
rect 43150 20850 43202 20862
rect 6470 20794 6522 20806
rect 6638 20802 6690 20814
rect 6190 20738 6242 20750
rect 6638 20738 6690 20750
rect 7422 20802 7474 20814
rect 9326 20802 9378 20814
rect 7858 20750 7870 20802
rect 7922 20750 7934 20802
rect 7422 20738 7474 20750
rect 9326 20738 9378 20750
rect 12350 20802 12402 20814
rect 12350 20738 12402 20750
rect 12574 20802 12626 20814
rect 12574 20738 12626 20750
rect 13358 20802 13410 20814
rect 17614 20802 17666 20814
rect 14578 20750 14590 20802
rect 14642 20750 14654 20802
rect 13358 20738 13410 20750
rect 15318 20712 15330 20764
rect 15382 20712 15394 20764
rect 15922 20722 15934 20774
rect 15986 20722 15998 20774
rect 17614 20738 17666 20750
rect 18398 20802 18450 20814
rect 22430 20802 22482 20814
rect 19262 20750 19274 20802
rect 19326 20750 19338 20802
rect 20850 20750 20862 20802
rect 20914 20750 20926 20802
rect 21590 20767 21642 20779
rect 18398 20738 18450 20750
rect 21590 20703 21642 20715
rect 21870 20774 21922 20786
rect 21870 20710 21922 20722
rect 22094 20774 22146 20786
rect 22094 20710 22146 20722
rect 22206 20746 22258 20758
rect 5910 20690 5962 20702
rect 4666 20638 4678 20690
rect 4730 20638 4742 20690
rect 3490 20582 3502 20634
rect 3554 20582 3566 20634
rect 5910 20626 5962 20638
rect 6302 20690 6354 20702
rect 6302 20626 6354 20638
rect 12014 20690 12066 20702
rect 22430 20738 22482 20750
rect 23102 20802 23154 20814
rect 23102 20738 23154 20750
rect 23774 20802 23826 20814
rect 23774 20738 23826 20750
rect 24446 20802 24498 20814
rect 24446 20738 24498 20750
rect 25118 20802 25170 20814
rect 25118 20738 25170 20750
rect 28702 20802 28754 20814
rect 28702 20738 28754 20750
rect 29206 20802 29258 20814
rect 33966 20802 34018 20814
rect 35422 20802 35474 20814
rect 29206 20738 29258 20750
rect 29486 20774 29538 20786
rect 29486 20710 29538 20722
rect 29710 20774 29762 20786
rect 29710 20710 29762 20722
rect 29934 20774 29986 20786
rect 29934 20710 29986 20722
rect 30046 20746 30098 20758
rect 33058 20750 33070 20802
rect 33122 20750 33134 20802
rect 12842 20638 12854 20690
rect 12906 20638 12918 20690
rect 22206 20682 22258 20694
rect 31378 20694 31390 20746
rect 31442 20694 31454 20746
rect 32050 20694 32062 20746
rect 32114 20694 32126 20746
rect 32386 20694 32398 20746
rect 32450 20694 32462 20746
rect 33734 20712 33746 20764
rect 33798 20712 33810 20764
rect 33966 20738 34018 20750
rect 34850 20735 34862 20787
rect 34914 20735 34926 20787
rect 35186 20750 35198 20802
rect 35250 20750 35262 20802
rect 35422 20738 35474 20750
rect 37438 20802 37490 20814
rect 37438 20738 37490 20750
rect 37998 20802 38050 20814
rect 44270 20802 44322 20814
rect 47742 20802 47794 20814
rect 48638 20802 48690 20814
rect 37998 20738 38050 20750
rect 41246 20763 41298 20775
rect 42366 20767 42418 20779
rect 30046 20682 30098 20694
rect 40686 20690 40738 20702
rect 41246 20699 41298 20711
rect 41750 20746 41802 20758
rect 12014 20626 12066 20638
rect 32622 20634 32674 20646
rect 20694 20578 20746 20590
rect 20694 20514 20746 20526
rect 23438 20578 23490 20590
rect 42018 20694 42030 20746
rect 42082 20694 42094 20746
rect 42242 20694 42254 20746
rect 42306 20694 42318 20746
rect 43381 20750 43393 20802
rect 43445 20750 43457 20802
rect 46946 20750 46958 20802
rect 47010 20750 47022 20802
rect 47954 20750 47966 20802
rect 48018 20750 48030 20802
rect 44270 20738 44322 20750
rect 47742 20738 47794 20750
rect 42366 20703 42418 20715
rect 48290 20694 48302 20746
rect 48354 20694 48366 20746
rect 48638 20738 48690 20750
rect 41750 20682 41802 20694
rect 40686 20626 40738 20638
rect 32622 20570 32674 20582
rect 35758 20578 35810 20590
rect 23438 20514 23490 20526
rect 35758 20514 35810 20526
rect 36374 20578 36426 20590
rect 36374 20514 36426 20526
rect 37102 20578 37154 20590
rect 37102 20514 37154 20526
rect 37830 20578 37882 20590
rect 48066 20582 48078 20634
rect 48130 20582 48142 20634
rect 37830 20514 37882 20526
rect 1344 20410 49616 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 49616 20410
rect 1344 20324 49616 20358
rect 8822 20242 8874 20254
rect 5282 20134 5294 20186
rect 5346 20134 5358 20186
rect 7186 20134 7198 20186
rect 7250 20134 7262 20186
rect 8822 20178 8874 20190
rect 23494 20242 23546 20254
rect 23494 20178 23546 20190
rect 46062 20242 46114 20254
rect 20246 20130 20298 20142
rect 12070 20074 12122 20086
rect 1598 20018 1650 20030
rect 4722 19966 4734 20018
rect 4786 19966 4798 20018
rect 5058 19993 5070 20045
rect 5122 19993 5134 20045
rect 5406 20018 5458 20030
rect 6638 20018 6690 20030
rect 6962 20022 6974 20074
rect 7026 20022 7038 20074
rect 7758 20056 7810 20068
rect 5842 19966 5854 20018
rect 5906 19966 5918 20018
rect 7298 19966 7310 20018
rect 7362 19966 7374 20018
rect 11510 20047 11562 20059
rect 8486 20018 8538 20030
rect 7758 19992 7810 20004
rect 8082 19966 8094 20018
rect 8146 19966 8158 20018
rect 8978 19966 8990 20018
rect 9042 19966 9054 20018
rect 12282 20022 12294 20074
rect 12346 20022 12358 20074
rect 12562 20022 12574 20074
rect 12626 20022 12638 20074
rect 20246 20066 20298 20078
rect 24054 20130 24106 20142
rect 29486 20130 29538 20142
rect 24054 20066 24106 20078
rect 28926 20074 28978 20086
rect 28366 20046 28418 20058
rect 11510 19983 11562 19995
rect 11778 19966 11790 20018
rect 11842 19966 11854 20018
rect 12070 20010 12122 20022
rect 13458 19993 13470 20045
rect 13522 19993 13534 20045
rect 16718 20018 16770 20030
rect 1598 19954 1650 19966
rect 5406 19954 5458 19966
rect 6638 19954 6690 19966
rect 8486 19954 8538 19966
rect 16718 19954 16770 19966
rect 16830 20018 16882 20030
rect 17378 19966 17390 20018
rect 17442 19966 17454 20018
rect 17714 19993 17726 20045
rect 17778 19993 17790 20045
rect 18062 20018 18114 20030
rect 19294 20018 19346 20030
rect 18722 19966 18734 20018
rect 18786 19966 18798 20018
rect 18946 19966 18958 20018
rect 19010 19966 19022 20018
rect 16830 19954 16882 19966
rect 18062 19954 18114 19966
rect 19294 19954 19346 19966
rect 21030 20018 21082 20030
rect 22542 20018 22594 20030
rect 21858 19966 21870 20018
rect 21922 19966 21934 20018
rect 22194 19966 22206 20018
rect 22258 19966 22270 20018
rect 21030 19954 21082 19966
rect 22542 19954 22594 19966
rect 24782 20018 24834 20030
rect 25218 19993 25230 20045
rect 25282 19993 25294 20045
rect 27458 19966 27470 20018
rect 27522 19966 27534 20018
rect 28366 19982 28418 19994
rect 28590 20046 28642 20058
rect 28802 20022 28814 20074
rect 28866 20022 28878 20074
rect 29486 20066 29538 20078
rect 33238 20130 33290 20142
rect 34358 20130 34410 20142
rect 40002 20134 40014 20186
rect 40066 20134 40078 20186
rect 46062 20178 46114 20190
rect 28926 20010 28978 20022
rect 29150 20018 29202 20030
rect 30146 20022 30158 20074
rect 30210 20022 30222 20074
rect 31278 20018 31330 20030
rect 31490 20022 31502 20074
rect 31554 20022 31566 20074
rect 33238 20066 33290 20078
rect 33518 20074 33570 20086
rect 33618 20022 33630 20074
rect 33682 20022 33694 20074
rect 34358 20066 34410 20078
rect 45334 20130 45386 20142
rect 33854 20046 33906 20058
rect 28590 19982 28642 19994
rect 30370 19966 30382 20018
rect 30434 19966 30446 20018
rect 24782 19954 24834 19966
rect 29150 19954 29202 19966
rect 30774 19962 30826 19974
rect 8318 19906 8370 19918
rect 21478 19906 21530 19918
rect 2370 19854 2382 19906
rect 2434 19854 2446 19906
rect 4274 19854 4286 19906
rect 4338 19854 4350 19906
rect 6022 19850 6074 19862
rect 11330 19854 11342 19906
rect 11394 19854 11406 19906
rect 17602 19854 17614 19906
rect 17666 19854 17678 19906
rect 8318 19842 8370 19854
rect 18622 19850 18674 19862
rect 6022 19786 6074 19798
rect 13022 19794 13074 19806
rect 13022 19730 13074 19742
rect 14478 19794 14530 19806
rect 21478 19842 21530 19854
rect 30606 19906 30658 19918
rect 31938 19966 31950 20018
rect 32002 19966 32014 20018
rect 33518 20010 33570 20022
rect 33854 19982 33906 19994
rect 34078 20046 34130 20058
rect 39902 20057 39954 20069
rect 34078 19982 34130 19994
rect 34638 20018 34690 20030
rect 31278 19954 31330 19966
rect 34638 19954 34690 19966
rect 34862 20018 34914 20030
rect 35130 19966 35142 20018
rect 35194 19966 35206 20018
rect 35970 19993 35982 20045
rect 36034 19993 36046 20045
rect 38546 19981 38558 20033
rect 38610 19981 38622 20033
rect 38882 19966 38894 20018
rect 38946 19966 38958 20018
rect 39554 19966 39566 20018
rect 39618 19966 39630 20018
rect 39902 19993 39954 20005
rect 40126 20018 40178 20030
rect 41178 20022 41190 20074
rect 41242 20022 41254 20074
rect 45334 20066 45386 20078
rect 41918 20018 41970 20030
rect 40898 19966 40910 20018
rect 40962 19966 40974 20018
rect 34862 19954 34914 19966
rect 40126 19954 40178 19966
rect 41918 19954 41970 19966
rect 42254 20018 42306 20030
rect 42910 20004 42922 20056
rect 42974 20004 42986 20056
rect 44046 20018 44098 20030
rect 44324 20018 44376 20030
rect 43586 19966 43598 20018
rect 43650 19966 43662 20018
rect 44146 19966 44158 20018
rect 44210 19966 44222 20018
rect 42254 19954 42306 19966
rect 44046 19954 44098 19966
rect 44324 19954 44376 19966
rect 46398 20018 46450 20030
rect 46722 20010 46734 20062
rect 46786 20010 46798 20062
rect 48638 20018 48690 20030
rect 47058 19966 47070 20018
rect 47122 19966 47134 20018
rect 47282 19966 47294 20018
rect 47346 19966 47358 20018
rect 46398 19954 46450 19966
rect 48638 19954 48690 19966
rect 48862 20018 48914 20030
rect 48862 19954 48914 19966
rect 30774 19898 30826 19910
rect 31614 19906 31666 19918
rect 16426 19742 16438 19794
rect 16490 19742 16502 19794
rect 18622 19786 18674 19798
rect 19630 19794 19682 19806
rect 21858 19798 21870 19850
rect 21922 19798 21934 19850
rect 30606 19842 30658 19854
rect 31614 19842 31666 19854
rect 32454 19906 32506 19918
rect 42646 19906 42698 19918
rect 38434 19854 38446 19906
rect 38498 19854 38510 19906
rect 41346 19854 41358 19906
rect 41410 19854 41422 19906
rect 32454 19842 32506 19854
rect 42646 19842 42698 19854
rect 43710 19850 43762 19862
rect 46610 19854 46622 19906
rect 46674 19854 46686 19906
rect 14478 19730 14530 19742
rect 19630 19730 19682 19742
rect 22878 19794 22930 19806
rect 22878 19730 22930 19742
rect 24446 19794 24498 19806
rect 24446 19730 24498 19742
rect 28086 19794 28138 19806
rect 28086 19730 28138 19742
rect 36990 19794 37042 19806
rect 43710 19786 43762 19798
rect 44718 19794 44770 19806
rect 36990 19730 37042 19742
rect 49130 19742 49142 19794
rect 49194 19742 49206 19794
rect 44718 19730 44770 19742
rect 1344 19626 49616 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 49616 19626
rect 1344 19540 49616 19574
rect 2046 19458 2098 19470
rect 2046 19394 2098 19406
rect 16998 19458 17050 19470
rect 16998 19394 17050 19406
rect 24558 19458 24610 19470
rect 24558 19394 24610 19406
rect 12966 19346 13018 19358
rect 4050 19294 4062 19346
rect 4114 19294 4126 19346
rect 5618 19294 5630 19346
rect 5682 19294 5694 19346
rect 9314 19294 9326 19346
rect 9378 19294 9390 19346
rect 10434 19294 10446 19346
rect 10498 19294 10510 19346
rect 12338 19294 12350 19346
rect 12402 19294 12414 19346
rect 12966 19282 13018 19294
rect 14590 19346 14642 19358
rect 17782 19346 17834 19358
rect 31042 19350 31054 19402
rect 31106 19350 31118 19402
rect 45446 19346 45498 19358
rect 14590 19282 14642 19294
rect 16438 19290 16490 19302
rect 2382 19234 2434 19246
rect 6638 19234 6690 19246
rect 9662 19234 9714 19246
rect 13918 19234 13970 19246
rect 14196 19234 14248 19246
rect 2382 19170 2434 19182
rect 4946 19154 4958 19206
rect 5010 19154 5022 19206
rect 5730 19138 5742 19190
rect 5794 19138 5806 19190
rect 5954 19182 5966 19234
rect 6018 19182 6030 19234
rect 7410 19182 7422 19234
rect 7474 19182 7486 19234
rect 13346 19182 13358 19234
rect 13410 19182 13422 19234
rect 14018 19182 14030 19234
rect 14082 19182 14094 19234
rect 6638 19170 6690 19182
rect 9662 19170 9714 19182
rect 13918 19170 13970 19182
rect 14196 19170 14248 19182
rect 15094 19234 15146 19246
rect 16270 19234 16322 19246
rect 15094 19170 15146 19182
rect 15318 19178 15370 19190
rect 15934 19178 15986 19190
rect 15586 19126 15598 19178
rect 15650 19126 15662 19178
rect 15810 19126 15822 19178
rect 15874 19126 15886 19178
rect 20066 19294 20078 19346
rect 20130 19294 20142 19346
rect 27570 19294 27582 19346
rect 27634 19294 27646 19346
rect 28466 19294 28478 19346
rect 28530 19294 28542 19346
rect 35746 19294 35758 19346
rect 35810 19294 35822 19346
rect 37874 19294 37886 19346
rect 37938 19294 37950 19346
rect 39778 19294 39790 19346
rect 39842 19294 39854 19346
rect 17782 19282 17834 19294
rect 45446 19282 45498 19294
rect 45894 19346 45946 19358
rect 49074 19294 49086 19346
rect 49138 19294 49150 19346
rect 45894 19282 45946 19294
rect 16438 19226 16490 19238
rect 16718 19234 16770 19246
rect 16270 19170 16322 19182
rect 16718 19170 16770 19182
rect 20862 19234 20914 19246
rect 20862 19170 20914 19182
rect 21198 19234 21250 19246
rect 24222 19234 24274 19246
rect 21970 19182 21982 19234
rect 22034 19182 22046 19234
rect 21198 19170 21250 19182
rect 24222 19170 24274 19182
rect 24894 19234 24946 19246
rect 36542 19234 36594 19246
rect 25666 19182 25678 19234
rect 25730 19182 25742 19234
rect 28130 19182 28142 19234
rect 28194 19182 28206 19234
rect 28310 19204 28362 19216
rect 24894 19170 24946 19182
rect 28310 19140 28362 19152
rect 29150 19199 29202 19211
rect 29150 19135 29202 19147
rect 29262 19206 29314 19218
rect 29262 19142 29314 19154
rect 29486 19206 29538 19218
rect 29486 19142 29538 19154
rect 29710 19206 29762 19218
rect 29710 19142 29762 19154
rect 30478 19144 30490 19196
rect 30542 19144 30554 19196
rect 31154 19182 31166 19234
rect 31218 19182 31230 19234
rect 15318 19114 15370 19126
rect 15934 19114 15986 19126
rect 16606 19122 16658 19134
rect 16606 19058 16658 19070
rect 18174 19122 18226 19134
rect 18174 19058 18226 19070
rect 23886 19122 23938 19134
rect 23886 19058 23938 19070
rect 29990 19122 30042 19134
rect 31714 19126 31726 19178
rect 31778 19126 31790 19178
rect 32162 19126 32174 19178
rect 32226 19126 32238 19178
rect 32834 19126 32846 19178
rect 32898 19126 32910 19178
rect 36542 19170 36594 19182
rect 37102 19234 37154 19246
rect 40574 19234 40626 19246
rect 40282 19182 40294 19234
rect 40346 19182 40358 19234
rect 37102 19170 37154 19182
rect 40574 19170 40626 19182
rect 40686 19234 40738 19246
rect 41470 19234 41522 19246
rect 46398 19234 46450 19246
rect 41010 19182 41022 19234
rect 41074 19182 41086 19234
rect 42242 19182 42254 19234
rect 42306 19182 42318 19234
rect 47170 19182 47182 19234
rect 47234 19182 47246 19234
rect 40686 19170 40738 19182
rect 41470 19170 41522 19182
rect 46398 19170 46450 19182
rect 29990 19058 30042 19070
rect 33854 19122 33906 19134
rect 13526 19010 13578 19022
rect 32722 19014 32734 19066
rect 32786 19014 32798 19066
rect 33854 19058 33906 19070
rect 44158 19122 44210 19134
rect 44158 19058 44210 19070
rect 13526 18946 13578 18958
rect 41190 19010 41242 19022
rect 41190 18946 41242 18958
rect 44998 19010 45050 19022
rect 44998 18946 45050 18958
rect 1344 18842 49616 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 49616 18842
rect 1344 18756 49616 18790
rect 8094 18674 8146 18686
rect 4274 18566 4286 18618
rect 4338 18566 4350 18618
rect 7410 18566 7422 18618
rect 7474 18566 7486 18618
rect 8094 18610 8146 18622
rect 19798 18674 19850 18686
rect 19798 18610 19850 18622
rect 24054 18674 24106 18686
rect 24054 18610 24106 18622
rect 26014 18674 26066 18686
rect 26014 18610 26066 18622
rect 27302 18674 27354 18686
rect 27302 18610 27354 18622
rect 43430 18674 43482 18686
rect 47070 18674 47122 18686
rect 43430 18610 43482 18622
rect 44046 18618 44098 18630
rect 11678 18562 11730 18574
rect 19238 18562 19290 18574
rect 17770 18510 17782 18562
rect 17834 18510 17846 18562
rect 3054 18450 3106 18462
rect 2034 18398 2046 18450
rect 2098 18398 2110 18450
rect 3490 18398 3502 18450
rect 3554 18398 3566 18450
rect 3714 18442 3726 18494
rect 3778 18442 3790 18494
rect 4398 18450 4450 18462
rect 4722 18454 4734 18506
rect 4786 18454 4798 18506
rect 7086 18489 7138 18501
rect 11678 18498 11730 18510
rect 18566 18506 18618 18518
rect 5742 18450 5794 18462
rect 4946 18398 4958 18450
rect 5010 18398 5022 18450
rect 3054 18386 3106 18398
rect 4398 18386 4450 18398
rect 5742 18386 5794 18398
rect 5854 18450 5906 18462
rect 6066 18398 6078 18450
rect 6130 18398 6142 18450
rect 6626 18398 6638 18450
rect 6690 18398 6702 18450
rect 18398 18485 18450 18497
rect 7086 18425 7138 18437
rect 7310 18450 7362 18462
rect 5854 18386 5906 18398
rect 7310 18386 7362 18398
rect 7758 18450 7810 18462
rect 12798 18450 12850 18462
rect 11909 18398 11921 18450
rect 11973 18398 11985 18450
rect 7758 18386 7810 18398
rect 12798 18386 12850 18398
rect 13358 18450 13410 18462
rect 13358 18386 13410 18398
rect 13470 18450 13522 18462
rect 14030 18450 14082 18462
rect 13738 18398 13750 18450
rect 13802 18398 13814 18450
rect 13470 18386 13522 18398
rect 14030 18386 14082 18398
rect 17278 18450 17330 18462
rect 17278 18386 17330 18398
rect 17502 18450 17554 18462
rect 18566 18442 18618 18454
rect 18790 18506 18842 18518
rect 47070 18610 47122 18622
rect 44046 18554 44098 18566
rect 19238 18498 19290 18510
rect 33070 18506 33122 18518
rect 18790 18442 18842 18454
rect 18958 18478 19010 18490
rect 18398 18421 18450 18433
rect 18958 18414 19010 18426
rect 20246 18450 20298 18462
rect 17502 18386 17554 18398
rect 20738 18398 20750 18450
rect 20802 18398 20814 18450
rect 21522 18398 21534 18450
rect 21586 18398 21598 18450
rect 22262 18436 22274 18488
rect 22326 18436 22338 18488
rect 22542 18450 22594 18462
rect 24222 18450 24274 18462
rect 23202 18398 23214 18450
rect 23266 18398 23278 18450
rect 20246 18386 20298 18398
rect 22542 18386 22594 18398
rect 24222 18386 24274 18398
rect 26350 18450 26402 18462
rect 26350 18386 26402 18398
rect 28030 18450 28082 18462
rect 28030 18386 28082 18398
rect 28142 18450 28194 18462
rect 28142 18386 28194 18398
rect 30830 18450 30882 18462
rect 31602 18398 31614 18450
rect 31666 18398 31678 18450
rect 31938 18425 31950 18477
rect 32002 18425 32014 18477
rect 32286 18450 32338 18462
rect 33462 18506 33514 18518
rect 33070 18442 33122 18454
rect 33238 18485 33290 18497
rect 33462 18442 33514 18454
rect 33630 18478 33682 18490
rect 33238 18421 33290 18433
rect 33630 18414 33682 18426
rect 33910 18450 33962 18462
rect 30830 18386 30882 18398
rect 32286 18386 32338 18398
rect 33910 18386 33962 18398
rect 34526 18450 34578 18462
rect 37214 18450 37266 18462
rect 36418 18398 36430 18450
rect 36482 18398 36494 18450
rect 37650 18398 37662 18450
rect 37714 18398 37726 18450
rect 39890 18425 39902 18477
rect 39954 18425 39966 18477
rect 41010 18398 41022 18450
rect 41074 18398 41086 18450
rect 41234 18413 41246 18465
rect 41298 18413 41310 18465
rect 41582 18450 41634 18462
rect 34526 18386 34578 18398
rect 37214 18386 37266 18398
rect 41582 18386 41634 18398
rect 41806 18450 41858 18462
rect 41806 18386 41858 18398
rect 42366 18450 42418 18462
rect 42366 18386 42418 18398
rect 42590 18450 42642 18462
rect 43810 18398 43822 18450
rect 43874 18398 43886 18450
rect 44034 18413 44046 18465
rect 44098 18413 44110 18465
rect 44494 18450 44546 18462
rect 45950 18450 46002 18462
rect 45358 18398 45370 18450
rect 45422 18398 45434 18450
rect 42590 18386 42642 18398
rect 44494 18386 44546 18398
rect 45950 18386 46002 18398
rect 46174 18450 46226 18462
rect 47406 18450 47458 18462
rect 46442 18398 46454 18450
rect 46506 18398 46518 18450
rect 46174 18386 46226 18398
rect 47406 18386 47458 18398
rect 47518 18450 47570 18462
rect 49086 18450 49138 18462
rect 48794 18398 48806 18450
rect 48858 18398 48870 18450
rect 47518 18386 47570 18398
rect 49086 18386 49138 18398
rect 49198 18450 49250 18462
rect 49198 18386 49250 18398
rect 24558 18338 24610 18350
rect 3826 18286 3838 18338
rect 3890 18286 3902 18338
rect 6246 18282 6298 18294
rect 14802 18286 14814 18338
rect 14866 18286 14878 18338
rect 16706 18286 16718 18338
rect 16770 18286 16782 18338
rect 2718 18226 2770 18238
rect 5450 18174 5462 18226
rect 5514 18174 5526 18226
rect 6246 18218 6298 18230
rect 20918 18282 20970 18294
rect 21746 18230 21758 18282
rect 21810 18230 21822 18282
rect 23314 18230 23326 18282
rect 23378 18230 23390 18282
rect 24558 18274 24610 18286
rect 27694 18338 27746 18350
rect 40406 18338 40458 18350
rect 28914 18286 28926 18338
rect 28978 18286 28990 18338
rect 31714 18286 31726 18338
rect 31778 18286 31790 18338
rect 41346 18286 41358 18338
rect 41410 18286 41422 18338
rect 27694 18274 27746 18286
rect 40406 18274 40458 18286
rect 20918 18218 20970 18230
rect 45614 18226 45666 18238
rect 42074 18174 42086 18226
rect 42138 18174 42150 18226
rect 42858 18174 42870 18226
rect 42922 18174 42934 18226
rect 2718 18162 2770 18174
rect 45614 18162 45666 18174
rect 47854 18226 47906 18238
rect 47854 18162 47906 18174
rect 1344 18058 49616 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 49616 18058
rect 1344 17972 49616 18006
rect 4846 17890 4898 17902
rect 4846 17826 4898 17838
rect 7646 17890 7698 17902
rect 42814 17890 42866 17902
rect 35018 17838 35030 17890
rect 35082 17838 35094 17890
rect 7646 17826 7698 17838
rect 42814 17826 42866 17838
rect 19350 17778 19402 17790
rect 2370 17726 2382 17778
rect 2434 17726 2446 17778
rect 7074 17726 7086 17778
rect 7138 17726 7150 17778
rect 8978 17726 8990 17778
rect 9042 17726 9054 17778
rect 11554 17726 11566 17778
rect 11618 17726 11630 17778
rect 15542 17722 15594 17734
rect 15810 17726 15822 17778
rect 15874 17726 15886 17778
rect 1598 17666 1650 17678
rect 1598 17602 1650 17614
rect 4286 17666 4338 17678
rect 4286 17602 4338 17614
rect 5182 17666 5234 17678
rect 5182 17602 5234 17614
rect 6190 17666 6242 17678
rect 6190 17602 6242 17614
rect 6302 17666 6354 17678
rect 7310 17666 7362 17678
rect 9942 17666 9994 17678
rect 12574 17666 12626 17678
rect 6626 17614 6638 17666
rect 6690 17614 6702 17666
rect 6302 17602 6354 17614
rect 6962 17570 6974 17622
rect 7026 17570 7038 17622
rect 7310 17602 7362 17614
rect 8306 17599 8318 17651
rect 8370 17599 8382 17651
rect 8642 17614 8654 17666
rect 8706 17614 8718 17666
rect 9090 17570 9102 17622
rect 9154 17570 9166 17622
rect 9314 17614 9326 17666
rect 9378 17614 9390 17666
rect 11218 17614 11230 17666
rect 11282 17614 11294 17666
rect 9942 17602 9994 17614
rect 11442 17599 11454 17651
rect 11506 17599 11518 17651
rect 11890 17614 11902 17666
rect 11954 17614 11966 17666
rect 12226 17587 12238 17639
rect 12290 17587 12302 17639
rect 12574 17602 12626 17614
rect 13358 17666 13410 17678
rect 13358 17602 13410 17614
rect 13582 17666 13634 17678
rect 19350 17714 19402 17726
rect 26238 17778 26290 17790
rect 45490 17782 45502 17834
rect 45554 17782 45566 17834
rect 41010 17726 41022 17778
rect 41074 17726 41086 17778
rect 43922 17726 43934 17778
rect 43986 17726 43998 17778
rect 48514 17726 48526 17778
rect 48578 17726 48590 17778
rect 26238 17714 26290 17726
rect 13850 17614 13862 17666
rect 13914 17614 13926 17666
rect 13582 17602 13634 17614
rect 14814 17610 14866 17622
rect 15138 17614 15150 17666
rect 15202 17614 15214 17666
rect 15542 17658 15594 17670
rect 16494 17666 16546 17678
rect 15922 17570 15934 17622
rect 15986 17570 15998 17622
rect 16146 17614 16158 17666
rect 16210 17614 16222 17666
rect 16494 17602 16546 17614
rect 16718 17666 16770 17678
rect 16718 17602 16770 17614
rect 17950 17666 18002 17678
rect 17950 17602 18002 17614
rect 18398 17666 18450 17678
rect 23102 17666 23154 17678
rect 18398 17602 18450 17614
rect 21310 17610 21362 17622
rect 5898 17502 5910 17554
rect 5962 17502 5974 17554
rect 14814 17546 14866 17558
rect 15374 17554 15426 17566
rect 16986 17502 16998 17554
rect 17050 17502 17062 17554
rect 21310 17546 21362 17558
rect 21422 17610 21474 17622
rect 22150 17610 22202 17622
rect 21422 17546 21474 17558
rect 21982 17554 22034 17566
rect 23102 17602 23154 17614
rect 23326 17666 23378 17678
rect 23326 17602 23378 17614
rect 23774 17666 23826 17678
rect 25846 17666 25898 17678
rect 26910 17666 26962 17678
rect 24770 17614 24782 17666
rect 24834 17614 24846 17666
rect 23482 17558 23494 17610
rect 23546 17558 23558 17610
rect 23774 17602 23826 17614
rect 25218 17586 25230 17638
rect 25282 17586 25294 17638
rect 25442 17614 25454 17666
rect 25506 17614 25518 17666
rect 26786 17614 26798 17666
rect 26850 17614 26862 17666
rect 25846 17602 25898 17614
rect 22150 17546 22202 17558
rect 23662 17554 23714 17566
rect 8418 17446 8430 17498
rect 8482 17446 8494 17498
rect 12002 17446 12014 17498
rect 12066 17446 12078 17498
rect 15374 17490 15426 17502
rect 21982 17490 22034 17502
rect 23662 17490 23714 17502
rect 24054 17554 24106 17566
rect 24054 17490 24106 17502
rect 25678 17554 25730 17566
rect 26620 17558 26632 17610
rect 26684 17558 26696 17610
rect 26910 17602 26962 17614
rect 27694 17666 27746 17678
rect 27694 17602 27746 17614
rect 28086 17666 28138 17678
rect 31950 17666 32002 17678
rect 31154 17614 31166 17666
rect 31218 17614 31230 17666
rect 35310 17666 35362 17678
rect 28086 17602 28138 17614
rect 31950 17602 32002 17614
rect 32162 17586 32174 17638
rect 32226 17586 32238 17638
rect 35310 17602 35362 17614
rect 35422 17666 35474 17678
rect 35422 17602 35474 17614
rect 35646 17666 35698 17678
rect 38222 17666 38274 17678
rect 36866 17614 36878 17666
rect 36930 17614 36942 17666
rect 35646 17602 35698 17614
rect 38222 17602 38274 17614
rect 38334 17666 38386 17678
rect 42142 17666 42194 17678
rect 39106 17614 39118 17666
rect 39170 17614 39182 17666
rect 41458 17614 41470 17666
rect 41522 17614 41534 17666
rect 38334 17602 38386 17614
rect 25678 17490 25730 17502
rect 29262 17554 29314 17566
rect 41738 17558 41750 17610
rect 41802 17558 41814 17610
rect 42142 17602 42194 17614
rect 43150 17666 43202 17678
rect 46622 17666 46674 17678
rect 43474 17614 43486 17666
rect 43538 17614 43550 17666
rect 43150 17602 43202 17614
rect 43810 17599 43822 17651
rect 43874 17599 43886 17651
rect 45266 17614 45278 17666
rect 45330 17614 45342 17666
rect 45490 17614 45502 17666
rect 45554 17614 45566 17666
rect 46622 17602 46674 17614
rect 49310 17666 49362 17678
rect 49310 17602 49362 17614
rect 29262 17490 29314 17502
rect 17614 17442 17666 17454
rect 17614 17378 17666 17390
rect 18734 17442 18786 17454
rect 18734 17378 18786 17390
rect 22766 17442 22818 17454
rect 22766 17378 22818 17390
rect 24614 17442 24666 17454
rect 24614 17378 24666 17390
rect 27358 17442 27410 17454
rect 27358 17378 27410 17390
rect 35982 17442 36034 17454
rect 35982 17378 36034 17390
rect 37886 17442 37938 17454
rect 41570 17446 41582 17498
rect 41634 17446 41646 17498
rect 37886 17378 37938 17390
rect 46118 17442 46170 17454
rect 46118 17378 46170 17390
rect 1344 17274 49616 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 49616 17274
rect 1344 17188 49616 17222
rect 6134 17106 6186 17118
rect 4286 16994 4338 17006
rect 5282 16998 5294 17050
rect 5346 16998 5358 17050
rect 6134 17042 6186 17054
rect 28590 17106 28642 17118
rect 28590 17042 28642 17054
rect 36710 17106 36762 17118
rect 36710 17042 36762 17054
rect 37158 17106 37210 17118
rect 37158 17042 37210 17054
rect 37886 17106 37938 17118
rect 37886 17042 37938 17054
rect 40126 17106 40178 17118
rect 40126 17042 40178 17054
rect 48974 17106 49026 17118
rect 48974 17042 49026 17054
rect 12798 16994 12850 17006
rect 8698 16942 8710 16994
rect 8762 16942 8774 16994
rect 4286 16930 4338 16942
rect 1598 16882 1650 16894
rect 4834 16830 4846 16882
rect 4898 16830 4910 16882
rect 5058 16857 5070 16909
rect 5122 16857 5134 16909
rect 5406 16882 5458 16894
rect 6850 16886 6862 16938
rect 6914 16886 6926 16938
rect 12798 16930 12850 16942
rect 13358 16994 13410 17006
rect 13358 16930 13410 16942
rect 23438 16994 23490 17006
rect 33238 16994 33290 17006
rect 7086 16882 7138 16894
rect 6402 16830 6414 16882
rect 6466 16830 6478 16882
rect 1598 16818 1650 16830
rect 5406 16818 5458 16830
rect 7086 16818 7138 16830
rect 7422 16882 7474 16894
rect 7422 16818 7474 16830
rect 8206 16882 8258 16894
rect 8206 16818 8258 16830
rect 8430 16882 8482 16894
rect 8430 16818 8482 16830
rect 9438 16882 9490 16894
rect 9438 16818 9490 16830
rect 10110 16882 10162 16894
rect 10110 16818 10162 16830
rect 16046 16882 16098 16894
rect 16370 16874 16382 16926
rect 16434 16874 16446 16926
rect 17838 16920 17890 16932
rect 16594 16830 16606 16882
rect 16658 16830 16670 16882
rect 19104 16920 19156 16932
rect 23438 16930 23490 16942
rect 24726 16938 24778 16950
rect 18846 16882 18898 16894
rect 17838 16856 17890 16868
rect 18162 16830 18174 16882
rect 18226 16830 18238 16882
rect 16046 16818 16098 16830
rect 18566 16826 18618 16838
rect 6750 16770 6802 16782
rect 18398 16770 18450 16782
rect 2370 16718 2382 16770
rect 2434 16718 2446 16770
rect 10882 16718 10894 16770
rect 10946 16718 10958 16770
rect 15250 16718 15262 16770
rect 15314 16718 15326 16770
rect 16258 16718 16270 16770
rect 16322 16718 16334 16770
rect 18946 16830 18958 16882
rect 19010 16830 19022 16882
rect 19104 16856 19156 16868
rect 20078 16882 20130 16894
rect 18846 16818 18898 16830
rect 20078 16818 20130 16830
rect 22766 16882 22818 16894
rect 22766 16818 22818 16830
rect 23102 16882 23154 16894
rect 24098 16886 24110 16938
rect 24162 16886 24174 16938
rect 26338 16886 26350 16938
rect 26402 16886 26414 16938
rect 27544 16920 27596 16932
rect 33238 16930 33290 16942
rect 41078 16994 41130 17006
rect 46330 16942 46342 16994
rect 46394 16942 46406 16994
rect 41078 16930 41130 16942
rect 24322 16830 24334 16882
rect 24386 16830 24398 16882
rect 24726 16874 24778 16886
rect 26798 16882 26850 16894
rect 26562 16830 26574 16882
rect 26626 16830 26638 16882
rect 23102 16818 23154 16830
rect 26798 16818 26850 16830
rect 26966 16882 27018 16894
rect 26966 16818 27018 16830
rect 27246 16882 27298 16894
rect 27346 16830 27358 16882
rect 27410 16830 27422 16882
rect 46902 16911 46954 16923
rect 27544 16856 27596 16868
rect 28926 16882 28978 16894
rect 27246 16818 27298 16830
rect 28926 16818 28978 16830
rect 29598 16882 29650 16894
rect 30370 16857 30382 16909
rect 30434 16857 30446 16909
rect 33406 16882 33458 16894
rect 29598 16818 29650 16830
rect 33406 16818 33458 16830
rect 37550 16882 37602 16894
rect 38546 16845 38558 16897
rect 38610 16845 38622 16897
rect 39230 16882 39282 16894
rect 38882 16830 38894 16882
rect 38946 16830 38958 16882
rect 37550 16818 37602 16830
rect 39230 16818 39282 16830
rect 39342 16882 39394 16894
rect 39342 16818 39394 16830
rect 40462 16882 40514 16894
rect 40462 16818 40514 16830
rect 42366 16882 42418 16894
rect 42366 16818 42418 16830
rect 42478 16882 42530 16894
rect 42478 16818 42530 16830
rect 42702 16882 42754 16894
rect 42702 16818 42754 16830
rect 42926 16882 42978 16894
rect 42926 16818 42978 16830
rect 44046 16882 44098 16894
rect 44046 16818 44098 16830
rect 44270 16882 44322 16894
rect 45166 16882 45218 16894
rect 44538 16830 44550 16882
rect 44602 16830 44614 16882
rect 44270 16818 44322 16830
rect 45166 16818 45218 16830
rect 45278 16882 45330 16894
rect 45950 16882 46002 16894
rect 45546 16830 45558 16882
rect 45610 16830 45622 16882
rect 49310 16882 49362 16894
rect 46902 16847 46954 16859
rect 45278 16818 45330 16830
rect 45950 16818 46002 16830
rect 46062 16826 46114 16838
rect 47058 16830 47070 16882
rect 47122 16830 47134 16882
rect 18566 16762 18618 16774
rect 19518 16770 19570 16782
rect 24558 16770 24610 16782
rect 6750 16706 6802 16718
rect 18398 16706 18450 16718
rect 20850 16718 20862 16770
rect 20914 16718 20926 16770
rect 19518 16706 19570 16718
rect 24558 16706 24610 16718
rect 27918 16770 27970 16782
rect 41750 16770 41802 16782
rect 34178 16718 34190 16770
rect 34242 16718 34254 16770
rect 36082 16718 36094 16770
rect 36146 16718 36158 16770
rect 38434 16718 38446 16770
rect 38498 16718 38510 16770
rect 49310 16818 49362 16830
rect 46062 16762 46114 16774
rect 46722 16718 46734 16770
rect 46786 16718 46798 16770
rect 27918 16706 27970 16718
rect 41750 16706 41802 16718
rect 9774 16658 9826 16670
rect 9774 16594 9826 16606
rect 29262 16658 29314 16670
rect 29262 16594 29314 16606
rect 31054 16658 31106 16670
rect 39610 16606 39622 16658
rect 39674 16606 39686 16658
rect 42074 16606 42086 16658
rect 42138 16606 42150 16658
rect 43194 16606 43206 16658
rect 43258 16606 43270 16658
rect 31054 16594 31106 16606
rect 1344 16490 49616 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 49616 16490
rect 1344 16404 49616 16438
rect 2494 16322 2546 16334
rect 11678 16322 11730 16334
rect 5002 16270 5014 16322
rect 5066 16270 5078 16322
rect 6122 16270 6134 16322
rect 6186 16270 6198 16322
rect 2494 16258 2546 16270
rect 11678 16258 11730 16270
rect 15038 16322 15090 16334
rect 15038 16258 15090 16270
rect 16662 16322 16714 16334
rect 20694 16322 20746 16334
rect 16662 16258 16714 16270
rect 20134 16266 20186 16278
rect 20694 16258 20746 16270
rect 21534 16322 21586 16334
rect 25510 16322 25562 16334
rect 21534 16258 21586 16270
rect 23326 16266 23378 16278
rect 3490 16158 3502 16210
rect 3554 16158 3566 16210
rect 4274 16158 4286 16210
rect 4338 16158 4350 16210
rect 6694 16154 6746 16166
rect 8530 16158 8542 16210
rect 8594 16158 8606 16210
rect 10434 16158 10446 16210
rect 10498 16158 10510 16210
rect 19058 16158 19070 16210
rect 19122 16158 19134 16210
rect 20134 16202 20186 16214
rect 25510 16258 25562 16270
rect 30146 16214 30158 16266
rect 30210 16214 30222 16266
rect 23326 16202 23378 16214
rect 36486 16210 36538 16222
rect 44214 16210 44266 16222
rect 49254 16210 49306 16222
rect 27906 16158 27918 16210
rect 27970 16158 27982 16210
rect 29586 16158 29598 16210
rect 29650 16158 29662 16210
rect 39554 16158 39566 16210
rect 39618 16158 39630 16210
rect 41122 16158 41134 16210
rect 41186 16158 41198 16210
rect 44930 16158 44942 16210
rect 44994 16158 45006 16210
rect 46834 16158 46846 16210
rect 46898 16158 46910 16210
rect 2830 16098 2882 16110
rect 4622 16098 4674 16110
rect 3154 16046 3166 16098
rect 3218 16046 3230 16098
rect 2830 16034 2882 16046
rect 3378 16031 3390 16083
rect 3442 16031 3454 16083
rect 3938 16046 3950 16098
rect 4002 16046 4014 16098
rect 4118 16068 4170 16080
rect 4622 16034 4674 16046
rect 4734 16098 4786 16110
rect 4734 16034 4786 16046
rect 5742 16098 5794 16110
rect 5742 16034 5794 16046
rect 5854 16098 5906 16110
rect 5854 16034 5906 16046
rect 6526 16098 6578 16110
rect 36486 16146 36538 16158
rect 44214 16146 44266 16158
rect 49254 16146 49306 16158
rect 6694 16090 6746 16102
rect 6974 16098 7026 16110
rect 6526 16034 6578 16046
rect 6974 16034 7026 16046
rect 11230 16098 11282 16110
rect 11230 16034 11282 16046
rect 12014 16098 12066 16110
rect 12014 16034 12066 16046
rect 13918 16098 13970 16110
rect 17166 16098 17218 16110
rect 14782 16046 14794 16098
rect 14846 16046 14858 16098
rect 16482 16046 16494 16098
rect 16546 16046 16558 16098
rect 13918 16034 13970 16046
rect 17166 16034 17218 16046
rect 19854 16098 19906 16110
rect 22206 16098 22258 16110
rect 23550 16098 23602 16110
rect 19854 16034 19906 16046
rect 19966 16077 20018 16089
rect 4118 16004 4170 16016
rect 20850 16046 20862 16098
rect 20914 16046 20926 16098
rect 22082 16046 22094 16098
rect 22146 16046 22158 16098
rect 22978 16046 22990 16098
rect 23042 16046 23054 16098
rect 23202 16046 23214 16098
rect 23266 16046 23278 16098
rect 19966 16013 20018 16025
rect 6862 15986 6914 15998
rect 6862 15922 6914 15934
rect 7254 15986 7306 15998
rect 21916 15990 21928 16042
rect 21980 15990 21992 16042
rect 22206 16034 22258 16046
rect 23550 16034 23602 16046
rect 24222 16098 24274 16110
rect 24222 16034 24274 16046
rect 24446 16098 24498 16110
rect 28702 16098 28754 16110
rect 30942 16098 30994 16110
rect 34526 16098 34578 16110
rect 35758 16098 35810 16110
rect 25330 16046 25342 16098
rect 25394 16046 25406 16098
rect 29250 16046 29262 16098
rect 29314 16046 29326 16098
rect 24446 16034 24498 16046
rect 28702 16034 28754 16046
rect 29474 16002 29486 16054
rect 29538 16002 29550 16054
rect 30034 16046 30046 16098
rect 30098 16046 30110 16098
rect 30774 16008 30786 16060
rect 30838 16008 30850 16060
rect 31714 16046 31726 16098
rect 31778 16046 31790 16098
rect 35074 16046 35086 16098
rect 35138 16046 35150 16098
rect 30942 16034 30994 16046
rect 34526 16034 34578 16046
rect 26014 15986 26066 15998
rect 24714 15934 24726 15986
rect 24778 15934 24790 15986
rect 7254 15922 7306 15934
rect 26014 15922 26066 15934
rect 33630 15986 33682 15998
rect 35522 15990 35534 16042
rect 35586 15990 35598 16042
rect 35758 16034 35810 16046
rect 36878 16098 36930 16110
rect 39902 16098 39954 16110
rect 37650 16046 37662 16098
rect 37714 16046 37726 16098
rect 36878 16034 36930 16046
rect 39902 16034 39954 16046
rect 40238 16098 40290 16110
rect 43822 16098 43874 16110
rect 43026 16046 43038 16098
rect 43090 16046 43102 16098
rect 40238 16034 40290 16046
rect 43822 16034 43874 16046
rect 47630 16098 47682 16110
rect 47630 16034 47682 16046
rect 47742 16098 47794 16110
rect 47742 16034 47794 16046
rect 33630 15922 33682 15934
rect 13638 15874 13690 15886
rect 13638 15810 13690 15822
rect 23886 15874 23938 15886
rect 23886 15810 23938 15822
rect 34190 15874 34242 15886
rect 35634 15878 35646 15930
rect 35698 15878 35710 15930
rect 34190 15810 34242 15822
rect 48078 15874 48130 15886
rect 48078 15810 48130 15822
rect 1344 15706 49616 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 49616 15706
rect 1344 15620 49616 15654
rect 9718 15538 9770 15550
rect 4610 15430 4622 15482
rect 4674 15430 4686 15482
rect 9718 15474 9770 15486
rect 20022 15538 20074 15550
rect 20022 15474 20074 15486
rect 24502 15538 24554 15550
rect 16494 15426 16546 15438
rect 23762 15430 23774 15482
rect 23826 15430 23838 15482
rect 24502 15474 24554 15486
rect 26406 15538 26458 15550
rect 37494 15538 37546 15550
rect 26406 15474 26458 15486
rect 31390 15482 31442 15494
rect 30494 15426 30546 15438
rect 2830 15314 2882 15326
rect 4778 15318 4790 15370
rect 4842 15318 4854 15370
rect 16494 15362 16546 15374
rect 18230 15370 18282 15382
rect 5182 15314 5234 15326
rect 4498 15262 4510 15314
rect 4562 15262 4574 15314
rect 5954 15262 5966 15314
rect 6018 15262 6030 15314
rect 6290 15306 6302 15358
rect 6354 15306 6366 15358
rect 9886 15334 9938 15346
rect 6974 15314 7026 15326
rect 2830 15250 2882 15262
rect 5182 15250 5234 15262
rect 6974 15250 7026 15262
rect 7198 15314 7250 15326
rect 7198 15250 7250 15262
rect 8038 15314 8090 15326
rect 9886 15270 9938 15282
rect 9986 15262 9998 15314
rect 10050 15262 10062 15314
rect 10994 15289 11006 15341
rect 11058 15289 11070 15341
rect 12238 15314 12290 15326
rect 8038 15250 8090 15262
rect 12238 15250 12290 15262
rect 13806 15314 13858 15326
rect 17602 15318 17614 15370
rect 17666 15318 17678 15370
rect 37494 15474 37546 15486
rect 44718 15538 44770 15550
rect 39106 15430 39118 15482
rect 39170 15430 39182 15482
rect 44718 15474 44770 15486
rect 31390 15418 31442 15430
rect 33114 15374 33126 15426
rect 33178 15374 33190 15426
rect 36810 15374 36822 15426
rect 36874 15374 36886 15426
rect 17826 15262 17838 15314
rect 17890 15262 17902 15314
rect 18230 15306 18282 15318
rect 19220 15352 19272 15364
rect 23662 15353 23714 15365
rect 30494 15362 30546 15374
rect 19518 15314 19570 15326
rect 19220 15288 19272 15300
rect 19394 15262 19406 15314
rect 19458 15262 19470 15314
rect 20290 15289 20302 15341
rect 20354 15289 20366 15341
rect 22530 15262 22542 15314
rect 22594 15262 22606 15314
rect 23202 15262 23214 15314
rect 23266 15262 23278 15314
rect 31502 15353 31554 15365
rect 23662 15289 23714 15301
rect 23886 15314 23938 15326
rect 25118 15314 25170 15326
rect 27806 15314 27858 15326
rect 24322 15262 24334 15314
rect 24386 15262 24398 15314
rect 26226 15262 26238 15314
rect 26290 15262 26302 15314
rect 28578 15262 28590 15314
rect 28642 15262 28654 15314
rect 31042 15262 31054 15314
rect 31106 15262 31118 15314
rect 31502 15289 31554 15301
rect 31726 15314 31778 15326
rect 13806 15250 13858 15262
rect 19518 15250 19570 15262
rect 23886 15250 23938 15262
rect 25118 15250 25170 15262
rect 27806 15250 27858 15262
rect 31726 15250 31778 15262
rect 33406 15314 33458 15326
rect 33406 15250 33458 15262
rect 33630 15314 33682 15326
rect 33630 15250 33682 15262
rect 33966 15314 34018 15326
rect 33966 15250 34018 15262
rect 34190 15314 34242 15326
rect 35198 15314 35250 15326
rect 34906 15262 34918 15314
rect 34970 15262 34982 15314
rect 34190 15250 34242 15262
rect 35198 15250 35250 15262
rect 35422 15314 35474 15326
rect 35746 15277 35758 15329
rect 35810 15277 35822 15329
rect 36318 15314 36370 15326
rect 36082 15262 36094 15314
rect 36146 15262 36158 15314
rect 35422 15250 35474 15262
rect 36318 15250 36370 15262
rect 36542 15314 36594 15326
rect 38770 15318 38782 15370
rect 38834 15318 38846 15370
rect 39006 15314 39058 15326
rect 38322 15262 38334 15314
rect 38386 15262 38398 15314
rect 36542 15250 36594 15262
rect 39006 15250 39058 15262
rect 39566 15314 39618 15326
rect 39566 15250 39618 15262
rect 39678 15314 39730 15326
rect 41906 15262 41918 15314
rect 41970 15262 41982 15314
rect 42242 15277 42254 15329
rect 42306 15277 42318 15329
rect 42802 15262 42814 15314
rect 42866 15262 42878 15314
rect 43026 15262 43038 15314
rect 43090 15262 43102 15314
rect 45714 15289 45726 15341
rect 45778 15289 45790 15341
rect 47350 15314 47402 15326
rect 46386 15262 46398 15314
rect 46450 15262 46462 15314
rect 46722 15262 46734 15314
rect 46786 15262 46798 15314
rect 47730 15277 47742 15329
rect 47794 15277 47806 15329
rect 48638 15314 48690 15326
rect 48066 15262 48078 15314
rect 48130 15262 48142 15314
rect 39678 15250 39730 15262
rect 47350 15250 47402 15262
rect 48638 15250 48690 15262
rect 18062 15202 18114 15214
rect 6402 15150 6414 15202
rect 6466 15150 6478 15202
rect 14578 15150 14590 15202
rect 14642 15150 14654 15202
rect 18062 15138 18114 15150
rect 18846 15202 18898 15214
rect 41638 15202 41690 15214
rect 35634 15150 35646 15202
rect 35698 15150 35710 15202
rect 42354 15150 42366 15202
rect 42418 15150 42430 15202
rect 18846 15138 18898 15150
rect 41638 15138 41690 15150
rect 42702 15146 42754 15158
rect 2494 15090 2546 15102
rect 25454 15090 25506 15102
rect 7466 15038 7478 15090
rect 7530 15038 7542 15090
rect 34458 15038 34470 15090
rect 34522 15038 34534 15090
rect 39946 15038 39958 15090
rect 40010 15038 40022 15090
rect 42702 15082 42754 15094
rect 46846 15146 46898 15158
rect 47618 15150 47630 15202
rect 47682 15150 47694 15202
rect 46846 15082 46898 15094
rect 48974 15090 49026 15102
rect 2494 15026 2546 15038
rect 25454 15026 25506 15038
rect 48974 15026 49026 15038
rect 1344 14922 49616 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 49616 14922
rect 1344 14836 49616 14870
rect 32622 14754 32674 14766
rect 30874 14702 30886 14754
rect 30938 14702 30950 14754
rect 42746 14702 42758 14754
rect 42810 14702 42822 14754
rect 32622 14690 32674 14702
rect 7422 14642 7474 14654
rect 20078 14642 20130 14654
rect 2370 14590 2382 14642
rect 2434 14590 2446 14642
rect 4274 14590 4286 14642
rect 4338 14590 4350 14642
rect 6402 14590 6414 14642
rect 6466 14590 6478 14642
rect 7422 14578 7474 14590
rect 7590 14586 7642 14598
rect 8530 14590 8542 14642
rect 8594 14590 8606 14642
rect 10434 14590 10446 14642
rect 10498 14590 10510 14642
rect 24882 14590 24894 14642
rect 24946 14590 24958 14642
rect 26786 14590 26798 14642
rect 26850 14590 26862 14642
rect 31602 14590 31614 14642
rect 31666 14590 31678 14642
rect 34178 14590 34190 14642
rect 34242 14590 34254 14642
rect 36978 14590 36990 14642
rect 37042 14590 37054 14642
rect 39778 14590 39790 14642
rect 39842 14590 39854 14642
rect 47170 14590 47182 14642
rect 47234 14590 47246 14642
rect 49074 14590 49086 14642
rect 49138 14590 49150 14642
rect 1598 14530 1650 14542
rect 1598 14466 1650 14478
rect 5182 14530 5234 14542
rect 20078 14578 20130 14590
rect 5954 14478 5966 14530
rect 6018 14478 6030 14530
rect 5182 14466 5234 14478
rect 6290 14463 6302 14515
rect 6354 14463 6366 14515
rect 6962 14450 6974 14502
rect 7026 14450 7038 14502
rect 7186 14478 7198 14530
rect 7250 14478 7262 14530
rect 7590 14522 7642 14534
rect 7758 14530 7810 14542
rect 7758 14466 7810 14478
rect 11790 14530 11842 14542
rect 13470 14530 13522 14542
rect 17278 14530 17330 14542
rect 11790 14466 11842 14478
rect 12114 14463 12126 14515
rect 12178 14463 12190 14515
rect 12450 14478 12462 14530
rect 12514 14478 12526 14530
rect 14242 14478 14254 14530
rect 14306 14478 14318 14530
rect 16594 14478 16606 14530
rect 16658 14478 16670 14530
rect 13470 14466 13522 14478
rect 16158 14418 16210 14430
rect 16930 14422 16942 14474
rect 16994 14422 17006 14474
rect 17278 14466 17330 14478
rect 18398 14530 18450 14542
rect 18398 14466 18450 14478
rect 18622 14530 18674 14542
rect 19686 14530 19738 14542
rect 18622 14466 18674 14478
rect 19058 14450 19070 14502
rect 19122 14450 19134 14502
rect 19282 14478 19294 14530
rect 19346 14478 19358 14530
rect 19686 14466 19738 14478
rect 20472 14530 20524 14542
rect 20750 14530 20802 14542
rect 20626 14478 20638 14530
rect 20690 14478 20702 14530
rect 27582 14530 27634 14542
rect 29934 14530 29986 14542
rect 20472 14466 20524 14478
rect 20750 14466 20802 14478
rect 21634 14450 21646 14502
rect 21698 14450 21710 14502
rect 29362 14478 29374 14530
rect 29426 14478 29438 14530
rect 29710 14491 29762 14503
rect 27582 14466 27634 14478
rect 29934 14466 29986 14478
rect 30494 14530 30546 14542
rect 30494 14466 30546 14478
rect 30606 14530 30658 14542
rect 32286 14530 32338 14542
rect 35870 14530 35922 14542
rect 37662 14530 37714 14542
rect 30606 14466 30658 14478
rect 31714 14463 31726 14515
rect 31778 14463 31790 14515
rect 31938 14478 31950 14530
rect 32002 14478 32014 14530
rect 33842 14478 33854 14530
rect 33906 14478 33918 14530
rect 32286 14466 32338 14478
rect 34066 14463 34078 14515
rect 34130 14463 34142 14515
rect 35186 14478 35198 14530
rect 35250 14478 35262 14530
rect 35646 14491 35698 14503
rect 19518 14418 19570 14430
rect 29710 14427 29762 14439
rect 35870 14466 35922 14478
rect 37090 14463 37102 14515
rect 37154 14463 37166 14515
rect 37314 14478 37326 14530
rect 37378 14478 37390 14530
rect 37662 14466 37714 14478
rect 38670 14530 38722 14542
rect 42478 14530 42530 14542
rect 39218 14478 39230 14530
rect 39282 14478 39294 14530
rect 41682 14478 41694 14530
rect 41746 14478 41758 14530
rect 38670 14466 38722 14478
rect 35646 14427 35698 14439
rect 39050 14422 39062 14474
rect 39114 14422 39126 14474
rect 42478 14466 42530 14478
rect 43038 14530 43090 14542
rect 43038 14466 43090 14478
rect 43262 14530 43314 14542
rect 46062 14530 46114 14542
rect 43362 14478 43374 14530
rect 43426 14478 43438 14530
rect 43262 14466 43314 14478
rect 12126 14362 12178 14374
rect 4846 14306 4898 14318
rect 4846 14242 4898 14254
rect 11454 14306 11506 14318
rect 18106 14366 18118 14418
rect 18170 14366 18182 14418
rect 16158 14354 16210 14366
rect 17378 14310 17390 14362
rect 17442 14310 17454 14362
rect 19518 14354 19570 14366
rect 44942 14418 44994 14430
rect 45173 14422 45185 14474
rect 45237 14422 45249 14474
rect 46062 14466 46114 14478
rect 46398 14530 46450 14542
rect 46398 14466 46450 14478
rect 29810 14310 29822 14362
rect 29874 14310 29886 14362
rect 35970 14310 35982 14362
rect 36034 14310 36046 14362
rect 12126 14298 12178 14310
rect 37998 14306 38050 14318
rect 39218 14310 39230 14362
rect 39282 14310 39294 14362
rect 44942 14354 44994 14366
rect 11454 14242 11506 14254
rect 37998 14242 38050 14254
rect 1344 14138 49616 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 49616 14138
rect 1344 14052 49616 14086
rect 8038 13970 8090 13982
rect 7410 13862 7422 13914
rect 7474 13862 7486 13914
rect 8038 13906 8090 13918
rect 19070 13970 19122 13982
rect 9650 13862 9662 13914
rect 9714 13862 9726 13914
rect 19070 13906 19122 13918
rect 40238 13970 40290 13982
rect 13806 13858 13858 13870
rect 22430 13858 22482 13870
rect 33730 13862 33742 13914
rect 33794 13862 33806 13914
rect 40238 13906 40290 13918
rect 41974 13970 42026 13982
rect 41974 13906 42026 13918
rect 2606 13746 2658 13758
rect 2606 13682 2658 13694
rect 5294 13746 5346 13758
rect 6066 13738 6078 13790
rect 6130 13738 6142 13790
rect 6974 13746 7026 13758
rect 7186 13750 7198 13802
rect 7250 13750 7262 13802
rect 13806 13794 13858 13806
rect 16494 13802 16546 13814
rect 9102 13746 9154 13758
rect 6402 13694 6414 13746
rect 6466 13694 6478 13746
rect 7522 13694 7534 13746
rect 7586 13694 7598 13746
rect 7858 13694 7870 13746
rect 7922 13694 7934 13746
rect 9538 13694 9550 13746
rect 9602 13694 9614 13746
rect 9874 13721 9886 13773
rect 9938 13721 9950 13773
rect 10222 13746 10274 13758
rect 5294 13682 5346 13694
rect 6974 13682 7026 13694
rect 9102 13682 9154 13694
rect 10222 13682 10274 13694
rect 11118 13746 11170 13758
rect 22430 13794 22482 13806
rect 35310 13858 35362 13870
rect 47394 13862 47406 13914
rect 47458 13862 47470 13914
rect 11890 13694 11902 13746
rect 11954 13694 11966 13746
rect 16494 13738 16546 13750
rect 17838 13746 17890 13758
rect 18118 13746 18170 13758
rect 16594 13694 16606 13746
rect 16658 13694 16670 13746
rect 17938 13694 17950 13746
rect 18002 13694 18014 13746
rect 11118 13682 11170 13694
rect 17838 13682 17890 13694
rect 18118 13682 18170 13694
rect 19406 13746 19458 13758
rect 19406 13682 19458 13694
rect 19742 13746 19794 13758
rect 20514 13694 20526 13746
rect 20578 13694 20590 13746
rect 22866 13727 22878 13779
rect 22930 13727 22942 13779
rect 23202 13750 23214 13802
rect 23266 13750 23278 13802
rect 23762 13750 23774 13802
rect 23826 13750 23838 13802
rect 23960 13734 23972 13786
rect 24024 13734 24036 13786
rect 25528 13784 25580 13796
rect 25230 13746 25282 13758
rect 25330 13694 25342 13746
rect 25394 13694 25406 13746
rect 25528 13720 25580 13732
rect 26798 13746 26850 13758
rect 19742 13682 19794 13694
rect 25230 13682 25282 13694
rect 26798 13682 26850 13694
rect 32622 13746 32674 13758
rect 34066 13750 34078 13802
rect 34130 13750 34142 13802
rect 35310 13794 35362 13806
rect 34302 13746 34354 13758
rect 37998 13746 38050 13758
rect 33618 13694 33630 13746
rect 33682 13694 33694 13746
rect 37202 13694 37214 13746
rect 37266 13694 37278 13746
rect 32622 13682 32674 13694
rect 34302 13682 34354 13694
rect 37998 13682 38050 13694
rect 38782 13746 38834 13758
rect 38782 13682 38834 13694
rect 38894 13746 38946 13758
rect 39330 13738 39342 13790
rect 39394 13738 39406 13790
rect 39902 13746 39954 13758
rect 39666 13694 39678 13746
rect 39730 13694 39742 13746
rect 38894 13682 38946 13694
rect 39902 13682 39954 13694
rect 42142 13746 42194 13758
rect 42142 13682 42194 13694
rect 42926 13746 42978 13758
rect 42926 13682 42978 13694
rect 45950 13746 46002 13758
rect 45950 13682 46002 13694
rect 46174 13746 46226 13758
rect 47170 13694 47182 13746
rect 47234 13694 47246 13746
rect 47506 13721 47518 13773
rect 47570 13721 47582 13773
rect 47854 13746 47906 13758
rect 46174 13682 46226 13694
rect 47854 13682 47906 13694
rect 48638 13746 48690 13758
rect 48638 13682 48690 13694
rect 48862 13746 48914 13758
rect 48862 13682 48914 13694
rect 3378 13582 3390 13634
rect 3442 13582 3454 13634
rect 5954 13582 5966 13634
rect 6018 13582 6030 13634
rect 16774 13578 16826 13590
rect 23986 13582 23998 13634
rect 24050 13582 24062 13634
rect 27570 13582 27582 13634
rect 27634 13582 27646 13634
rect 29474 13582 29486 13634
rect 29538 13582 29550 13634
rect 39218 13582 39230 13634
rect 39282 13582 39294 13634
rect 43698 13582 43710 13634
rect 43762 13582 43774 13634
rect 45602 13582 45614 13634
rect 45666 13582 45678 13634
rect 49130 13582 49142 13634
rect 49194 13582 49206 13634
rect 8766 13522 8818 13534
rect 8766 13458 8818 13470
rect 16326 13522 16378 13534
rect 16774 13514 16826 13526
rect 18510 13522 18562 13534
rect 16326 13458 16378 13470
rect 18510 13458 18562 13470
rect 25902 13522 25954 13534
rect 25902 13458 25954 13470
rect 32286 13522 32338 13534
rect 42478 13522 42530 13534
rect 38490 13470 38502 13522
rect 38554 13470 38566 13522
rect 46442 13470 46454 13522
rect 46506 13470 46518 13522
rect 32286 13458 32338 13470
rect 42478 13458 42530 13470
rect 1344 13354 49616 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 49616 13354
rect 1344 13268 49616 13302
rect 3390 13186 3442 13198
rect 21422 13186 21474 13198
rect 3390 13122 3442 13134
rect 7310 13130 7362 13142
rect 7802 13134 7814 13186
rect 7866 13134 7878 13186
rect 2550 13074 2602 13086
rect 21422 13122 21474 13134
rect 23102 13186 23154 13198
rect 23102 13122 23154 13134
rect 27918 13186 27970 13198
rect 27918 13122 27970 13134
rect 4610 13022 4622 13074
rect 4674 13022 4686 13074
rect 7310 13066 7362 13078
rect 18062 13074 18114 13086
rect 9202 13022 9214 13074
rect 9266 13022 9278 13074
rect 16370 13022 16382 13074
rect 16434 13022 16446 13074
rect 19182 13074 19234 13086
rect 2550 13010 2602 13022
rect 18062 13010 18114 13022
rect 18230 13018 18282 13030
rect 3726 12962 3778 12974
rect 2706 12910 2718 12962
rect 2770 12910 2782 12962
rect 3726 12898 3778 12910
rect 4398 12962 4450 12974
rect 6302 12962 6354 12974
rect 8094 12962 8146 12974
rect 5058 12910 5070 12962
rect 5122 12910 5134 12962
rect 5618 12910 5630 12962
rect 5682 12910 5694 12962
rect 4398 12898 4450 12910
rect 4778 12854 4790 12906
rect 4842 12854 4854 12906
rect 5954 12883 5966 12935
rect 6018 12883 6030 12935
rect 6962 12910 6974 12962
rect 7026 12910 7038 12962
rect 7186 12910 7198 12962
rect 7250 12910 7262 12962
rect 6302 12898 6354 12910
rect 8094 12898 8146 12910
rect 8318 12962 8370 12974
rect 8318 12898 8370 12910
rect 8430 12962 8482 12974
rect 12462 12962 12514 12974
rect 11890 12910 11902 12962
rect 11954 12910 11966 12962
rect 8430 12898 8482 12910
rect 12114 12883 12126 12935
rect 12178 12883 12190 12935
rect 12462 12898 12514 12910
rect 13694 12962 13746 12974
rect 19182 13010 19234 13022
rect 26742 13074 26794 13086
rect 39398 13074 39450 13086
rect 30370 13022 30382 13074
rect 30434 13022 30446 13074
rect 31826 13022 31838 13074
rect 31890 13022 31902 13074
rect 33730 13022 33742 13074
rect 33794 13022 33806 13074
rect 37762 13022 37774 13074
rect 37826 13022 37838 13074
rect 26742 13010 26794 13022
rect 39398 13010 39450 13022
rect 39902 13074 39954 13086
rect 43810 13022 43822 13074
rect 43874 13022 43886 13074
rect 39902 13010 39954 13022
rect 45670 13018 45722 13030
rect 14466 12910 14478 12962
rect 14530 12910 14542 12962
rect 17502 12924 17554 12936
rect 13694 12898 13746 12910
rect 17826 12910 17838 12962
rect 17890 12910 17902 12962
rect 18230 12954 18282 12966
rect 18510 12962 18562 12974
rect 19966 12962 20018 12974
rect 18610 12910 18622 12962
rect 18674 12910 18686 12962
rect 18510 12898 18562 12910
rect 11118 12850 11170 12862
rect 17502 12860 17554 12872
rect 18778 12854 18790 12906
rect 18842 12854 18854 12906
rect 19966 12898 20018 12910
rect 20302 12962 20354 12974
rect 20302 12898 20354 12910
rect 21758 12962 21810 12974
rect 21758 12898 21810 12910
rect 22430 12962 22482 12974
rect 22430 12898 22482 12910
rect 22766 12962 22818 12974
rect 22766 12898 22818 12910
rect 23438 12962 23490 12974
rect 28254 12962 28306 12974
rect 29374 12962 29426 12974
rect 31054 12962 31106 12974
rect 34862 12962 34914 12974
rect 24210 12910 24222 12962
rect 24274 12910 24286 12962
rect 28354 12910 28366 12962
rect 28418 12910 28430 12962
rect 23438 12898 23490 12910
rect 28254 12898 28306 12910
rect 29374 12898 29426 12910
rect 29698 12883 29710 12935
rect 29762 12883 29774 12935
rect 30034 12910 30046 12962
rect 30098 12910 30110 12962
rect 30482 12895 30494 12947
rect 30546 12895 30558 12947
rect 30706 12910 30718 12962
rect 30770 12910 30782 12962
rect 34178 12910 34190 12962
rect 34242 12910 34254 12962
rect 31054 12898 31106 12910
rect 4062 12738 4114 12750
rect 5730 12742 5742 12794
rect 5794 12742 5806 12794
rect 11118 12786 11170 12798
rect 26126 12850 26178 12862
rect 34458 12854 34470 12906
rect 34522 12854 34534 12906
rect 34862 12898 34914 12910
rect 35982 12962 36034 12974
rect 38334 12962 38386 12974
rect 37314 12910 37326 12962
rect 37378 12910 37390 12962
rect 35982 12898 36034 12910
rect 37650 12866 37662 12918
rect 37714 12866 37726 12918
rect 38334 12898 38386 12910
rect 38558 12962 38610 12974
rect 38558 12898 38610 12910
rect 39566 12962 39618 12974
rect 39566 12898 39618 12910
rect 41358 12962 41410 12974
rect 42254 12962 42306 12974
rect 41682 12910 41694 12962
rect 41746 12910 41758 12962
rect 41358 12898 41410 12910
rect 41906 12895 41918 12947
rect 41970 12895 41982 12947
rect 42254 12898 42306 12910
rect 42478 12962 42530 12974
rect 42478 12898 42530 12910
rect 43598 12962 43650 12974
rect 45502 12962 45554 12974
rect 43598 12898 43650 12910
rect 43922 12895 43934 12947
rect 43986 12895 43998 12947
rect 44258 12910 44270 12962
rect 44322 12910 44334 12962
rect 44942 12906 44994 12918
rect 45266 12910 45278 12962
rect 45330 12910 45342 12962
rect 45670 12954 45722 12966
rect 49310 12962 49362 12974
rect 48514 12910 48526 12962
rect 48578 12910 48590 12962
rect 45502 12898 45554 12910
rect 49310 12898 49362 12910
rect 38826 12798 38838 12850
rect 38890 12798 38902 12850
rect 12002 12742 12014 12794
rect 12066 12742 12078 12794
rect 26126 12786 26178 12798
rect 41918 12794 41970 12806
rect 42746 12798 42758 12850
rect 42810 12798 42822 12850
rect 44942 12842 44994 12854
rect 46622 12850 46674 12862
rect 4062 12674 4114 12686
rect 22094 12738 22146 12750
rect 29250 12742 29262 12794
rect 29314 12742 29326 12794
rect 34290 12742 34302 12794
rect 34354 12742 34366 12794
rect 22094 12674 22146 12686
rect 36318 12738 36370 12750
rect 36318 12674 36370 12686
rect 40518 12738 40570 12750
rect 40518 12674 40570 12686
rect 41022 12738 41074 12750
rect 46622 12786 46674 12798
rect 41918 12730 41970 12742
rect 43262 12738 43314 12750
rect 41022 12674 41074 12686
rect 43262 12674 43314 12686
rect 1344 12570 49616 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 49616 12570
rect 1344 12484 49616 12518
rect 6414 12402 6466 12414
rect 6414 12338 6466 12350
rect 9718 12402 9770 12414
rect 9718 12338 9770 12350
rect 26742 12402 26794 12414
rect 10210 12294 10222 12346
rect 10274 12294 10286 12346
rect 26742 12338 26794 12350
rect 32566 12402 32618 12414
rect 32566 12338 32618 12350
rect 48974 12402 49026 12414
rect 18062 12290 18114 12302
rect 24446 12290 24498 12302
rect 13178 12238 13190 12290
rect 13242 12238 13254 12290
rect 17502 12234 17554 12246
rect 1598 12178 1650 12190
rect 1598 12114 1650 12126
rect 4286 12178 4338 12190
rect 4946 12153 4958 12205
rect 5010 12153 5022 12205
rect 7534 12178 7586 12190
rect 4286 12114 4338 12126
rect 7534 12114 7586 12126
rect 7646 12178 7698 12190
rect 8642 12126 8654 12178
rect 8706 12126 8718 12178
rect 8866 12170 8878 12222
rect 8930 12170 8942 12222
rect 11006 12178 11058 12190
rect 10434 12126 10446 12178
rect 10498 12126 10510 12178
rect 11554 12126 11566 12178
rect 11618 12126 11630 12178
rect 11890 12153 11902 12205
rect 11954 12153 11966 12205
rect 12238 12178 12290 12190
rect 7646 12114 7698 12126
rect 11006 12114 11058 12126
rect 12238 12114 12290 12126
rect 12798 12178 12850 12190
rect 12798 12114 12850 12126
rect 12910 12178 12962 12190
rect 12910 12114 12962 12126
rect 14030 12178 14082 12190
rect 18062 12226 18114 12238
rect 18230 12234 18282 12246
rect 21914 12238 21926 12290
rect 21978 12238 21990 12290
rect 23774 12234 23826 12246
rect 17502 12170 17554 12182
rect 18808 12215 18860 12227
rect 17826 12126 17838 12178
rect 17890 12126 17902 12178
rect 18230 12170 18282 12182
rect 18510 12178 18562 12190
rect 18610 12126 18622 12178
rect 18674 12126 18686 12178
rect 18808 12151 18860 12163
rect 19574 12178 19626 12190
rect 20178 12154 20190 12206
rect 20242 12154 20254 12206
rect 21310 12178 21362 12190
rect 14030 12114 14082 12126
rect 18510 12114 18562 12126
rect 19574 12114 19626 12126
rect 19182 12066 19234 12078
rect 2370 12014 2382 12066
rect 2434 12014 2446 12066
rect 7914 12014 7926 12066
rect 7978 12014 7990 12066
rect 8978 12014 8990 12066
rect 9042 12014 9054 12066
rect 11666 12014 11678 12066
rect 11730 12014 11742 12066
rect 14802 12014 14814 12066
rect 14866 12014 14878 12066
rect 16706 12014 16718 12066
rect 16770 12014 16782 12066
rect 19182 12002 19234 12014
rect 19742 12066 19794 12078
rect 20402 12070 20414 12122
rect 20466 12070 20478 12122
rect 21310 12114 21362 12126
rect 21422 12178 21474 12190
rect 21422 12114 21474 12126
rect 21646 12178 21698 12190
rect 22922 12182 22934 12234
rect 22986 12182 22998 12234
rect 23986 12182 23998 12234
rect 24050 12182 24062 12234
rect 24446 12226 24498 12238
rect 27582 12290 27634 12302
rect 27582 12226 27634 12238
rect 45838 12290 45890 12302
rect 47842 12294 47854 12346
rect 47906 12294 47918 12346
rect 48974 12338 49026 12350
rect 45838 12226 45890 12238
rect 23090 12126 23102 12178
rect 23154 12126 23166 12178
rect 23774 12170 23826 12182
rect 25454 12178 25506 12190
rect 21646 12114 21698 12126
rect 23494 12122 23546 12134
rect 19742 12002 19794 12014
rect 23326 12066 23378 12078
rect 23494 12058 23546 12070
rect 24614 12122 24666 12134
rect 25454 12114 25506 12126
rect 25790 12178 25842 12190
rect 27246 12178 27298 12190
rect 26114 12126 26126 12178
rect 26178 12126 26190 12178
rect 26562 12126 26574 12178
rect 26626 12126 26638 12178
rect 28130 12126 28142 12178
rect 28194 12126 28206 12178
rect 28354 12170 28366 12222
rect 28418 12170 28430 12222
rect 29138 12153 29150 12205
rect 29202 12153 29214 12205
rect 31502 12178 31554 12190
rect 25790 12114 25842 12126
rect 27246 12114 27298 12126
rect 31502 12114 31554 12126
rect 31726 12178 31778 12190
rect 32958 12178 33010 12190
rect 31994 12126 32006 12178
rect 32058 12126 32070 12178
rect 31726 12114 31778 12126
rect 32958 12114 33010 12126
rect 35982 12178 36034 12190
rect 39006 12178 39058 12190
rect 36754 12126 36766 12178
rect 36818 12126 36830 12178
rect 35982 12114 36034 12126
rect 39006 12114 39058 12126
rect 39230 12178 39282 12190
rect 39230 12114 39282 12126
rect 39790 12178 39842 12190
rect 39790 12114 39842 12126
rect 42030 12178 42082 12190
rect 42030 12114 42082 12126
rect 42142 12178 42194 12190
rect 42578 12170 42590 12222
rect 42642 12170 42654 12222
rect 43150 12178 43202 12190
rect 42802 12126 42814 12178
rect 42866 12126 42878 12178
rect 43922 12126 43934 12178
rect 43986 12126 43998 12178
rect 46274 12126 46286 12178
rect 46338 12126 46350 12178
rect 46610 12141 46622 12193
rect 46674 12141 46686 12193
rect 47170 12126 47182 12178
rect 47234 12126 47246 12178
rect 47394 12153 47406 12205
rect 47458 12153 47470 12205
rect 47742 12178 47794 12190
rect 42142 12114 42194 12126
rect 43150 12114 43202 12126
rect 47742 12114 47794 12126
rect 48638 12178 48690 12190
rect 48638 12114 48690 12126
rect 24614 12058 24666 12070
rect 41414 12066 41466 12078
rect 28466 12014 28478 12066
rect 28530 12014 28542 12066
rect 33730 12014 33742 12066
rect 33794 12014 33806 12066
rect 35634 12014 35646 12066
rect 35698 12014 35710 12066
rect 38658 12014 38670 12066
rect 38722 12014 38734 12066
rect 42466 12014 42478 12066
rect 42530 12014 42542 12066
rect 46722 12014 46734 12066
rect 46786 12014 46798 12066
rect 23326 12002 23378 12014
rect 41414 12002 41466 12014
rect 20974 11954 21026 11966
rect 20974 11890 21026 11902
rect 26294 11954 26346 11966
rect 26294 11890 26346 11902
rect 29822 11954 29874 11966
rect 40126 11954 40178 11966
rect 39498 11902 39510 11954
rect 39562 11902 39574 11954
rect 41738 11902 41750 11954
rect 41802 11902 41814 11954
rect 29822 11890 29874 11902
rect 40126 11890 40178 11902
rect 1344 11786 49616 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 49616 11786
rect 1344 11700 49616 11734
rect 2382 11618 2434 11630
rect 19742 11618 19794 11630
rect 32622 11618 32674 11630
rect 2382 11554 2434 11566
rect 7198 11562 7250 11574
rect 18106 11566 18118 11618
rect 18170 11566 18182 11618
rect 21690 11566 21702 11618
rect 21754 11566 21766 11618
rect 34682 11566 34694 11618
rect 34746 11566 34758 11618
rect 48234 11566 48246 11618
rect 48298 11566 48310 11618
rect 19742 11554 19794 11566
rect 32622 11554 32674 11566
rect 3490 11454 3502 11506
rect 3554 11454 3566 11506
rect 5730 11454 5742 11506
rect 5794 11454 5806 11506
rect 7198 11498 7250 11510
rect 15878 11506 15930 11518
rect 14242 11454 14254 11506
rect 14306 11454 14318 11506
rect 15878 11442 15930 11454
rect 16326 11506 16378 11518
rect 16326 11442 16378 11454
rect 18622 11506 18674 11518
rect 23538 11454 23550 11506
rect 23602 11454 23614 11506
rect 25442 11454 25454 11506
rect 25506 11454 25518 11506
rect 31714 11454 31726 11506
rect 31778 11454 31790 11506
rect 40114 11454 40126 11506
rect 40178 11454 40190 11506
rect 18622 11442 18674 11454
rect 2718 11394 2770 11406
rect 4062 11394 4114 11406
rect 6302 11394 6354 11406
rect 3154 11342 3166 11394
rect 3218 11342 3230 11394
rect 2718 11330 2770 11342
rect 3378 11298 3390 11350
rect 3442 11298 3454 11350
rect 4062 11330 4114 11342
rect 4286 11355 4338 11367
rect 4610 11342 4622 11394
rect 4674 11342 4686 11394
rect 5618 11342 5630 11394
rect 5682 11342 5694 11394
rect 4286 11291 4338 11303
rect 5954 11286 5966 11338
rect 6018 11286 6030 11338
rect 6302 11330 6354 11342
rect 6638 11394 6690 11406
rect 7870 11394 7922 11406
rect 7298 11342 7310 11394
rect 7362 11342 7374 11394
rect 7522 11342 7534 11394
rect 7586 11342 7598 11394
rect 6638 11330 6690 11342
rect 7870 11330 7922 11342
rect 8542 11394 8594 11406
rect 12574 11394 12626 11406
rect 9314 11342 9326 11394
rect 9378 11342 9390 11394
rect 11890 11342 11902 11394
rect 11954 11342 11966 11394
rect 12350 11355 12402 11367
rect 8542 11330 8594 11342
rect 12574 11330 12626 11342
rect 13806 11394 13858 11406
rect 13806 11330 13858 11342
rect 13918 11394 13970 11406
rect 16942 11394 16994 11406
rect 13918 11330 13970 11342
rect 14354 11327 14366 11379
rect 14418 11327 14430 11379
rect 14578 11342 14590 11394
rect 14642 11342 14654 11394
rect 16818 11342 16830 11394
rect 16882 11342 16894 11394
rect 16942 11330 16994 11342
rect 17614 11394 17666 11406
rect 17614 11330 17666 11342
rect 17838 11394 17890 11406
rect 17838 11330 17890 11342
rect 19016 11394 19068 11406
rect 19294 11394 19346 11406
rect 19170 11342 19182 11394
rect 19234 11342 19246 11394
rect 19016 11330 19068 11342
rect 19294 11330 19346 11342
rect 20078 11394 20130 11406
rect 20078 11330 20130 11342
rect 20414 11394 20466 11406
rect 20414 11330 20466 11342
rect 20750 11394 20802 11406
rect 20750 11330 20802 11342
rect 21982 11394 22034 11406
rect 21982 11330 22034 11342
rect 22094 11394 22146 11406
rect 22094 11330 22146 11342
rect 22766 11394 22818 11406
rect 22766 11330 22818 11342
rect 25790 11394 25842 11406
rect 29374 11394 29426 11406
rect 31166 11394 31218 11406
rect 32958 11394 33010 11406
rect 34302 11394 34354 11406
rect 26562 11342 26574 11394
rect 26626 11342 26638 11394
rect 25790 11330 25842 11342
rect 29374 11330 29426 11342
rect 29598 11355 29650 11367
rect 8206 11282 8258 11294
rect 3938 11174 3950 11226
rect 4002 11174 4014 11226
rect 8206 11218 8258 11230
rect 11230 11282 11282 11294
rect 12350 11291 12402 11303
rect 30034 11342 30046 11394
rect 30098 11342 30110 11394
rect 30482 11342 30494 11394
rect 30546 11342 30558 11394
rect 30942 11355 30994 11367
rect 28478 11282 28530 11294
rect 29598 11291 29650 11303
rect 31166 11330 31218 11342
rect 31826 11327 31838 11379
rect 31890 11327 31902 11379
rect 32162 11342 32174 11394
rect 32226 11342 32238 11394
rect 32958 11330 33010 11342
rect 30942 11291 30994 11303
rect 33618 11298 33630 11350
rect 33682 11298 33694 11350
rect 33954 11342 33966 11394
rect 34018 11342 34030 11394
rect 34302 11330 34354 11342
rect 34414 11394 34466 11406
rect 34414 11330 34466 11342
rect 36318 11394 36370 11406
rect 36318 11330 36370 11342
rect 36542 11394 36594 11406
rect 40910 11394 40962 11406
rect 36866 11342 36878 11394
rect 36930 11342 36942 11394
rect 36542 11330 36594 11342
rect 40910 11330 40962 11342
rect 41022 11394 41074 11406
rect 44718 11394 44770 11406
rect 47854 11394 47906 11406
rect 41794 11342 41806 11394
rect 41858 11342 41870 11394
rect 45490 11342 45502 11394
rect 45554 11342 45566 11394
rect 41022 11330 41074 11342
rect 44718 11330 44770 11342
rect 47854 11330 47906 11342
rect 47966 11394 48018 11406
rect 47966 11330 48018 11342
rect 48526 11394 48578 11406
rect 48526 11330 48578 11342
rect 38222 11282 38274 11294
rect 13514 11230 13526 11282
rect 13578 11230 13590 11282
rect 36026 11230 36038 11282
rect 36090 11230 36102 11282
rect 11230 11218 11282 11230
rect 12002 11174 12014 11226
rect 12066 11174 12078 11226
rect 28478 11218 28530 11230
rect 16662 11170 16714 11182
rect 16662 11106 16714 11118
rect 17278 11170 17330 11182
rect 29250 11174 29262 11226
rect 29314 11174 29326 11226
rect 31266 11174 31278 11226
rect 31330 11174 31342 11226
rect 33842 11174 33854 11226
rect 33906 11174 33918 11226
rect 38222 11218 38274 11230
rect 43710 11282 43762 11294
rect 43710 11218 43762 11230
rect 47406 11282 47458 11294
rect 47406 11218 47458 11230
rect 17278 11106 17330 11118
rect 35254 11170 35306 11182
rect 35254 11106 35306 11118
rect 35702 11170 35754 11182
rect 35702 11106 35754 11118
rect 44326 11170 44378 11182
rect 44326 11106 44378 11118
rect 48862 11170 48914 11182
rect 48862 11106 48914 11118
rect 1344 11002 49616 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 49616 11002
rect 1344 10916 49616 10950
rect 8094 10834 8146 10846
rect 8094 10770 8146 10782
rect 8878 10834 8930 10846
rect 8878 10770 8930 10782
rect 21142 10834 21194 10846
rect 4286 10722 4338 10734
rect 9650 10726 9662 10778
rect 9714 10726 9726 10778
rect 21142 10770 21194 10782
rect 27806 10834 27858 10846
rect 4286 10658 4338 10670
rect 11230 10722 11282 10734
rect 25330 10726 25342 10778
rect 25394 10726 25406 10778
rect 27806 10770 27858 10782
rect 34358 10834 34410 10846
rect 34358 10770 34410 10782
rect 36766 10834 36818 10846
rect 36766 10770 36818 10782
rect 39554 10726 39566 10778
rect 39618 10726 39630 10778
rect 43038 10722 43090 10734
rect 11230 10658 11282 10670
rect 17558 10666 17610 10678
rect 1598 10610 1650 10622
rect 5070 10610 5122 10622
rect 4778 10558 4790 10610
rect 4842 10558 4854 10610
rect 1598 10546 1650 10558
rect 5070 10546 5122 10558
rect 5294 10610 5346 10622
rect 5294 10546 5346 10558
rect 5854 10610 5906 10622
rect 5854 10546 5906 10558
rect 5966 10610 6018 10622
rect 5966 10546 6018 10558
rect 6190 10610 6242 10622
rect 6190 10546 6242 10558
rect 6414 10610 6466 10622
rect 6414 10546 6466 10558
rect 7534 10610 7586 10622
rect 7534 10546 7586 10558
rect 8430 10610 8482 10622
rect 8430 10546 8482 10558
rect 8542 10610 8594 10622
rect 8542 10546 8594 10558
rect 9774 10610 9826 10622
rect 10098 10585 10110 10637
rect 10162 10585 10174 10637
rect 13918 10610 13970 10622
rect 10434 10558 10446 10610
rect 10498 10558 10510 10610
rect 9774 10546 9826 10558
rect 13918 10546 13970 10558
rect 14030 10610 14082 10622
rect 17558 10602 17610 10614
rect 18286 10666 18338 10678
rect 29082 10670 29094 10722
rect 29146 10670 29158 10722
rect 33450 10670 33462 10722
rect 33514 10670 33526 10722
rect 17938 10558 17950 10610
rect 18002 10558 18014 10610
rect 18286 10602 18338 10614
rect 18734 10610 18786 10622
rect 18834 10558 18846 10610
rect 18898 10558 18910 10610
rect 18992 10608 19004 10660
rect 19056 10608 19068 10660
rect 20340 10648 20392 10660
rect 21680 10648 21732 10660
rect 20638 10610 20690 10622
rect 20340 10584 20392 10596
rect 20514 10558 20526 10610
rect 20578 10558 20590 10610
rect 14030 10546 14082 10558
rect 18734 10546 18786 10558
rect 20638 10546 20690 10558
rect 21422 10610 21474 10622
rect 21522 10558 21534 10610
rect 21586 10558 21598 10610
rect 21680 10584 21732 10596
rect 22486 10610 22538 10622
rect 22866 10558 22878 10610
rect 22930 10558 22942 10610
rect 23090 10586 23102 10638
rect 23154 10586 23166 10638
rect 24164 10608 24176 10660
rect 24228 10608 24240 10660
rect 24446 10610 24498 10622
rect 24322 10558 24334 10610
rect 24386 10558 24398 10610
rect 21422 10546 21474 10558
rect 22486 10546 22538 10558
rect 24446 10546 24498 10558
rect 25454 10610 25506 10622
rect 25666 10614 25678 10666
rect 25730 10614 25742 10666
rect 43038 10658 43090 10670
rect 28142 10610 28194 10622
rect 26114 10558 26126 10610
rect 26178 10558 26190 10610
rect 26338 10558 26350 10610
rect 26402 10558 26414 10610
rect 25454 10546 25506 10558
rect 28142 10546 28194 10558
rect 28590 10610 28642 10622
rect 28590 10546 28642 10558
rect 28814 10610 28866 10622
rect 28814 10546 28866 10558
rect 29374 10610 29426 10622
rect 29374 10546 29426 10558
rect 32062 10610 32114 10622
rect 32062 10546 32114 10558
rect 32958 10610 33010 10622
rect 32958 10546 33010 10558
rect 33182 10610 33234 10622
rect 34626 10558 34638 10610
rect 34690 10558 34702 10610
rect 34962 10573 34974 10625
rect 35026 10573 35038 10625
rect 35298 10558 35310 10610
rect 35362 10558 35374 10610
rect 38434 10585 38446 10637
rect 38498 10585 38510 10637
rect 39006 10610 39058 10622
rect 39330 10585 39342 10637
rect 39394 10585 39406 10637
rect 39902 10610 39954 10622
rect 39666 10558 39678 10610
rect 39730 10558 39742 10610
rect 41010 10573 41022 10625
rect 41074 10573 41086 10625
rect 42124 10610 42176 10622
rect 41234 10558 41246 10610
rect 41298 10558 41310 10610
rect 33182 10546 33234 10558
rect 39006 10546 39058 10558
rect 39902 10546 39954 10558
rect 42124 10546 42176 10558
rect 42366 10610 42418 10622
rect 43374 10610 43426 10622
rect 42366 10546 42418 10558
rect 42870 10554 42922 10566
rect 17726 10498 17778 10510
rect 2370 10446 2382 10498
rect 2434 10446 2446 10498
rect 13122 10446 13134 10498
rect 13186 10446 13198 10498
rect 14802 10446 14814 10498
rect 14866 10446 14878 10498
rect 16706 10446 16718 10498
rect 16770 10446 16782 10498
rect 17726 10434 17778 10446
rect 22094 10498 22146 10510
rect 22094 10434 22146 10446
rect 22654 10498 22706 10510
rect 22654 10434 22706 10446
rect 23774 10498 23826 10510
rect 43922 10558 43934 10610
rect 43986 10558 43998 10610
rect 44594 10602 44606 10654
rect 44658 10602 44670 10654
rect 44930 10558 44942 10610
rect 44994 10558 45006 10610
rect 47394 10585 47406 10637
rect 47458 10585 47470 10637
rect 48246 10610 48298 10622
rect 43374 10546 43426 10558
rect 48246 10546 48298 10558
rect 48638 10610 48690 10622
rect 48638 10546 48690 10558
rect 23774 10434 23826 10446
rect 26518 10442 26570 10454
rect 30146 10446 30158 10498
rect 30210 10446 30222 10498
rect 35074 10446 35086 10498
rect 35138 10446 35150 10498
rect 40898 10446 40910 10498
rect 40962 10446 40974 10498
rect 41570 10446 41582 10498
rect 41634 10495 41646 10498
rect 41794 10495 41806 10498
rect 41634 10449 41806 10495
rect 41634 10446 41646 10449
rect 41794 10446 41806 10449
rect 41858 10446 41870 10498
rect 42870 10490 42922 10502
rect 44482 10446 44494 10498
rect 44546 10446 44558 10498
rect 7198 10386 7250 10398
rect 5562 10334 5574 10386
rect 5626 10334 5638 10386
rect 6682 10334 6694 10386
rect 6746 10334 6758 10386
rect 7198 10322 7250 10334
rect 19406 10386 19458 10398
rect 19406 10322 19458 10334
rect 19966 10386 20018 10398
rect 26518 10378 26570 10390
rect 35478 10386 35530 10398
rect 19966 10322 20018 10334
rect 35478 10322 35530 10334
rect 40238 10386 40290 10398
rect 44146 10390 44158 10442
rect 44210 10390 44222 10442
rect 40238 10322 40290 10334
rect 46062 10386 46114 10398
rect 46062 10322 46114 10334
rect 48974 10386 49026 10398
rect 48974 10322 49026 10334
rect 1344 10218 49616 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 49616 10218
rect 1344 10132 49616 10166
rect 2382 10050 2434 10062
rect 2382 9986 2434 9998
rect 30494 10050 30546 10062
rect 30494 9986 30546 9998
rect 34862 10050 34914 10062
rect 41470 10050 41522 10062
rect 36250 9998 36262 10050
rect 36314 9998 36326 10050
rect 34862 9986 34914 9998
rect 41470 9986 41522 9998
rect 21422 9938 21474 9950
rect 37158 9938 37210 9950
rect 12338 9886 12350 9938
rect 12402 9886 12414 9938
rect 19686 9882 19738 9894
rect 2718 9826 2770 9838
rect 2718 9762 2770 9774
rect 3726 9826 3778 9838
rect 6302 9826 6354 9838
rect 3726 9762 3778 9774
rect 3950 9787 4002 9799
rect 4274 9774 4286 9826
rect 4338 9774 4350 9826
rect 5618 9774 5630 9826
rect 5682 9774 5694 9826
rect 10782 9826 10834 9838
rect 14366 9826 14418 9838
rect 17726 9826 17778 9838
rect 23650 9886 23662 9938
rect 23714 9886 23726 9938
rect 25554 9886 25566 9938
rect 25618 9886 25630 9938
rect 28130 9886 28142 9938
rect 28194 9886 28206 9938
rect 21422 9874 21474 9886
rect 37158 9874 37210 9886
rect 38334 9938 38386 9950
rect 38334 9874 38386 9886
rect 40294 9938 40346 9950
rect 48638 9938 48690 9950
rect 45490 9886 45502 9938
rect 45554 9886 45566 9938
rect 47394 9886 47406 9938
rect 47458 9886 47470 9938
rect 40294 9874 40346 9886
rect 48638 9874 48690 9886
rect 3950 9723 4002 9735
rect 6066 9718 6078 9770
rect 6130 9718 6142 9770
rect 6302 9762 6354 9774
rect 7298 9741 7310 9793
rect 7362 9741 7374 9793
rect 7746 9718 7758 9770
rect 7810 9718 7822 9770
rect 8082 9718 8094 9770
rect 8146 9718 8158 9770
rect 8392 9741 8404 9793
rect 8456 9741 8468 9793
rect 11330 9774 11342 9826
rect 11394 9774 11406 9826
rect 11890 9774 11902 9826
rect 11954 9774 11966 9826
rect 10782 9762 10834 9774
rect 12226 9759 12238 9811
rect 12290 9759 12302 9811
rect 13570 9774 13582 9826
rect 13634 9774 13646 9826
rect 15138 9774 15150 9826
rect 15202 9774 15214 9826
rect 18274 9774 18286 9826
rect 18338 9774 18350 9826
rect 18958 9788 19010 9800
rect 14366 9762 14418 9774
rect 17726 9762 17778 9774
rect 8542 9714 8594 9726
rect 3602 9606 3614 9658
rect 3666 9606 3678 9658
rect 6402 9606 6414 9658
rect 6466 9606 6478 9658
rect 8542 9650 8594 9662
rect 17054 9714 17106 9726
rect 18050 9718 18062 9770
rect 18114 9718 18126 9770
rect 19282 9774 19294 9826
rect 19346 9774 19358 9826
rect 19686 9818 19738 9830
rect 20806 9826 20858 9838
rect 20178 9746 20190 9798
rect 20242 9746 20254 9798
rect 20402 9774 20414 9826
rect 20466 9774 20478 9826
rect 20806 9762 20858 9774
rect 21814 9826 21866 9838
rect 22094 9826 22146 9838
rect 22878 9826 22930 9838
rect 21970 9774 21982 9826
rect 22034 9774 22046 9826
rect 22306 9774 22318 9826
rect 22370 9774 22382 9826
rect 21814 9762 21866 9774
rect 22094 9762 22146 9774
rect 22878 9762 22930 9774
rect 27582 9826 27634 9838
rect 30830 9826 30882 9838
rect 27582 9762 27634 9774
rect 28242 9759 28254 9811
rect 28306 9759 28318 9811
rect 28578 9774 28590 9826
rect 28642 9774 28654 9826
rect 30830 9762 30882 9774
rect 31614 9826 31666 9838
rect 35254 9826 35306 9838
rect 35534 9826 35586 9838
rect 32478 9774 32490 9826
rect 32542 9774 32554 9826
rect 31614 9762 31666 9774
rect 33126 9770 33178 9782
rect 18958 9724 19010 9736
rect 11554 9606 11566 9658
rect 11618 9606 11630 9658
rect 17054 9650 17106 9662
rect 19518 9714 19570 9726
rect 17826 9606 17838 9658
rect 17890 9606 17902 9658
rect 19518 9650 19570 9662
rect 20638 9714 20690 9726
rect 20638 9650 20690 9662
rect 32734 9714 32786 9726
rect 33282 9718 33294 9770
rect 33346 9718 33358 9770
rect 33506 9735 33518 9787
rect 33570 9735 33582 9787
rect 35410 9774 35422 9826
rect 35474 9774 35486 9826
rect 35254 9762 35306 9774
rect 35534 9762 35586 9774
rect 35870 9826 35922 9838
rect 35870 9762 35922 9774
rect 35982 9826 36034 9838
rect 35982 9762 36034 9774
rect 37662 9826 37714 9838
rect 37662 9762 37714 9774
rect 37998 9826 38050 9838
rect 39678 9826 39730 9838
rect 37998 9762 38050 9774
rect 38222 9787 38274 9799
rect 38658 9774 38670 9826
rect 38722 9774 38734 9826
rect 38994 9774 39006 9826
rect 39058 9774 39070 9826
rect 39330 9747 39342 9799
rect 39394 9747 39406 9799
rect 39678 9762 39730 9774
rect 40574 9826 40626 9838
rect 40574 9762 40626 9774
rect 41022 9826 41074 9838
rect 33126 9706 33178 9718
rect 34078 9714 34130 9726
rect 38222 9723 38274 9735
rect 32734 9650 32786 9662
rect 34078 9650 34130 9662
rect 40686 9714 40738 9726
rect 40842 9718 40854 9770
rect 40906 9718 40918 9770
rect 41022 9762 41074 9774
rect 41806 9826 41858 9838
rect 41806 9762 41858 9774
rect 41918 9826 41970 9838
rect 43598 9826 43650 9838
rect 43306 9774 43318 9826
rect 43370 9774 43382 9826
rect 41918 9762 41970 9774
rect 43598 9762 43650 9774
rect 43822 9826 43874 9838
rect 43822 9762 43874 9774
rect 48190 9826 48242 9838
rect 48190 9762 48242 9774
rect 48302 9826 48354 9838
rect 48302 9762 48354 9774
rect 27246 9602 27298 9614
rect 39106 9606 39118 9658
rect 39170 9606 39182 9658
rect 40686 9650 40738 9662
rect 27246 9538 27298 9550
rect 42254 9602 42306 9614
rect 42254 9538 42306 9550
rect 42870 9602 42922 9614
rect 42870 9538 42922 9550
rect 44214 9602 44266 9614
rect 44214 9538 44266 9550
rect 44998 9602 45050 9614
rect 44998 9538 45050 9550
rect 49142 9602 49194 9614
rect 49142 9538 49194 9550
rect 1344 9434 49616 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 49616 9434
rect 1344 9348 49616 9382
rect 6582 9266 6634 9278
rect 4902 9210 4954 9222
rect 6582 9202 6634 9214
rect 7086 9266 7138 9278
rect 24726 9266 24778 9278
rect 7086 9202 7138 9214
rect 19910 9210 19962 9222
rect 4902 9146 4954 9158
rect 10894 9154 10946 9166
rect 5820 9080 5872 9092
rect 10894 9090 10946 9102
rect 19406 9154 19458 9166
rect 24726 9202 24778 9214
rect 48134 9210 48186 9222
rect 19910 9146 19962 9158
rect 28702 9154 28754 9166
rect 1598 9042 1650 9054
rect 1598 8978 1650 8990
rect 4286 9042 4338 9054
rect 4722 8990 4734 9042
rect 4786 8990 4798 9042
rect 6078 9042 6130 9054
rect 5820 9016 5872 9028
rect 5954 8990 5966 9042
rect 6018 8990 6030 9042
rect 4286 8978 4338 8990
rect 6078 8978 6130 8990
rect 7422 9042 7474 9054
rect 7422 8978 7474 8990
rect 8206 9042 8258 9054
rect 8206 8978 8258 8990
rect 8318 9042 8370 9054
rect 8318 8978 8370 8990
rect 9998 9042 10050 9054
rect 13582 9042 13634 9054
rect 12786 8990 12798 9042
rect 12850 8990 12862 9042
rect 9998 8978 10050 8990
rect 13582 8978 13634 8990
rect 14030 9042 14082 9054
rect 17278 9042 17330 9054
rect 18946 9046 18958 9098
rect 19010 9046 19022 9098
rect 19406 9090 19458 9102
rect 19574 9098 19626 9110
rect 28702 9090 28754 9102
rect 33406 9154 33458 9166
rect 33406 9090 33458 9102
rect 38894 9154 38946 9166
rect 38894 9090 38946 9102
rect 39510 9154 39562 9166
rect 39510 9090 39562 9102
rect 43486 9154 43538 9166
rect 48134 9146 48186 9158
rect 43486 9090 43538 9102
rect 14802 8990 14814 9042
rect 14866 8990 14878 9042
rect 17938 8990 17950 9042
rect 18002 8990 18014 9042
rect 19170 8990 19182 9042
rect 19234 8990 19246 9042
rect 19574 9034 19626 9046
rect 20526 9042 20578 9054
rect 24110 9042 24162 9054
rect 19730 8990 19742 9042
rect 19794 8990 19806 9042
rect 21298 8990 21310 9042
rect 21362 8990 21374 9042
rect 14030 8978 14082 8990
rect 17278 8978 17330 8990
rect 20526 8978 20578 8990
rect 24110 8978 24162 8990
rect 25118 9042 25170 9054
rect 25118 8978 25170 8990
rect 26014 9042 26066 9054
rect 29038 9042 29090 9054
rect 26786 8990 26798 9042
rect 26850 8990 26862 9042
rect 26014 8978 26066 8990
rect 29038 8978 29090 8990
rect 29262 9042 29314 9054
rect 29262 8978 29314 8990
rect 30830 9042 30882 9054
rect 31490 9005 31502 9057
rect 31554 9005 31566 9057
rect 36094 9042 36146 9054
rect 31826 8990 31838 9042
rect 31890 8990 31902 9042
rect 35298 8990 35310 9042
rect 35362 8990 35374 9042
rect 30830 8978 30882 8990
rect 36094 8978 36146 8990
rect 36206 9042 36258 9054
rect 36206 8978 36258 8990
rect 39790 9042 39842 9054
rect 40070 9042 40122 9054
rect 39890 8990 39902 9042
rect 39954 8990 39966 9042
rect 39790 8978 39842 8990
rect 40070 8978 40122 8990
rect 40238 9042 40290 9054
rect 40238 8978 40290 8990
rect 40798 9042 40850 9054
rect 43990 9042 44042 9054
rect 44258 9046 44270 9098
rect 44322 9046 44334 9098
rect 44494 9070 44546 9082
rect 41570 8990 41582 9042
rect 41634 8990 41646 9042
rect 44494 9006 44546 9018
rect 44718 9070 44770 9082
rect 44718 9006 44770 9018
rect 44830 9077 44882 9089
rect 44830 9013 44882 9025
rect 45602 9017 45614 9069
rect 45666 9017 45678 9069
rect 48638 9042 48690 9054
rect 40798 8978 40850 8990
rect 43990 8978 44042 8990
rect 48638 8978 48690 8990
rect 2370 8878 2382 8930
rect 2434 8878 2446 8930
rect 16706 8878 16718 8930
rect 16770 8878 16782 8930
rect 23202 8878 23214 8930
rect 23266 8878 23278 8930
rect 31378 8878 31390 8930
rect 31442 8878 31454 8930
rect 36978 8878 36990 8930
rect 37042 8878 37054 8930
rect 5406 8818 5458 8830
rect 5406 8754 5458 8766
rect 7870 8818 7922 8830
rect 7870 8754 7922 8766
rect 8654 8818 8706 8830
rect 8654 8754 8706 8766
rect 9662 8818 9714 8830
rect 9662 8754 9714 8766
rect 17614 8818 17666 8830
rect 17614 8754 17666 8766
rect 18118 8818 18170 8830
rect 18118 8754 18170 8766
rect 23774 8818 23826 8830
rect 23774 8754 23826 8766
rect 25454 8818 25506 8830
rect 30494 8818 30546 8830
rect 29530 8766 29542 8818
rect 29594 8766 29606 8818
rect 25454 8754 25506 8766
rect 30494 8754 30546 8766
rect 48974 8818 49026 8830
rect 48974 8754 49026 8766
rect 1344 8650 49616 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 49616 8650
rect 1344 8564 49616 8598
rect 21926 8482 21978 8494
rect 21926 8418 21978 8430
rect 23326 8482 23378 8494
rect 23326 8418 23378 8430
rect 37214 8482 37266 8494
rect 39274 8430 39286 8482
rect 39338 8430 39350 8482
rect 37214 8418 37266 8430
rect 4958 8370 5010 8382
rect 7254 8370 7306 8382
rect 4958 8306 5010 8318
rect 5126 8314 5178 8326
rect 7254 8306 7306 8318
rect 12798 8370 12850 8382
rect 44326 8370 44378 8382
rect 30034 8318 30046 8370
rect 30098 8318 30110 8370
rect 36306 8318 36318 8370
rect 36370 8318 36382 8370
rect 41122 8318 41134 8370
rect 41186 8318 41198 8370
rect 43026 8318 43038 8370
rect 43090 8318 43102 8370
rect 12798 8306 12850 8318
rect 44326 8306 44378 8318
rect 3378 8178 3390 8230
rect 3442 8178 3454 8230
rect 3602 8206 3614 8258
rect 3666 8206 3678 8258
rect 4398 8220 4450 8232
rect 4006 8202 4058 8214
rect 3838 8146 3890 8158
rect 4722 8206 4734 8258
rect 4786 8206 4798 8258
rect 5126 8250 5178 8262
rect 6302 8258 6354 8270
rect 5618 8206 5630 8258
rect 5682 8206 5694 8258
rect 4398 8156 4450 8168
rect 6066 8150 6078 8202
rect 6130 8150 6142 8202
rect 6302 8194 6354 8206
rect 7422 8258 7474 8270
rect 11230 8258 11282 8270
rect 12462 8258 12514 8270
rect 19854 8258 19906 8270
rect 8194 8206 8206 8258
rect 8258 8206 8270 8258
rect 10546 8206 10558 8258
rect 10610 8206 10622 8258
rect 12338 8206 12350 8258
rect 12402 8206 12414 8258
rect 13906 8206 13918 8258
rect 13970 8206 13982 8258
rect 7422 8194 7474 8206
rect 4006 8138 4058 8150
rect 10110 8146 10162 8158
rect 10882 8150 10894 8202
rect 10946 8150 10958 8202
rect 11230 8194 11282 8206
rect 12462 8194 12514 8206
rect 16146 8178 16158 8230
rect 16210 8178 16222 8230
rect 18610 8178 18622 8230
rect 18674 8178 18686 8230
rect 19854 8194 19906 8206
rect 20078 8258 20130 8270
rect 20078 8194 20130 8206
rect 20190 8258 20242 8270
rect 20190 8194 20242 8206
rect 21590 8258 21642 8270
rect 25006 8258 25058 8270
rect 22082 8206 22094 8258
rect 22146 8206 22158 8258
rect 21590 8194 21642 8206
rect 22306 8178 22318 8230
rect 22370 8178 22382 8230
rect 25006 8194 25058 8206
rect 25230 8258 25282 8270
rect 25230 8194 25282 8206
rect 26574 8258 26626 8270
rect 26574 8194 26626 8206
rect 26966 8258 27018 8270
rect 26966 8194 27018 8206
rect 27470 8258 27522 8270
rect 29262 8258 29314 8270
rect 28018 8206 28030 8258
rect 28082 8206 28094 8258
rect 27470 8194 27522 8206
rect 27794 8150 27806 8202
rect 27858 8150 27870 8202
rect 29262 8194 29314 8206
rect 32398 8258 32450 8270
rect 33854 8258 33906 8270
rect 33262 8206 33274 8258
rect 33326 8206 33338 8258
rect 32398 8194 32450 8206
rect 33854 8194 33906 8206
rect 34918 8258 34970 8270
rect 34918 8194 34970 8206
rect 35646 8258 35698 8270
rect 37550 8258 37602 8270
rect 35858 8206 35870 8258
rect 35922 8206 35934 8258
rect 36150 8228 36202 8240
rect 35646 8194 35698 8206
rect 37550 8194 37602 8206
rect 37774 8258 37826 8270
rect 38222 8258 38274 8270
rect 38098 8206 38110 8258
rect 38162 8206 38174 8258
rect 37774 8194 37826 8206
rect 36150 8164 36202 8176
rect 31950 8146 32002 8158
rect 3838 8082 3890 8094
rect 19562 8094 19574 8146
rect 19626 8094 19638 8146
rect 25498 8094 25510 8146
rect 25562 8094 25574 8146
rect 6178 8038 6190 8090
rect 6242 8038 6254 8090
rect 10110 8082 10162 8094
rect 10658 8038 10670 8090
rect 10722 8038 10734 8090
rect 12182 8034 12234 8046
rect 12182 7970 12234 7982
rect 17614 8034 17666 8046
rect 17614 7970 17666 7982
rect 20526 8034 20578 8046
rect 20526 7970 20578 7982
rect 26238 8034 26290 8046
rect 27906 8038 27918 8090
rect 27970 8038 27982 8090
rect 31950 8082 32002 8094
rect 33518 8146 33570 8158
rect 37930 8150 37942 8202
rect 37994 8150 38006 8202
rect 38222 8194 38274 8206
rect 38502 8258 38554 8270
rect 38502 8194 38554 8206
rect 38894 8258 38946 8270
rect 38894 8194 38946 8206
rect 39006 8258 39058 8270
rect 39006 8194 39058 8206
rect 39566 8258 39618 8270
rect 39566 8194 39618 8206
rect 39790 8258 39842 8270
rect 39790 8194 39842 8206
rect 40350 8258 40402 8270
rect 40350 8194 40402 8206
rect 43374 8258 43426 8270
rect 49310 8258 49362 8270
rect 45278 8230 45330 8242
rect 43374 8194 43426 8206
rect 45166 8202 45218 8214
rect 48514 8206 48526 8258
rect 48578 8206 48590 8258
rect 45278 8166 45330 8178
rect 45490 8150 45502 8202
rect 45554 8150 45566 8202
rect 45737 8150 45749 8202
rect 45801 8150 45813 8202
rect 49310 8194 49362 8206
rect 40058 8094 40070 8146
rect 40122 8094 40134 8146
rect 45166 8138 45218 8150
rect 46006 8146 46058 8158
rect 33518 8082 33570 8094
rect 46006 8082 46058 8094
rect 46622 8146 46674 8158
rect 46622 8082 46674 8094
rect 26238 7970 26290 7982
rect 34190 8034 34242 8046
rect 34190 7970 34242 7982
rect 35310 8034 35362 8046
rect 35310 7970 35362 7982
rect 43710 8034 43762 8046
rect 43710 7970 43762 7982
rect 1344 7866 49616 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 49616 7866
rect 1344 7780 49616 7814
rect 5854 7698 5906 7710
rect 5854 7634 5906 7646
rect 7590 7698 7642 7710
rect 7590 7634 7642 7646
rect 48974 7698 49026 7710
rect 8654 7586 8706 7598
rect 10994 7590 11006 7642
rect 11058 7590 11070 7642
rect 7982 7530 8034 7542
rect 1598 7474 1650 7486
rect 7186 7449 7198 7501
rect 7250 7449 7262 7501
rect 7746 7422 7758 7474
rect 7810 7422 7822 7474
rect 7982 7466 8034 7478
rect 8094 7512 8146 7524
rect 8654 7522 8706 7534
rect 11846 7586 11898 7598
rect 11846 7522 11898 7534
rect 12294 7586 12346 7598
rect 12294 7522 12346 7534
rect 20302 7586 20354 7598
rect 8094 7448 8146 7460
rect 1598 7410 1650 7422
rect 8822 7418 8874 7430
rect 9650 7422 9662 7474
rect 9714 7422 9726 7474
rect 9986 7437 9998 7489
rect 10050 7437 10062 7489
rect 10434 7422 10446 7474
rect 10498 7422 10510 7474
rect 10770 7449 10782 7501
rect 10834 7449 10846 7501
rect 11118 7474 11170 7486
rect 11118 7410 11170 7422
rect 12574 7474 12626 7486
rect 13438 7478 13450 7530
rect 13502 7478 13514 7530
rect 20302 7522 20354 7534
rect 24446 7586 24498 7598
rect 24446 7522 24498 7534
rect 29262 7586 29314 7598
rect 31154 7590 31166 7642
rect 31218 7590 31230 7642
rect 48974 7634 49026 7646
rect 29262 7522 29314 7534
rect 38558 7586 38610 7598
rect 38558 7522 38610 7534
rect 45465 7530 45517 7542
rect 44774 7509 44826 7521
rect 12574 7410 12626 7422
rect 14030 7474 14082 7486
rect 17614 7474 17666 7486
rect 14802 7422 14814 7474
rect 14866 7422 14878 7474
rect 18386 7422 18398 7474
rect 18450 7422 18462 7474
rect 20850 7437 20862 7489
rect 20914 7437 20926 7489
rect 21758 7474 21810 7486
rect 21074 7422 21086 7474
rect 21138 7422 21150 7474
rect 14030 7410 14082 7422
rect 17614 7410 17666 7422
rect 21758 7410 21810 7422
rect 25118 7474 25170 7486
rect 27806 7474 27858 7486
rect 25890 7422 25902 7474
rect 25954 7422 25966 7474
rect 25118 7410 25170 7422
rect 27806 7410 27858 7422
rect 28142 7474 28194 7486
rect 28142 7410 28194 7422
rect 28366 7474 28418 7486
rect 28366 7410 28418 7422
rect 28926 7474 28978 7486
rect 28926 7410 28978 7422
rect 30718 7474 30770 7486
rect 31042 7449 31054 7501
rect 31106 7449 31118 7501
rect 32062 7474 32114 7486
rect 31266 7422 31278 7474
rect 31330 7422 31342 7474
rect 31770 7422 31782 7474
rect 31834 7422 31846 7474
rect 30718 7410 30770 7422
rect 32062 7410 32114 7422
rect 32174 7474 32226 7486
rect 32174 7410 32226 7422
rect 34862 7474 34914 7486
rect 34862 7410 34914 7422
rect 34974 7474 35026 7486
rect 34974 7410 35026 7422
rect 35198 7474 35250 7486
rect 35198 7410 35250 7422
rect 35422 7474 35474 7486
rect 37438 7474 37490 7486
rect 35690 7422 35702 7474
rect 35754 7422 35766 7474
rect 36194 7422 36206 7474
rect 36258 7422 36270 7474
rect 36530 7422 36542 7474
rect 36594 7422 36606 7474
rect 38302 7422 38314 7474
rect 38366 7422 38378 7474
rect 39442 7422 39454 7474
rect 39506 7422 39518 7474
rect 41122 7422 41134 7474
rect 41186 7422 41198 7474
rect 43026 7449 43038 7501
rect 43090 7449 43102 7501
rect 43598 7474 43650 7486
rect 44774 7445 44826 7457
rect 45054 7502 45106 7514
rect 45266 7478 45278 7530
rect 45330 7478 45342 7530
rect 45465 7466 45517 7478
rect 45054 7438 45106 7450
rect 45714 7449 45726 7501
rect 45778 7449 45790 7501
rect 48638 7474 48690 7486
rect 35422 7410 35474 7422
rect 37438 7410 37490 7422
rect 43598 7410 43650 7422
rect 48638 7410 48690 7422
rect 2370 7310 2382 7362
rect 2434 7310 2446 7362
rect 4274 7310 4286 7362
rect 4338 7310 4350 7362
rect 8822 7354 8874 7366
rect 33238 7362 33290 7374
rect 10098 7310 10110 7362
rect 10162 7310 10174 7362
rect 16706 7310 16718 7362
rect 16770 7310 16782 7362
rect 20738 7310 20750 7362
rect 20802 7310 20814 7362
rect 22530 7310 22542 7362
rect 22594 7310 22606 7362
rect 33238 7298 33290 7310
rect 33686 7362 33738 7374
rect 33686 7298 33738 7310
rect 34246 7362 34298 7374
rect 37046 7362 37098 7374
rect 34246 7298 34298 7310
rect 36094 7306 36146 7318
rect 13694 7250 13746 7262
rect 37046 7298 37098 7310
rect 39174 7362 39226 7374
rect 39174 7298 39226 7310
rect 28634 7198 28646 7250
rect 28698 7198 28710 7250
rect 34570 7198 34582 7250
rect 34634 7198 34646 7250
rect 36094 7242 36146 7254
rect 43934 7250 43986 7262
rect 13694 7186 13746 7198
rect 43934 7186 43986 7198
rect 44550 7250 44602 7262
rect 44550 7186 44602 7198
rect 47070 7250 47122 7262
rect 47070 7186 47122 7198
rect 1344 7082 49616 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 49616 7082
rect 1344 6996 49616 7030
rect 2494 6914 2546 6926
rect 2494 6850 2546 6862
rect 23102 6914 23154 6926
rect 23102 6850 23154 6862
rect 37158 6914 37210 6926
rect 37930 6862 37942 6914
rect 37994 6862 38006 6914
rect 37158 6850 37210 6862
rect 7758 6802 7810 6814
rect 5058 6750 5070 6802
rect 5122 6750 5134 6802
rect 9762 6750 9774 6802
rect 9826 6750 9838 6802
rect 12226 6750 12238 6802
rect 12290 6750 12302 6802
rect 14130 6750 14142 6802
rect 14194 6750 14206 6802
rect 25442 6750 25454 6802
rect 25506 6750 25518 6802
rect 27458 6750 27470 6802
rect 27522 6750 27534 6802
rect 30258 6750 30270 6802
rect 30322 6750 30334 6802
rect 33170 6750 33182 6802
rect 33234 6750 33246 6802
rect 40450 6750 40462 6802
rect 40514 6750 40526 6802
rect 7758 6738 7810 6750
rect 2830 6690 2882 6702
rect 6302 6690 6354 6702
rect 8094 6690 8146 6702
rect 3714 6638 3726 6690
rect 3778 6638 3790 6690
rect 4610 6638 4622 6690
rect 4674 6638 4686 6690
rect 2830 6626 2882 6638
rect 4946 6623 4958 6675
rect 5010 6623 5022 6675
rect 5618 6638 5630 6690
rect 5682 6638 5694 6690
rect 7074 6638 7086 6690
rect 7138 6638 7150 6690
rect 7410 6638 7422 6690
rect 7474 6638 7486 6690
rect 13022 6690 13074 6702
rect 5954 6582 5966 6634
rect 6018 6582 6030 6634
rect 6302 6626 6354 6638
rect 7746 6582 7758 6634
rect 7810 6582 7822 6634
rect 8094 6626 8146 6638
rect 8642 6605 8654 6657
rect 8706 6605 8718 6657
rect 8978 6582 8990 6634
rect 9042 6582 9054 6634
rect 9426 6582 9438 6634
rect 9490 6582 9502 6634
rect 9736 6598 9748 6650
rect 9800 6598 9812 6650
rect 13022 6626 13074 6638
rect 13358 6690 13410 6702
rect 17166 6690 17218 6702
rect 16594 6638 16606 6690
rect 16658 6638 16670 6690
rect 13358 6626 13410 6638
rect 10334 6578 10386 6590
rect 6918 6522 6970 6534
rect 5730 6470 5742 6522
rect 5794 6470 5806 6522
rect 10334 6514 10386 6526
rect 16046 6578 16098 6590
rect 16930 6582 16942 6634
rect 16994 6582 17006 6634
rect 17166 6626 17218 6638
rect 17614 6690 17666 6702
rect 17614 6626 17666 6638
rect 17838 6690 17890 6702
rect 19630 6690 19682 6702
rect 18386 6638 18398 6690
rect 18450 6638 18462 6690
rect 19058 6638 19070 6690
rect 19122 6638 19134 6690
rect 19406 6651 19458 6663
rect 17838 6626 17890 6638
rect 19630 6626 19682 6638
rect 20078 6690 20130 6702
rect 20078 6626 20130 6638
rect 20302 6690 20354 6702
rect 20302 6626 20354 6638
rect 21198 6690 21250 6702
rect 21198 6626 21250 6638
rect 22430 6690 22482 6702
rect 22430 6626 22482 6638
rect 23438 6690 23490 6702
rect 23438 6626 23490 6638
rect 23998 6690 24050 6702
rect 25958 6690 26010 6702
rect 23998 6626 24050 6638
rect 24322 6611 24334 6663
rect 24386 6611 24398 6663
rect 24546 6638 24558 6690
rect 24610 6638 24622 6690
rect 24994 6638 25006 6690
rect 25058 6638 25070 6690
rect 25330 6623 25342 6675
rect 25394 6623 25406 6675
rect 25958 6626 26010 6638
rect 26462 6690 26514 6702
rect 29598 6690 29650 6702
rect 30494 6690 30546 6702
rect 26462 6626 26514 6638
rect 26786 6611 26798 6663
rect 26850 6611 26862 6663
rect 27122 6638 27134 6690
rect 27186 6638 27198 6690
rect 27570 6623 27582 6675
rect 27634 6623 27646 6675
rect 27906 6638 27918 6690
rect 27970 6638 27982 6690
rect 29922 6638 29934 6690
rect 29986 6638 29998 6690
rect 29598 6626 29650 6638
rect 19406 6587 19458 6599
rect 30146 6594 30158 6646
rect 30210 6594 30222 6646
rect 30494 6626 30546 6638
rect 30718 6690 30770 6702
rect 30718 6626 30770 6638
rect 31838 6690 31890 6702
rect 32622 6690 32674 6702
rect 32330 6638 32342 6690
rect 32394 6638 32406 6690
rect 31838 6626 31890 6638
rect 32622 6626 32674 6638
rect 32846 6690 32898 6702
rect 35870 6690 35922 6702
rect 35074 6638 35086 6690
rect 35138 6638 35150 6690
rect 32846 6626 32898 6638
rect 35870 6626 35922 6638
rect 36542 6690 36594 6702
rect 37550 6690 37602 6702
rect 37314 6638 37326 6690
rect 37378 6638 37390 6690
rect 36542 6626 36594 6638
rect 37550 6626 37602 6638
rect 37662 6690 37714 6702
rect 37662 6626 37714 6638
rect 38558 6690 38610 6702
rect 38558 6626 38610 6638
rect 41246 6690 41298 6702
rect 41246 6626 41298 6638
rect 41358 6690 41410 6702
rect 41358 6626 41410 6638
rect 41694 6690 41746 6702
rect 41694 6626 41746 6638
rect 42590 6690 42642 6702
rect 49310 6690 49362 6702
rect 42590 6626 42642 6638
rect 43150 6662 43202 6674
rect 45558 6655 45610 6667
rect 43710 6634 43762 6646
rect 43150 6598 43202 6610
rect 42870 6578 42922 6590
rect 43362 6582 43374 6634
rect 43426 6582 43438 6634
rect 43586 6582 43598 6634
rect 43650 6582 43662 6634
rect 45110 6634 45162 6646
rect 18106 6526 18118 6578
rect 18170 6526 18182 6578
rect 16046 6514 16098 6526
rect 18566 6522 18618 6534
rect 20570 6526 20582 6578
rect 20634 6526 20646 6578
rect 30986 6526 30998 6578
rect 31050 6526 31062 6578
rect 43710 6570 43762 6582
rect 44886 6578 44938 6590
rect 17266 6470 17278 6522
rect 17330 6470 17342 6522
rect 19506 6470 19518 6522
rect 19570 6470 19582 6522
rect 6918 6458 6970 6470
rect 18566 6458 18618 6470
rect 21534 6466 21586 6478
rect 21534 6402 21586 6414
rect 22094 6466 22146 6478
rect 23874 6470 23886 6522
rect 23938 6470 23950 6522
rect 26338 6470 26350 6522
rect 26402 6470 26414 6522
rect 42870 6514 42922 6526
rect 45378 6582 45390 6634
rect 45442 6582 45454 6634
rect 45558 6591 45610 6603
rect 45726 6634 45778 6646
rect 48514 6638 48526 6690
rect 48578 6638 48590 6690
rect 49310 6626 49362 6638
rect 45110 6570 45162 6582
rect 45726 6570 45778 6582
rect 46622 6578 46674 6590
rect 44886 6514 44938 6526
rect 46622 6514 46674 6526
rect 22094 6402 22146 6414
rect 29262 6466 29314 6478
rect 29262 6402 29314 6414
rect 31502 6466 31554 6478
rect 31502 6402 31554 6414
rect 36206 6466 36258 6478
rect 36206 6402 36258 6414
rect 42254 6466 42306 6478
rect 42254 6402 42306 6414
rect 44214 6466 44266 6478
rect 44214 6402 44266 6414
rect 46118 6466 46170 6478
rect 46118 6402 46170 6414
rect 1344 6298 49616 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 49616 6298
rect 1344 6212 49616 6246
rect 11454 6130 11506 6142
rect 5058 6022 5070 6074
rect 5122 6022 5134 6074
rect 11454 6066 11506 6078
rect 18342 6130 18394 6142
rect 18342 6066 18394 6078
rect 18734 6130 18786 6142
rect 18734 6066 18786 6078
rect 25398 6130 25450 6142
rect 25398 6066 25450 6078
rect 25846 6130 25898 6142
rect 25846 6066 25898 6078
rect 26518 6130 26570 6142
rect 26518 6066 26570 6078
rect 8430 6018 8482 6030
rect 6570 5966 6582 6018
rect 6634 5966 6646 6018
rect 4734 5906 4786 5918
rect 5226 5910 5238 5962
rect 5290 5910 5302 5962
rect 5630 5906 5682 5918
rect 4946 5854 4958 5906
rect 5010 5854 5022 5906
rect 4734 5842 4786 5854
rect 5630 5842 5682 5854
rect 6078 5906 6130 5918
rect 6078 5842 6130 5854
rect 6302 5906 6354 5918
rect 6302 5842 6354 5854
rect 6974 5906 7026 5918
rect 7422 5906 7474 5918
rect 6974 5842 7026 5854
rect 7142 5850 7194 5862
rect 7298 5854 7310 5906
rect 7362 5854 7374 5906
rect 7422 5842 7474 5854
rect 8094 5906 8146 5918
rect 8250 5910 8262 5962
rect 8314 5910 8326 5962
rect 8430 5954 8482 5966
rect 8822 6018 8874 6030
rect 8822 5954 8874 5966
rect 29822 6018 29874 6030
rect 30370 6022 30382 6074
rect 30434 6022 30446 6074
rect 31714 6022 31726 6074
rect 31778 6022 31790 6074
rect 39118 6018 39170 6030
rect 8094 5842 8146 5854
rect 8542 5906 8594 5918
rect 11118 5906 11170 5918
rect 9986 5854 9998 5906
rect 10050 5854 10062 5906
rect 10322 5854 10334 5906
rect 10386 5854 10398 5906
rect 8542 5842 8594 5854
rect 11118 5842 11170 5854
rect 15374 5906 15426 5918
rect 15698 5854 15710 5906
rect 15762 5854 15774 5906
rect 15922 5869 15934 5921
rect 15986 5869 15998 5921
rect 16382 5906 16434 5918
rect 15374 5842 15426 5854
rect 16382 5842 16434 5854
rect 16494 5906 16546 5918
rect 17490 5869 17502 5921
rect 17554 5869 17566 5921
rect 19070 5906 19122 5918
rect 17714 5854 17726 5906
rect 17778 5854 17790 5906
rect 19282 5881 19294 5933
rect 19346 5881 19358 5933
rect 22188 5906 22240 5918
rect 16494 5842 16546 5854
rect 19070 5842 19122 5854
rect 22188 5842 22240 5854
rect 22430 5906 22482 5918
rect 22922 5910 22934 5962
rect 22986 5910 22998 5962
rect 29822 5954 29874 5966
rect 38558 5962 38610 5974
rect 22430 5842 22482 5854
rect 23102 5906 23154 5918
rect 23102 5842 23154 5854
rect 24446 5906 24498 5918
rect 24446 5842 24498 5854
rect 24558 5906 24610 5918
rect 24558 5842 24610 5854
rect 27134 5906 27186 5918
rect 30538 5910 30550 5962
rect 30602 5910 30614 5962
rect 32062 5945 32114 5957
rect 30942 5906 30994 5918
rect 27906 5854 27918 5906
rect 27970 5854 27982 5906
rect 30258 5854 30270 5906
rect 30322 5854 30334 5906
rect 31602 5854 31614 5906
rect 31666 5854 31678 5906
rect 32062 5881 32114 5893
rect 32286 5906 32338 5918
rect 33406 5906 33458 5918
rect 33114 5854 33126 5906
rect 33178 5854 33190 5906
rect 27134 5842 27186 5854
rect 30942 5842 30994 5854
rect 32286 5842 32338 5854
rect 33406 5842 33458 5854
rect 33518 5906 33570 5918
rect 33842 5854 33854 5906
rect 33906 5854 33918 5906
rect 34178 5869 34190 5921
rect 34242 5869 34254 5921
rect 34738 5854 34750 5906
rect 34802 5854 34814 5906
rect 34962 5898 34974 5950
rect 35026 5898 35038 5950
rect 35634 5854 35646 5906
rect 35698 5854 35710 5906
rect 37874 5881 37886 5933
rect 37938 5881 37950 5933
rect 39118 5954 39170 5966
rect 43598 6018 43650 6030
rect 43598 5954 43650 5966
rect 44102 6018 44154 6030
rect 44102 5954 44154 5966
rect 38558 5898 38610 5910
rect 40910 5906 40962 5918
rect 44370 5910 44382 5962
rect 44434 5910 44446 5962
rect 44594 5910 44606 5962
rect 44658 5910 44670 5962
rect 44830 5934 44882 5946
rect 38882 5854 38894 5906
rect 38946 5854 38958 5906
rect 33518 5842 33570 5854
rect 39286 5850 39338 5862
rect 39666 5854 39678 5906
rect 39730 5854 39742 5906
rect 39890 5854 39902 5906
rect 39954 5854 39966 5906
rect 44830 5870 44882 5882
rect 44942 5941 44994 5953
rect 48302 5906 48354 5918
rect 44942 5877 44994 5889
rect 47506 5854 47518 5906
rect 47570 5854 47582 5906
rect 48626 5854 48638 5906
rect 48690 5854 48702 5906
rect 7142 5786 7194 5798
rect 23606 5794 23658 5806
rect 40910 5842 40962 5854
rect 48302 5842 48354 5854
rect 16034 5742 16046 5794
rect 16098 5742 16110 5794
rect 17378 5742 17390 5794
rect 17442 5742 17454 5794
rect 34290 5742 34302 5794
rect 34354 5742 34366 5794
rect 35074 5742 35086 5794
rect 35138 5742 35150 5794
rect 39286 5786 39338 5798
rect 4398 5682 4450 5694
rect 4398 5618 4450 5630
rect 7702 5682 7754 5694
rect 10098 5686 10110 5738
rect 10162 5686 10174 5738
rect 23606 5730 23658 5742
rect 39566 5738 39618 5750
rect 41682 5742 41694 5794
rect 41746 5742 41758 5794
rect 45602 5742 45614 5794
rect 45666 5742 45678 5794
rect 7702 5618 7754 5630
rect 15038 5682 15090 5694
rect 20302 5682 20354 5694
rect 16762 5630 16774 5682
rect 16826 5630 16838 5682
rect 24154 5630 24166 5682
rect 24218 5630 24230 5682
rect 39566 5674 39618 5686
rect 15038 5618 15090 5630
rect 20302 5618 20354 5630
rect 1344 5514 49616 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 49616 5514
rect 1344 5428 49616 5462
rect 6190 5346 6242 5358
rect 6190 5282 6242 5294
rect 6862 5346 6914 5358
rect 10334 5346 10386 5358
rect 9706 5294 9718 5346
rect 9770 5294 9782 5346
rect 6862 5282 6914 5294
rect 10334 5282 10386 5294
rect 29318 5234 29370 5246
rect 37158 5234 37210 5246
rect 3042 5182 3054 5234
rect 3106 5182 3118 5234
rect 4946 5182 4958 5234
rect 5010 5182 5022 5234
rect 7970 5182 7982 5234
rect 8034 5182 8046 5234
rect 8306 5182 8318 5234
rect 8370 5182 8382 5234
rect 14802 5182 14814 5234
rect 14866 5182 14878 5234
rect 16706 5182 16718 5234
rect 16770 5182 16782 5234
rect 18498 5182 18510 5234
rect 18562 5182 18574 5234
rect 20738 5182 20750 5234
rect 20802 5182 20814 5234
rect 22934 5178 22986 5190
rect 2270 5122 2322 5134
rect 2270 5058 2322 5070
rect 5854 5122 5906 5134
rect 5854 5058 5906 5070
rect 6526 5122 6578 5134
rect 9214 5122 9266 5134
rect 7522 5070 7534 5122
rect 7586 5070 7598 5122
rect 6526 5058 6578 5070
rect 7858 5055 7870 5107
rect 7922 5055 7934 5107
rect 8418 5055 8430 5107
rect 8482 5055 8494 5107
rect 8642 5070 8654 5122
rect 8706 5070 8718 5122
rect 9214 5058 9266 5070
rect 9438 5122 9490 5134
rect 9438 5058 9490 5070
rect 9998 5122 10050 5134
rect 9998 5058 10050 5070
rect 14030 5122 14082 5134
rect 21198 5122 21250 5134
rect 14030 5058 14082 5070
rect 17490 5042 17502 5094
rect 17554 5042 17566 5094
rect 20290 5070 20302 5122
rect 20354 5070 20366 5122
rect 20626 5055 20638 5107
rect 20690 5055 20702 5107
rect 21198 5058 21250 5070
rect 22430 5122 22482 5134
rect 33170 5182 33182 5234
rect 33234 5182 33246 5234
rect 36306 5182 36318 5234
rect 36370 5182 36382 5234
rect 39330 5182 39342 5234
rect 39394 5182 39406 5234
rect 44930 5182 44942 5234
rect 44994 5182 45006 5234
rect 29318 5170 29370 5182
rect 37158 5170 37210 5182
rect 22934 5114 22986 5126
rect 23102 5122 23154 5134
rect 22430 5058 22482 5070
rect 23102 5058 23154 5070
rect 23662 5122 23714 5134
rect 26350 5122 26402 5134
rect 25554 5070 25566 5122
rect 25618 5070 25630 5122
rect 23662 5058 23714 5070
rect 26350 5058 26402 5070
rect 27022 5122 27074 5134
rect 27022 5058 27074 5070
rect 27918 5122 27970 5134
rect 28478 5122 28530 5134
rect 28186 5070 28198 5122
rect 28250 5070 28262 5122
rect 27918 5058 27970 5070
rect 28478 5058 28530 5070
rect 28702 5122 28754 5134
rect 28702 5058 28754 5070
rect 29486 5122 29538 5134
rect 29486 5058 29538 5070
rect 30494 5122 30546 5134
rect 33630 5122 33682 5134
rect 38110 5122 38162 5134
rect 31266 5070 31278 5122
rect 31330 5070 31342 5122
rect 34402 5070 34414 5122
rect 34466 5070 34478 5122
rect 37426 5070 37438 5122
rect 37490 5070 37502 5122
rect 30494 5058 30546 5070
rect 33630 5058 33682 5070
rect 22188 5010 22240 5022
rect 37874 5014 37886 5066
rect 37938 5014 37950 5066
rect 38110 5058 38162 5070
rect 38558 5122 38610 5134
rect 38558 5058 38610 5070
rect 41246 5122 41298 5134
rect 47630 5122 47682 5134
rect 41246 5058 41298 5070
rect 41682 5042 41694 5094
rect 41746 5042 41758 5094
rect 46834 5070 46846 5122
rect 46898 5070 46910 5122
rect 47630 5058 47682 5070
rect 47854 5087 47906 5099
rect 47854 5023 47906 5035
rect 47966 5094 48018 5106
rect 47966 5030 48018 5042
rect 48190 5094 48242 5106
rect 48190 5030 48242 5042
rect 48414 5094 48466 5106
rect 48414 5030 48466 5042
rect 22188 4946 22240 4958
rect 48694 5010 48746 5022
rect 21534 4898 21586 4910
rect 21534 4834 21586 4846
rect 26686 4898 26738 4910
rect 26686 4834 26738 4846
rect 27582 4898 27634 4910
rect 38210 4902 38222 4954
rect 38274 4902 38286 4954
rect 48694 4946 48746 4958
rect 27582 4834 27634 4846
rect 43038 4898 43090 4910
rect 43038 4834 43090 4846
rect 49142 4898 49194 4910
rect 49142 4834 49194 4846
rect 1344 4730 49616 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 49616 4730
rect 1344 4644 49616 4678
rect 15374 4562 15426 4574
rect 15374 4498 15426 4510
rect 24558 4562 24610 4574
rect 31166 4562 31218 4574
rect 8878 4450 8930 4462
rect 16034 4454 16046 4506
rect 16098 4454 16110 4506
rect 18498 4454 18510 4506
rect 18562 4454 18574 4506
rect 24558 4498 24610 4510
rect 26630 4506 26682 4518
rect 8878 4386 8930 4398
rect 22318 4450 22370 4462
rect 6190 4338 6242 4350
rect 14366 4338 14418 4350
rect 6962 4286 6974 4338
rect 7026 4286 7038 4338
rect 6190 4274 6242 4286
rect 14366 4274 14418 4286
rect 15038 4338 15090 4350
rect 15038 4274 15090 4286
rect 15710 4338 15762 4350
rect 16202 4342 16214 4394
rect 16266 4342 16278 4394
rect 16606 4338 16658 4350
rect 16034 4286 16046 4338
rect 16098 4286 16110 4338
rect 15710 4274 15762 4286
rect 16606 4274 16658 4286
rect 17726 4338 17778 4350
rect 17726 4274 17778 4286
rect 17950 4338 18002 4350
rect 17950 4274 18002 4286
rect 18398 4338 18450 4350
rect 18722 4342 18734 4394
rect 18786 4342 18798 4394
rect 22318 4386 22370 4398
rect 22860 4450 22912 4462
rect 22860 4386 22912 4398
rect 23774 4450 23826 4462
rect 19630 4338 19682 4350
rect 23102 4338 23154 4350
rect 23594 4342 23606 4394
rect 23658 4342 23670 4394
rect 23774 4386 23826 4398
rect 25230 4450 25282 4462
rect 25230 4386 25282 4398
rect 26144 4450 26196 4462
rect 47742 4562 47794 4574
rect 31166 4498 31218 4510
rect 40966 4506 41018 4518
rect 26630 4442 26682 4454
rect 29598 4450 29650 4462
rect 18946 4286 18958 4338
rect 19010 4286 19022 4338
rect 20402 4286 20414 4338
rect 20466 4286 20478 4338
rect 18398 4274 18450 4286
rect 19630 4274 19682 4286
rect 23102 4274 23154 4286
rect 24222 4338 24274 4350
rect 25386 4342 25398 4394
rect 25450 4342 25462 4394
rect 26144 4386 26196 4398
rect 29598 4386 29650 4398
rect 38670 4450 38722 4462
rect 47742 4498 47794 4510
rect 48974 4562 49026 4574
rect 48974 4498 49026 4510
rect 40966 4442 41018 4454
rect 44046 4450 44098 4462
rect 38670 4386 38722 4398
rect 44046 4386 44098 4398
rect 44606 4450 44658 4462
rect 44606 4386 44658 4398
rect 24222 4274 24274 4286
rect 25902 4338 25954 4350
rect 25902 4274 25954 4286
rect 26910 4338 26962 4350
rect 27682 4286 27694 4338
rect 27746 4286 27758 4338
rect 32498 4313 32510 4365
rect 32562 4313 32574 4365
rect 33182 4338 33234 4350
rect 35870 4338 35922 4350
rect 35074 4286 35086 4338
rect 35138 4286 35150 4338
rect 26910 4274 26962 4286
rect 33182 4274 33234 4286
rect 35870 4274 35922 4286
rect 35982 4338 36034 4350
rect 36754 4286 36766 4338
rect 36818 4286 36830 4338
rect 39218 4330 39230 4382
rect 39282 4330 39294 4382
rect 39790 4338 39842 4350
rect 39442 4286 39454 4338
rect 39506 4286 39518 4338
rect 35982 4274 36034 4286
rect 39790 4274 39842 4286
rect 40126 4338 40178 4350
rect 40126 4274 40178 4286
rect 41358 4338 41410 4350
rect 47294 4338 47346 4350
rect 42130 4286 42142 4338
rect 42194 4286 42206 4338
rect 41358 4274 41410 4286
rect 47294 4274 47346 4286
rect 47406 4338 47458 4350
rect 47406 4274 47458 4286
rect 48638 4338 48690 4350
rect 48638 4274 48690 4286
rect 17434 4174 17446 4226
rect 17498 4174 17510 4226
rect 39106 4174 39118 4226
rect 39170 4174 39182 4226
rect 46498 4174 46510 4226
rect 46562 4174 46574 4226
rect 14030 4114 14082 4126
rect 14030 4050 14082 4062
rect 14702 4114 14754 4126
rect 14702 4050 14754 4062
rect 1344 3946 49616 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 49616 3946
rect 1344 3860 49616 3894
rect 31054 3778 31106 3790
rect 42702 3778 42754 3790
rect 31054 3714 31106 3726
rect 34974 3722 35026 3734
rect 38826 3726 38838 3778
rect 38890 3726 38902 3778
rect 42702 3714 42754 3726
rect 48302 3778 48354 3790
rect 48302 3714 48354 3726
rect 48974 3778 49026 3790
rect 48974 3714 49026 3726
rect 17714 3614 17726 3666
rect 17778 3614 17790 3666
rect 19618 3614 19630 3666
rect 19682 3614 19694 3666
rect 22082 3614 22094 3666
rect 22146 3614 22158 3666
rect 24770 3614 24782 3666
rect 24834 3614 24846 3666
rect 26674 3614 26686 3666
rect 26738 3614 26750 3666
rect 30594 3614 30606 3666
rect 30658 3614 30670 3666
rect 34974 3658 35026 3670
rect 47630 3666 47682 3678
rect 36978 3614 36990 3666
rect 37042 3614 37054 3666
rect 47630 3602 47682 3614
rect 16942 3554 16994 3566
rect 14018 3474 14030 3526
rect 14082 3474 14094 3526
rect 27470 3554 27522 3566
rect 16942 3490 16994 3502
rect 21410 3474 21422 3526
rect 21474 3474 21486 3526
rect 27470 3490 27522 3502
rect 29150 3554 29202 3566
rect 31390 3554 31442 3566
rect 39118 3554 39170 3566
rect 29150 3490 29202 3502
rect 29474 3475 29486 3527
rect 29538 3475 29550 3527
rect 29698 3502 29710 3554
rect 29762 3502 29774 3554
rect 30146 3502 30158 3554
rect 30210 3502 30222 3554
rect 30482 3487 30494 3539
rect 30546 3487 30558 3539
rect 32386 3502 32398 3554
rect 32450 3502 32462 3554
rect 31390 3490 31442 3502
rect 34626 3474 34638 3526
rect 34690 3474 34702 3526
rect 35074 3502 35086 3554
rect 35138 3502 35150 3554
rect 35410 3502 35422 3554
rect 35474 3502 35486 3554
rect 36194 3474 36206 3526
rect 36258 3474 36270 3526
rect 39118 3490 39170 3502
rect 39342 3554 39394 3566
rect 43038 3554 43090 3566
rect 39342 3490 39394 3502
rect 42018 3474 42030 3526
rect 42082 3474 42094 3526
rect 43038 3490 43090 3502
rect 43766 3554 43818 3566
rect 46958 3554 47010 3566
rect 43766 3490 43818 3502
rect 44046 3526 44098 3538
rect 44494 3526 44546 3538
rect 44046 3462 44098 3474
rect 44258 3446 44270 3498
rect 44322 3446 44334 3498
rect 44494 3462 44546 3474
rect 44606 3519 44658 3531
rect 44606 3455 44658 3467
rect 45558 3519 45610 3531
rect 45558 3455 45610 3467
rect 45838 3526 45890 3538
rect 45838 3462 45890 3474
rect 45334 3442 45386 3454
rect 46050 3446 46062 3498
rect 46114 3446 46126 3498
rect 46218 3486 46230 3538
rect 46282 3486 46294 3538
rect 46958 3490 47010 3502
rect 47294 3554 47346 3566
rect 47294 3490 47346 3502
rect 47966 3554 48018 3566
rect 47966 3490 48018 3502
rect 48638 3554 48690 3566
rect 48638 3490 48690 3502
rect 5574 3386 5626 3398
rect 1766 3330 1818 3342
rect 1766 3266 1818 3278
rect 3222 3330 3274 3342
rect 20134 3386 20186 3398
rect 5574 3322 5626 3334
rect 6806 3330 6858 3342
rect 3222 3266 3274 3278
rect 6806 3266 6858 3278
rect 8598 3330 8650 3342
rect 8598 3266 8650 3278
rect 10390 3330 10442 3342
rect 10390 3266 10442 3278
rect 12182 3330 12234 3342
rect 12182 3266 12234 3278
rect 13526 3330 13578 3342
rect 13526 3266 13578 3278
rect 15598 3330 15650 3342
rect 27750 3386 27802 3398
rect 40562 3390 40574 3442
rect 40626 3390 40638 3442
rect 20134 3322 20186 3334
rect 23942 3330 23994 3342
rect 15598 3266 15650 3278
rect 27750 3322 27802 3334
rect 28422 3330 28474 3342
rect 29026 3334 29038 3386
rect 29090 3334 29102 3386
rect 45334 3378 45386 3390
rect 23942 3266 23994 3278
rect 28422 3266 28474 3278
rect 46622 3330 46674 3342
rect 46622 3266 46674 3278
rect 1344 3162 49616 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 49616 3162
rect 1344 3076 49616 3110
rect 23930 2718 23942 2770
rect 23994 2767 24006 2770
rect 24434 2767 24446 2770
rect 23994 2721 24446 2767
rect 23994 2718 24006 2721
rect 24434 2718 24446 2721
rect 24498 2718 24510 2770
<< via1 >>
rect 30662 47966 30714 48018
rect 31838 47966 31890 48018
rect 43374 47966 43426 48018
rect 43822 47966 43874 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 14366 47630 14418 47682
rect 14814 47518 14866 47570
rect 19014 47518 19066 47570
rect 22430 47518 22482 47570
rect 30662 47518 30714 47570
rect 32622 47518 32674 47570
rect 35982 47518 36034 47570
rect 38838 47518 38890 47570
rect 39286 47518 39338 47570
rect 46398 47518 46450 47570
rect 11790 47406 11842 47458
rect 13246 47406 13298 47458
rect 14122 47350 14174 47402
rect 14926 47391 14978 47443
rect 15150 47406 15202 47458
rect 19182 47406 19234 47458
rect 21198 47406 21250 47458
rect 22766 47406 22818 47458
rect 23102 47406 23154 47458
rect 22598 47350 22650 47402
rect 24670 47362 24722 47414
rect 24894 47406 24946 47458
rect 26238 47406 26290 47458
rect 26350 47406 26402 47458
rect 26630 47406 26682 47458
rect 28366 47406 28418 47458
rect 29242 47406 29294 47458
rect 30830 47406 30882 47458
rect 32174 47406 32226 47458
rect 32510 47362 32562 47414
rect 35198 47378 35250 47430
rect 36094 47362 36146 47414
rect 36318 47406 36370 47458
rect 37326 47406 37378 47458
rect 38278 47406 38330 47458
rect 39678 47406 39730 47458
rect 40462 47406 40514 47458
rect 42814 47406 42866 47458
rect 43822 47406 43874 47458
rect 45838 47378 45890 47430
rect 46510 47362 46562 47414
rect 46734 47406 46786 47458
rect 47294 47406 47346 47458
rect 47966 47406 48018 47458
rect 49310 47406 49362 47458
rect 29486 47294 29538 47346
rect 11454 47182 11506 47234
rect 19518 47182 19570 47234
rect 20918 47182 20970 47234
rect 21366 47182 21418 47234
rect 21926 47182 21978 47234
rect 24782 47238 24834 47290
rect 42366 47294 42418 47346
rect 23270 47182 23322 47234
rect 30214 47182 30266 47234
rect 31166 47182 31218 47234
rect 33742 47182 33794 47234
rect 36934 47182 36986 47234
rect 37662 47182 37714 47234
rect 42982 47238 43034 47290
rect 47630 47182 47682 47234
rect 48134 47182 48186 47234
rect 48974 47182 49026 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 22878 46734 22930 46786
rect 23438 46734 23490 46786
rect 25342 46734 25394 46786
rect 40238 46790 40290 46842
rect 10222 46622 10274 46674
rect 11006 46622 11058 46674
rect 13358 46622 13410 46674
rect 13470 46622 13522 46674
rect 14030 46622 14082 46674
rect 14814 46622 14866 46674
rect 17614 46622 17666 46674
rect 19966 46622 20018 46674
rect 20190 46622 20242 46674
rect 20974 46622 21026 46674
rect 23681 46622 23733 46674
rect 24558 46622 24610 46674
rect 25585 46653 25637 46705
rect 26462 46622 26514 46674
rect 27582 46622 27634 46674
rect 30270 46622 30322 46674
rect 30382 46622 30434 46674
rect 30606 46622 30658 46674
rect 31446 46651 31498 46703
rect 31726 46622 31778 46674
rect 32062 46622 32114 46674
rect 32958 46622 33010 46674
rect 35534 46622 35586 46674
rect 36318 46622 36370 46674
rect 39342 46622 39394 46674
rect 40014 46622 40066 46674
rect 40238 46637 40290 46689
rect 41750 46678 41802 46730
rect 41470 46622 41522 46674
rect 41582 46622 41634 46674
rect 41918 46622 41970 46674
rect 44494 46622 44546 46674
rect 45278 46622 45330 46674
rect 45390 46622 45442 46674
rect 48638 46622 48690 46674
rect 12910 46510 12962 46562
rect 16718 46510 16770 46562
rect 29486 46510 29538 46562
rect 31278 46510 31330 46562
rect 33630 46510 33682 46562
rect 36654 46510 36706 46562
rect 38558 46510 38610 46562
rect 42590 46510 42642 46562
rect 46174 46510 46226 46562
rect 48078 46510 48130 46562
rect 48974 46510 49026 46562
rect 13750 46398 13802 46450
rect 17446 46398 17498 46450
rect 19630 46398 19682 46450
rect 30886 46398 30938 46450
rect 32398 46398 32450 46450
rect 33126 46398 33178 46450
rect 41190 46398 41242 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 40350 46006 40402 46058
rect 43822 46062 43874 46114
rect 11454 45950 11506 46002
rect 18734 45950 18786 46002
rect 22654 45950 22706 46002
rect 24446 45950 24498 46002
rect 29598 45950 29650 46002
rect 30830 45950 30882 46002
rect 37662 45950 37714 46002
rect 41358 45950 41410 46002
rect 9550 45838 9602 45890
rect 11118 45838 11170 45890
rect 11342 45794 11394 45846
rect 12014 45838 12066 45890
rect 12350 45811 12402 45863
rect 12574 45838 12626 45890
rect 14702 45838 14754 45890
rect 13825 45782 13877 45834
rect 14926 45838 14978 45890
rect 15710 45838 15762 45890
rect 17950 45838 18002 45890
rect 21310 45838 21362 45890
rect 22766 45794 22818 45846
rect 23102 45838 23154 45890
rect 23662 45838 23714 45890
rect 26350 45838 26402 45890
rect 27694 45838 27746 45890
rect 27806 45838 27858 45890
rect 28646 45838 28698 45890
rect 29150 45838 29202 45890
rect 29430 45808 29482 45860
rect 30046 45838 30098 45890
rect 33518 45810 33570 45862
rect 36878 45838 36930 45890
rect 40462 45838 40514 45890
rect 40798 45838 40850 45890
rect 41246 45838 41298 45890
rect 41470 45811 41522 45863
rect 41806 45838 41858 45890
rect 42142 45838 42194 45890
rect 42702 45838 42754 45890
rect 45054 45838 45106 45890
rect 45278 45838 45330 45890
rect 45950 45838 46002 45890
rect 13582 45726 13634 45778
rect 12126 45670 12178 45722
rect 17614 45726 17666 45778
rect 20638 45726 20690 45778
rect 32734 45726 32786 45778
rect 43578 45782 43630 45834
rect 45614 45782 45666 45834
rect 46398 45838 46450 45890
rect 47182 45838 47234 45890
rect 39566 45726 39618 45778
rect 49086 45726 49138 45778
rect 27358 45614 27410 45666
rect 27974 45614 28026 45666
rect 36486 45614 36538 45666
rect 46062 45670 46114 45722
rect 44886 45614 44938 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 38894 45278 38946 45330
rect 30718 45222 30770 45274
rect 39958 45278 40010 45330
rect 40406 45278 40458 45330
rect 12126 45166 12178 45218
rect 47518 45222 47570 45274
rect 37494 45166 37546 45218
rect 9438 45054 9490 45106
rect 13470 45054 13522 45106
rect 13694 45093 13746 45145
rect 14030 45054 14082 45106
rect 14590 45098 14642 45150
rect 14814 45054 14866 45106
rect 15374 45054 15426 45106
rect 15598 45098 15650 45150
rect 16942 45054 16994 45106
rect 17726 45054 17778 45106
rect 17838 45054 17890 45106
rect 18398 45054 18450 45106
rect 21534 45054 21586 45106
rect 22318 45054 22370 45106
rect 25230 45054 25282 45106
rect 25566 45069 25618 45121
rect 25902 45054 25954 45106
rect 26686 45054 26738 45106
rect 30606 45054 30658 45106
rect 31054 45093 31106 45145
rect 31278 45054 31330 45106
rect 31726 45054 31778 45106
rect 31950 45054 32002 45106
rect 32230 45054 32282 45106
rect 32958 45054 33010 45106
rect 33742 45054 33794 45106
rect 36206 45089 36258 45141
rect 36318 45110 36370 45162
rect 36542 45082 36594 45134
rect 36766 45110 36818 45162
rect 37046 45054 37098 45106
rect 37774 45082 37826 45134
rect 37998 45082 38050 45134
rect 38222 45110 38274 45162
rect 38334 45110 38386 45162
rect 38558 45054 38610 45106
rect 40910 45054 40962 45106
rect 41786 45054 41838 45106
rect 42702 45054 42754 45106
rect 43262 45081 43314 45133
rect 45726 45089 45778 45141
rect 45838 45110 45890 45162
rect 46062 45082 46114 45134
rect 46286 45110 46338 45162
rect 47294 45054 47346 45106
rect 47742 45093 47794 45145
rect 47966 45054 48018 45106
rect 48638 45054 48690 45106
rect 48862 45054 48914 45106
rect 49142 45054 49194 45106
rect 10222 44942 10274 44994
rect 12742 44942 12794 44994
rect 13918 44942 13970 44994
rect 14478 44942 14530 44994
rect 15710 44942 15762 44994
rect 19182 44942 19234 44994
rect 21086 44942 21138 44994
rect 24222 44942 24274 44994
rect 25678 44942 25730 44994
rect 28590 44942 28642 44994
rect 29542 44942 29594 44994
rect 35646 44942 35698 44994
rect 39510 44942 39562 44994
rect 16774 44830 16826 44882
rect 17446 44830 17498 44882
rect 42030 44830 42082 44882
rect 42534 44830 42586 44882
rect 46566 44830 46618 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 9102 44494 9154 44546
rect 19070 44494 19122 44546
rect 7422 44382 7474 44434
rect 12462 44382 12514 44434
rect 15822 44382 15874 44434
rect 24782 44382 24834 44434
rect 28534 44382 28586 44434
rect 30606 44438 30658 44490
rect 34638 44494 34690 44546
rect 37998 44494 38050 44546
rect 42534 44494 42586 44546
rect 43486 44494 43538 44546
rect 44046 44494 44098 44546
rect 45670 44494 45722 44546
rect 44830 44438 44882 44490
rect 35758 44382 35810 44434
rect 36990 44382 37042 44434
rect 40462 44382 40514 44434
rect 41470 44382 41522 44434
rect 46398 44382 46450 44434
rect 47742 44382 47794 44434
rect 7534 44226 7586 44278
rect 7870 44270 7922 44322
rect 9438 44270 9490 44322
rect 9886 44270 9938 44322
rect 12126 44242 12178 44294
rect 12574 44226 12626 44278
rect 12910 44270 12962 44322
rect 13358 44270 13410 44322
rect 13806 44270 13858 44322
rect 14926 44270 14978 44322
rect 15934 44226 15986 44278
rect 16158 44270 16210 44322
rect 17054 44270 17106 44322
rect 17614 44242 17666 44294
rect 17838 44242 17890 44294
rect 18062 44242 18114 44294
rect 18230 44254 18282 44306
rect 19406 44270 19458 44322
rect 19686 44270 19738 44322
rect 19966 44242 20018 44294
rect 20190 44214 20242 44266
rect 20414 44214 20466 44266
rect 20526 44235 20578 44287
rect 21758 44242 21810 44294
rect 23438 44270 23490 44322
rect 24446 44270 24498 44322
rect 25006 44270 25058 44322
rect 24670 44214 24722 44266
rect 27694 44214 27746 44266
rect 27806 44214 27858 44266
rect 28030 44242 28082 44294
rect 28254 44242 28306 44294
rect 29038 44270 29090 44322
rect 29262 44270 29314 44322
rect 29542 44270 29594 44322
rect 30158 44270 30210 44322
rect 30494 44270 30546 44322
rect 31166 44270 31218 44322
rect 31390 44214 31442 44266
rect 17334 44158 17386 44210
rect 31558 44214 31610 44266
rect 31726 44242 31778 44294
rect 32006 44235 32058 44287
rect 32622 44270 32674 44322
rect 32734 44270 32786 44322
rect 33518 44270 33570 44322
rect 34394 44270 34446 44322
rect 35198 44232 35250 44284
rect 35534 44270 35586 44322
rect 36094 44270 36146 44322
rect 35926 44214 35978 44266
rect 37102 44226 37154 44278
rect 37326 44270 37378 44322
rect 37662 44270 37714 44322
rect 41246 44270 41298 44322
rect 41806 44270 41858 44322
rect 42814 44270 42866 44322
rect 32230 44158 32282 44210
rect 33014 44158 33066 44210
rect 41638 44214 41690 44266
rect 42926 44270 42978 44322
rect 43150 44270 43202 44322
rect 44382 44270 44434 44322
rect 44942 44270 44994 44322
rect 45278 44270 45330 44322
rect 45950 44270 46002 44322
rect 46062 44270 46114 44322
rect 46510 44255 46562 44307
rect 46846 44270 46898 44322
rect 47294 44270 47346 44322
rect 47630 44255 47682 44307
rect 48302 44270 48354 44322
rect 38558 44158 38610 44210
rect 13526 44046 13578 44098
rect 13974 44046 14026 44098
rect 16718 44046 16770 44098
rect 18678 44046 18730 44098
rect 27414 44046 27466 44098
rect 30998 44046 31050 44098
rect 36262 44046 36314 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 11342 43654 11394 43706
rect 21982 43654 22034 43706
rect 6190 43486 6242 43538
rect 6974 43486 7026 43538
rect 9998 43486 10050 43538
rect 10558 43486 10610 43538
rect 10782 43530 10834 43582
rect 11678 43542 11730 43594
rect 11342 43486 11394 43538
rect 11902 43486 11954 43538
rect 12798 43486 12850 43538
rect 12910 43486 12962 43538
rect 13694 43486 13746 43538
rect 13806 43486 13858 43538
rect 14030 43486 14082 43538
rect 14814 43486 14866 43538
rect 16718 43486 16770 43538
rect 17278 43486 17330 43538
rect 17502 43486 17554 43538
rect 18174 43486 18226 43538
rect 18510 43486 18562 43538
rect 19406 43486 19458 43538
rect 19910 43542 19962 43594
rect 22766 43598 22818 43650
rect 20190 43514 20242 43566
rect 20414 43514 20466 43566
rect 20601 43542 20653 43594
rect 21870 43542 21922 43594
rect 28422 43598 28474 43650
rect 23009 43542 23061 43594
rect 21534 43486 21586 43538
rect 22094 43486 22146 43538
rect 24390 43542 24442 43594
rect 33406 43598 33458 43650
rect 43094 43654 43146 43706
rect 28702 43542 28754 43594
rect 23886 43486 23938 43538
rect 24558 43486 24610 43538
rect 25230 43486 25282 43538
rect 28926 43514 28978 43566
rect 29150 43514 29202 43566
rect 29262 43521 29314 43573
rect 29822 43486 29874 43538
rect 30158 43486 30210 43538
rect 30270 43486 30322 43538
rect 8878 43374 8930 43426
rect 10894 43374 10946 43426
rect 19686 43374 19738 43426
rect 18398 43318 18450 43370
rect 29990 43430 30042 43482
rect 31166 43486 31218 43538
rect 31838 43542 31890 43594
rect 31502 43486 31554 43538
rect 32174 43486 32226 43538
rect 33070 43486 33122 43538
rect 34750 43542 34802 43594
rect 21030 43374 21082 43426
rect 24222 43374 24274 43426
rect 26014 43374 26066 43426
rect 27918 43374 27970 43426
rect 30550 43374 30602 43426
rect 31838 43374 31890 43426
rect 33238 43430 33290 43482
rect 33518 43486 33570 43538
rect 34974 43514 35026 43566
rect 35142 43521 35194 43573
rect 35385 43542 35437 43594
rect 35758 43486 35810 43538
rect 36094 43486 36146 43538
rect 36542 43486 36594 43538
rect 37326 43486 37378 43538
rect 40462 43486 40514 43538
rect 40798 43486 40850 43538
rect 41470 43516 41522 43568
rect 41694 43542 41746 43594
rect 42926 43486 42978 43538
rect 43710 43514 43762 43566
rect 43934 43486 43986 43538
rect 44158 43486 44210 43538
rect 44326 43542 44378 43594
rect 44606 43542 44658 43594
rect 44718 43514 44770 43566
rect 44942 43542 44994 43594
rect 45166 43542 45218 43594
rect 41974 43430 42026 43482
rect 45726 43486 45778 43538
rect 45950 43486 46002 43538
rect 47294 43486 47346 43538
rect 47518 43486 47570 43538
rect 47854 43501 47906 43553
rect 48638 43486 48690 43538
rect 39230 43374 39282 43426
rect 9662 43262 9714 43314
rect 12518 43262 12570 43314
rect 13414 43262 13466 43314
rect 17782 43262 17834 43314
rect 19070 43262 19122 43314
rect 33798 43262 33850 43314
rect 34470 43262 34522 43314
rect 35646 43318 35698 43370
rect 47966 43374 48018 43426
rect 40126 43262 40178 43314
rect 40966 43318 41018 43370
rect 42254 43262 42306 43314
rect 45446 43262 45498 43314
rect 46230 43262 46282 43314
rect 46958 43262 47010 43314
rect 48974 43262 49026 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 7198 42926 7250 42978
rect 14590 42926 14642 42978
rect 16046 42926 16098 42978
rect 25454 42926 25506 42978
rect 29542 42926 29594 42978
rect 30326 42926 30378 42978
rect 37830 42926 37882 42978
rect 38446 42926 38498 42978
rect 42030 42926 42082 42978
rect 44102 42926 44154 42978
rect 18734 42814 18786 42866
rect 35310 42814 35362 42866
rect 47182 42814 47234 42866
rect 7441 42702 7493 42754
rect 8318 42702 8370 42754
rect 8766 42702 8818 42754
rect 9550 42702 9602 42754
rect 12238 42702 12290 42754
rect 12910 42702 12962 42754
rect 13470 42702 13522 42754
rect 14346 42702 14398 42754
rect 12574 42646 12626 42698
rect 15374 42674 15426 42726
rect 17950 42702 18002 42754
rect 21198 42702 21250 42754
rect 21646 42702 21698 42754
rect 22430 42702 22482 42754
rect 24782 42702 24834 42754
rect 25790 42702 25842 42754
rect 25902 42702 25954 42754
rect 27414 42702 27466 42754
rect 27694 42674 27746 42726
rect 27918 42674 27970 42726
rect 28142 42674 28194 42726
rect 11454 42590 11506 42642
rect 20638 42590 20690 42642
rect 12126 42534 12178 42586
rect 24334 42590 24386 42642
rect 28254 42646 28306 42698
rect 29038 42702 29090 42754
rect 29262 42702 29314 42754
rect 29822 42702 29874 42754
rect 30046 42702 30098 42754
rect 31166 42702 31218 42754
rect 31390 42663 31442 42715
rect 31838 42702 31890 42754
rect 32510 42702 32562 42754
rect 32790 42758 32842 42810
rect 32958 42702 33010 42754
rect 34078 42702 34130 42754
rect 32230 42590 32282 42642
rect 21366 42478 21418 42530
rect 24950 42534 25002 42586
rect 31278 42534 31330 42586
rect 34526 42646 34578 42698
rect 34750 42646 34802 42698
rect 35030 42646 35082 42698
rect 35422 42687 35474 42739
rect 35646 42702 35698 42754
rect 35982 42702 36034 42754
rect 32622 42590 32674 42642
rect 36990 42646 37042 42698
rect 37102 42674 37154 42726
rect 37326 42646 37378 42698
rect 37550 42674 37602 42726
rect 38110 42702 38162 42754
rect 38782 42702 38834 42754
rect 39790 42702 39842 42754
rect 40350 42702 40402 42754
rect 40910 42702 40962 42754
rect 41786 42702 41838 42754
rect 42366 42702 42418 42754
rect 42590 42702 42642 42754
rect 43374 42702 43426 42754
rect 43822 42702 43874 42754
rect 43542 42646 43594 42698
rect 45166 42702 45218 42754
rect 45390 42663 45442 42715
rect 45726 42702 45778 42754
rect 46398 42702 46450 42754
rect 42870 42590 42922 42642
rect 43710 42590 43762 42642
rect 36318 42478 36370 42530
rect 40462 42534 40514 42586
rect 49086 42590 49138 42642
rect 45614 42534 45666 42586
rect 39118 42478 39170 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 9998 42142 10050 42194
rect 34694 42142 34746 42194
rect 11230 42086 11282 42138
rect 18958 42030 19010 42082
rect 5854 41918 5906 41970
rect 6414 41918 6466 41970
rect 6638 41918 6690 41970
rect 6918 41918 6970 41970
rect 7198 41918 7250 41970
rect 7422 41918 7474 41970
rect 7758 41933 7810 41985
rect 8094 41918 8146 41970
rect 8878 41918 8930 41970
rect 9102 41918 9154 41970
rect 11566 41974 11618 42026
rect 10334 41918 10386 41970
rect 10894 41918 10946 41970
rect 11230 41918 11282 41970
rect 11790 41918 11842 41970
rect 12346 41956 12398 42008
rect 13582 41974 13634 42026
rect 13022 41918 13074 41970
rect 13694 41946 13746 41998
rect 13918 41946 13970 41998
rect 14142 41974 14194 42026
rect 15598 41953 15650 42005
rect 15710 41946 15762 41998
rect 15934 41946 15986 41998
rect 16158 41974 16210 42026
rect 16438 41918 16490 41970
rect 17390 41953 17442 42005
rect 17502 41974 17554 42026
rect 17726 41974 17778 42026
rect 17950 41974 18002 42026
rect 19798 42030 19850 42082
rect 18622 41918 18674 41970
rect 20078 41974 20130 42026
rect 20246 41974 20298 42026
rect 22262 42030 22314 42082
rect 29542 42030 29594 42082
rect 18790 41862 18842 41914
rect 19070 41918 19122 41970
rect 20526 41946 20578 41998
rect 20713 41974 20765 42026
rect 35590 42030 35642 42082
rect 42030 42030 42082 42082
rect 21646 41918 21698 41970
rect 21982 41918 22034 41970
rect 22542 41918 22594 41970
rect 22766 41918 22818 41970
rect 23774 41918 23826 41970
rect 25230 41918 25282 41970
rect 26462 41918 26514 41970
rect 28478 41945 28530 41997
rect 29766 41953 29818 42005
rect 30046 41946 30098 41998
rect 30270 41946 30322 41998
rect 30438 41934 30490 41986
rect 30718 41918 30770 41970
rect 31054 41918 31106 41970
rect 31502 41918 31554 41970
rect 31726 41918 31778 41970
rect 33742 41918 33794 41970
rect 34862 41918 34914 41970
rect 35870 41946 35922 41998
rect 36094 41974 36146 42026
rect 36318 41974 36370 42026
rect 36430 41953 36482 42005
rect 36654 41918 36706 41970
rect 37438 41918 37490 41970
rect 39678 41918 39730 41970
rect 41786 41974 41838 42026
rect 40910 41918 40962 41970
rect 42478 41918 42530 41970
rect 42590 41918 42642 41970
rect 42870 41918 42922 41970
rect 43486 41918 43538 41970
rect 44046 41974 44098 42026
rect 43822 41918 43874 41970
rect 44494 41918 44546 41970
rect 44718 41918 44770 41970
rect 45166 41918 45218 41970
rect 45838 41945 45890 41997
rect 47966 41918 48018 41970
rect 48638 41918 48690 41970
rect 7646 41806 7698 41858
rect 21142 41806 21194 41858
rect 10726 41750 10778 41802
rect 12798 41750 12850 41802
rect 28982 41806 29034 41858
rect 35254 41806 35306 41858
rect 39342 41806 39394 41858
rect 44270 41806 44322 41858
rect 5518 41694 5570 41746
rect 6134 41694 6186 41746
rect 8598 41694 8650 41746
rect 14422 41694 14474 41746
rect 18230 41694 18282 41746
rect 19350 41694 19402 41746
rect 23942 41694 23994 41746
rect 30942 41750 30994 41802
rect 25398 41694 25450 41746
rect 32006 41694 32058 41746
rect 34078 41694 34130 41746
rect 40014 41694 40066 41746
rect 44886 41694 44938 41746
rect 45334 41694 45386 41746
rect 48974 41694 49026 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 10222 41302 10274 41354
rect 10614 41358 10666 41410
rect 17502 41358 17554 41410
rect 6302 41246 6354 41298
rect 31390 41302 31442 41354
rect 40462 41358 40514 41410
rect 43094 41358 43146 41410
rect 15486 41246 15538 41298
rect 16046 41246 16098 41298
rect 29542 41246 29594 41298
rect 35198 41246 35250 41298
rect 45502 41246 45554 41298
rect 5518 41134 5570 41186
rect 8542 41134 8594 41186
rect 8766 41134 8818 41186
rect 9886 41134 9938 41186
rect 10110 41134 10162 41186
rect 10446 41134 10498 41186
rect 10894 41134 10946 41186
rect 11678 41134 11730 41186
rect 12554 41078 12606 41130
rect 13470 41101 13522 41153
rect 13806 41101 13858 41153
rect 14310 41078 14362 41130
rect 14564 41094 14616 41146
rect 15038 41134 15090 41186
rect 15374 41090 15426 41142
rect 16158 41119 16210 41171
rect 16494 41134 16546 41186
rect 16830 41134 16882 41186
rect 16942 41134 16994 41186
rect 17110 41134 17162 41186
rect 19966 41134 20018 41186
rect 21870 41134 21922 41186
rect 22878 41134 22930 41186
rect 23550 41134 23602 41186
rect 23774 41134 23826 41186
rect 8206 41022 8258 41074
rect 9046 41022 9098 41074
rect 12798 41022 12850 41074
rect 23214 41078 23266 41130
rect 24446 41134 24498 41186
rect 25230 41134 25282 41186
rect 27918 41106 27970 41158
rect 14702 41022 14754 41074
rect 27134 41022 27186 41074
rect 11062 40910 11114 40962
rect 18118 40910 18170 40962
rect 19630 40910 19682 40962
rect 20358 40910 20410 40962
rect 20806 40910 20858 40962
rect 23438 40966 23490 41018
rect 28142 41078 28194 41130
rect 28366 41078 28418 41130
rect 28478 41078 28530 41130
rect 29038 41134 29090 41186
rect 29262 41134 29314 41186
rect 29822 41134 29874 41186
rect 30046 41134 30098 41186
rect 30942 41134 30994 41186
rect 31278 41134 31330 41186
rect 31614 41134 31666 41186
rect 31838 41134 31890 41186
rect 33294 41134 33346 41186
rect 35982 41134 36034 41186
rect 37662 41134 37714 41186
rect 39902 41106 39954 41158
rect 40126 41134 40178 41186
rect 42254 41099 42306 41151
rect 44382 41134 44434 41186
rect 44942 41134 44994 41186
rect 45166 41134 45218 41186
rect 45726 41134 45778 41186
rect 45950 41134 46002 41186
rect 48526 41134 48578 41186
rect 49310 41134 49362 41186
rect 42366 41078 42418 41130
rect 42590 41078 42642 41130
rect 42814 41078 42866 41130
rect 27638 41022 27690 41074
rect 30326 41022 30378 41074
rect 32118 41022 32170 41074
rect 46622 41022 46674 41074
rect 22374 40910 22426 40962
rect 24110 40910 24162 40962
rect 36486 40910 36538 40962
rect 37158 40910 37210 40962
rect 41078 40910 41130 40962
rect 41526 40910 41578 40962
rect 41974 40910 42026 40962
rect 43878 40910 43930 40962
rect 44214 40910 44266 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 24110 40518 24162 40570
rect 25790 40518 25842 40570
rect 20750 40462 20802 40514
rect 34470 40574 34522 40626
rect 26630 40518 26682 40570
rect 30270 40518 30322 40570
rect 41526 40574 41578 40626
rect 41974 40574 42026 40626
rect 46454 40574 46506 40626
rect 5406 40350 5458 40402
rect 6638 40377 6690 40429
rect 11454 40406 11506 40458
rect 13246 40406 13298 40458
rect 28142 40462 28194 40514
rect 28982 40462 29034 40514
rect 8318 40350 8370 40402
rect 9550 40350 9602 40402
rect 9886 40350 9938 40402
rect 10446 40350 10498 40402
rect 10670 40350 10722 40402
rect 11118 40350 11170 40402
rect 11790 40350 11842 40402
rect 12910 40350 12962 40402
rect 13582 40350 13634 40402
rect 13918 40350 13970 40402
rect 14478 40350 14530 40402
rect 14814 40350 14866 40402
rect 15822 40350 15874 40402
rect 16158 40350 16210 40402
rect 16382 40389 16434 40441
rect 33910 40462 33962 40514
rect 16830 40350 16882 40402
rect 17726 40350 17778 40402
rect 19630 40350 19682 40402
rect 20414 40350 20466 40402
rect 23438 40350 23490 40402
rect 23998 40350 24050 40402
rect 24334 40377 24386 40429
rect 24558 40350 24610 40402
rect 25454 40350 25506 40402
rect 25678 40389 25730 40441
rect 26126 40350 26178 40402
rect 26798 40350 26850 40402
rect 27022 40350 27074 40402
rect 27898 40350 27950 40402
rect 28478 40350 28530 40402
rect 28702 40350 28754 40402
rect 29934 40406 29986 40458
rect 31222 40406 31274 40458
rect 29710 40350 29762 40402
rect 30382 40350 30434 40402
rect 31054 40350 31106 40402
rect 31614 40350 31666 40402
rect 31950 40350 32002 40402
rect 33070 40406 33122 40458
rect 33182 40378 33234 40430
rect 33406 40378 33458 40430
rect 33630 40406 33682 40458
rect 34862 40350 34914 40402
rect 35198 40350 35250 40402
rect 35310 40350 35362 40402
rect 36430 40406 36482 40458
rect 37270 40462 37322 40514
rect 40238 40462 40290 40514
rect 36542 40378 36594 40430
rect 36766 40378 36818 40430
rect 36990 40378 37042 40430
rect 42926 40406 42978 40458
rect 37550 40350 37602 40402
rect 38334 40350 38386 40402
rect 41358 40350 41410 40402
rect 41806 40350 41858 40402
rect 42590 40350 42642 40402
rect 43654 40350 43706 40402
rect 10110 40238 10162 40290
rect 42814 40294 42866 40346
rect 43990 40350 44042 40402
rect 44214 40406 44266 40458
rect 48078 40462 48130 40514
rect 44494 40378 44546 40430
rect 44718 40378 44770 40430
rect 44886 40366 44938 40418
rect 45091 40406 45143 40458
rect 45278 40378 45330 40430
rect 45502 40406 45554 40458
rect 45782 40406 45834 40458
rect 47834 40406 47886 40458
rect 46286 40350 46338 40402
rect 46958 40350 47010 40402
rect 48862 40365 48914 40417
rect 49086 40350 49138 40402
rect 11454 40238 11506 40290
rect 13134 40238 13186 40290
rect 16494 40238 16546 40290
rect 22654 40238 22706 40290
rect 31278 40238 31330 40290
rect 14814 40182 14866 40234
rect 43486 40238 43538 40290
rect 48750 40238 48802 40290
rect 42422 40126 42474 40178
rect 46006 40126 46058 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 8822 39734 8874 39786
rect 17278 39790 17330 39842
rect 19686 39790 19738 39842
rect 24950 39790 25002 39842
rect 25454 39790 25506 39842
rect 29486 39790 29538 39842
rect 5630 39678 5682 39730
rect 11454 39678 11506 39730
rect 16158 39678 16210 39730
rect 24278 39678 24330 39730
rect 30606 39734 30658 39786
rect 31278 39734 31330 39786
rect 37830 39790 37882 39842
rect 44886 39790 44938 39842
rect 26406 39678 26458 39730
rect 5742 39522 5794 39574
rect 5966 39566 6018 39618
rect 6638 39566 6690 39618
rect 6862 39527 6914 39579
rect 7310 39566 7362 39618
rect 7646 39510 7698 39562
rect 7758 39528 7810 39580
rect 8486 39566 8538 39618
rect 8654 39566 8706 39618
rect 9214 39531 9266 39583
rect 9382 39531 9434 39583
rect 9550 39510 9602 39562
rect 9774 39538 9826 39590
rect 10782 39566 10834 39618
rect 10894 39566 10946 39618
rect 8318 39454 8370 39506
rect 6526 39398 6578 39450
rect 11060 39510 11112 39562
rect 12014 39531 12066 39583
rect 12126 39510 12178 39562
rect 12406 39510 12458 39562
rect 12574 39538 12626 39590
rect 14254 39566 14306 39618
rect 14926 39566 14978 39618
rect 15486 39566 15538 39618
rect 15598 39566 15650 39618
rect 15764 39566 15816 39618
rect 10054 39454 10106 39506
rect 14646 39510 14698 39562
rect 16606 39566 16658 39618
rect 16718 39566 16770 39618
rect 18174 39566 18226 39618
rect 16884 39510 16936 39562
rect 19406 39566 19458 39618
rect 19966 39538 20018 39590
rect 12854 39454 12906 39506
rect 20190 39510 20242 39562
rect 20414 39510 20466 39562
rect 20526 39510 20578 39562
rect 21646 39538 21698 39590
rect 23326 39566 23378 39618
rect 24446 39566 24498 39618
rect 24670 39566 24722 39618
rect 25790 39566 25842 39618
rect 27694 39566 27746 39618
rect 27862 39622 27914 39674
rect 32174 39678 32226 39730
rect 35086 39678 35138 39730
rect 38894 39678 38946 39730
rect 40798 39678 40850 39730
rect 46398 39678 46450 39730
rect 47630 39678 47682 39730
rect 48750 39678 48802 39730
rect 28142 39566 28194 39618
rect 28422 39566 28474 39618
rect 29878 39566 29930 39618
rect 30046 39566 30098 39618
rect 30158 39566 30210 39618
rect 30494 39566 30546 39618
rect 30830 39566 30882 39618
rect 31390 39566 31442 39618
rect 31614 39566 31666 39618
rect 32734 39566 32786 39618
rect 32846 39566 32898 39618
rect 34638 39566 34690 39618
rect 19070 39454 19122 39506
rect 32568 39510 32620 39562
rect 34974 39551 35026 39603
rect 35422 39566 35474 39618
rect 36990 39531 37042 39583
rect 37102 39510 37154 39562
rect 37326 39538 37378 39590
rect 38110 39566 38162 39618
rect 42814 39566 42866 39618
rect 43486 39566 43538 39618
rect 45054 39566 45106 39618
rect 45614 39566 45666 39618
rect 37550 39510 37602 39562
rect 43262 39510 43314 39562
rect 48918 39622 48970 39674
rect 45950 39566 46002 39618
rect 46510 39566 46562 39618
rect 46958 39566 47010 39618
rect 47070 39566 47122 39618
rect 46174 39510 46226 39562
rect 47236 39510 47288 39562
rect 48190 39528 48242 39580
rect 48526 39566 48578 39618
rect 14142 39398 14194 39450
rect 28030 39454 28082 39506
rect 18510 39342 18562 39394
rect 33350 39342 33402 39394
rect 33798 39342 33850 39394
rect 34358 39342 34410 39394
rect 35758 39342 35810 39394
rect 36486 39342 36538 39394
rect 41638 39342 41690 39394
rect 42086 39342 42138 39394
rect 43038 39398 43090 39450
rect 42534 39342 42586 39394
rect 44326 39342 44378 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 11790 39006 11842 39058
rect 6526 38894 6578 38946
rect 12574 38950 12626 39002
rect 14646 38950 14698 39002
rect 25454 39006 25506 39058
rect 26126 39006 26178 39058
rect 29262 39006 29314 39058
rect 29934 39006 29986 39058
rect 10446 38894 10498 38946
rect 44606 38950 44658 39002
rect 48974 39006 49026 39058
rect 6769 38838 6821 38890
rect 5406 38782 5458 38834
rect 6190 38782 6242 38834
rect 7646 38782 7698 38834
rect 8598 38782 8650 38834
rect 8878 38782 8930 38834
rect 9102 38782 9154 38834
rect 9494 38838 9546 38890
rect 9662 38838 9714 38890
rect 15710 38894 15762 38946
rect 9886 38821 9938 38873
rect 12910 38838 12962 38890
rect 16438 38894 16490 38946
rect 11006 38782 11058 38834
rect 11342 38782 11394 38834
rect 12126 38782 12178 38834
rect 12462 38782 12514 38834
rect 13134 38782 13186 38834
rect 14814 38782 14866 38834
rect 15262 38810 15314 38862
rect 15878 38838 15930 38890
rect 15486 38782 15538 38834
rect 16718 38782 16770 38834
rect 16942 38782 16994 38834
rect 20638 38782 20690 38834
rect 20974 38826 21026 38878
rect 21310 38782 21362 38834
rect 22094 38782 22146 38834
rect 22318 38797 22370 38849
rect 22934 38838 22986 38890
rect 23102 38782 23154 38834
rect 23886 38797 23938 38849
rect 24222 38782 24274 38834
rect 25118 38782 25170 38834
rect 25790 38782 25842 38834
rect 26462 38782 26514 38834
rect 26686 38782 26738 38834
rect 26966 38782 27018 38834
rect 27246 38782 27298 38834
rect 28814 38782 28866 38834
rect 28926 38782 28978 38834
rect 30662 38838 30714 38890
rect 31222 38838 31274 38890
rect 29598 38782 29650 38834
rect 30830 38782 30882 38834
rect 31614 38838 31666 38890
rect 31726 38838 31778 38890
rect 31950 38838 32002 38890
rect 32174 38810 32226 38862
rect 33182 38782 33234 38834
rect 35870 38782 35922 38834
rect 35982 38782 36034 38834
rect 36766 38817 36818 38869
rect 36878 38838 36930 38890
rect 37102 38838 37154 38890
rect 37364 38798 37416 38850
rect 37606 38782 37658 38834
rect 37998 38782 38050 38834
rect 40798 38782 40850 38834
rect 44270 38782 44322 38834
rect 44606 38809 44658 38861
rect 44830 38782 44882 38834
rect 45278 38782 45330 38834
rect 45390 38782 45442 38834
rect 45576 38819 45628 38871
rect 46846 38782 46898 38834
rect 47070 38817 47122 38869
rect 47238 38817 47290 38869
rect 47406 38810 47458 38862
rect 47680 38810 47732 38862
rect 48638 38782 48690 38834
rect 3502 38670 3554 38722
rect 8262 38670 8314 38722
rect 17558 38670 17610 38722
rect 17950 38670 18002 38722
rect 19854 38670 19906 38722
rect 20862 38670 20914 38722
rect 22430 38670 22482 38722
rect 22766 38670 22818 38722
rect 23774 38670 23826 38722
rect 24726 38670 24778 38722
rect 11118 38614 11170 38666
rect 27582 38670 27634 38722
rect 28478 38670 28530 38722
rect 31054 38670 31106 38722
rect 32454 38670 32506 38722
rect 35086 38670 35138 38722
rect 38950 38670 39002 38722
rect 41582 38670 41634 38722
rect 43486 38670 43538 38722
rect 45950 38670 46002 38722
rect 46510 38670 46562 38722
rect 36318 38558 36370 38610
rect 38334 38558 38386 38610
rect 47910 38558 47962 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 10614 38222 10666 38274
rect 11678 38222 11730 38274
rect 16550 38222 16602 38274
rect 23214 38166 23266 38218
rect 30102 38222 30154 38274
rect 30886 38222 30938 38274
rect 31782 38222 31834 38274
rect 33294 38222 33346 38274
rect 34806 38222 34858 38274
rect 45950 38222 46002 38274
rect 8206 38110 8258 38162
rect 9214 38110 9266 38162
rect 18734 38110 18786 38162
rect 21422 38110 21474 38162
rect 24110 38110 24162 38162
rect 26574 38110 26626 38162
rect 28478 38110 28530 38162
rect 38558 38110 38610 38162
rect 40462 38110 40514 38162
rect 41694 38110 41746 38162
rect 43710 38110 43762 38162
rect 46622 38110 46674 38162
rect 48526 38110 48578 38162
rect 5518 37998 5570 38050
rect 6302 37998 6354 38050
rect 8654 37998 8706 38050
rect 8990 37998 9042 38050
rect 9550 37998 9602 38050
rect 9774 37998 9826 38050
rect 10110 37998 10162 38050
rect 10334 37998 10386 38050
rect 12014 37998 12066 38050
rect 12350 37998 12402 38050
rect 12574 37998 12626 38050
rect 13358 37998 13410 38050
rect 14142 37998 14194 38050
rect 16046 37998 16098 38050
rect 16830 37970 16882 38022
rect 16998 37963 17050 38015
rect 17278 37942 17330 37994
rect 17390 37963 17442 38015
rect 17614 37998 17666 38050
rect 18398 37998 18450 38050
rect 18622 37954 18674 38006
rect 18958 37998 19010 38050
rect 19294 37998 19346 38050
rect 20302 37998 20354 38050
rect 20582 37998 20634 38050
rect 20750 37998 20802 38050
rect 21310 37998 21362 38050
rect 21982 37998 22034 38050
rect 12854 37886 12906 37938
rect 20022 37886 20074 37938
rect 21646 37942 21698 37994
rect 22318 37998 22370 38050
rect 23326 37998 23378 38050
rect 23662 37998 23714 38050
rect 23998 37998 24050 38050
rect 24446 37959 24498 38011
rect 24670 37998 24722 38050
rect 25006 37998 25058 38050
rect 25790 37998 25842 38050
rect 29262 37963 29314 38015
rect 29374 37942 29426 37994
rect 29598 37970 29650 38022
rect 30382 37998 30434 38050
rect 29822 37942 29874 37994
rect 30606 37998 30658 38050
rect 31614 37998 31666 38050
rect 32958 37998 33010 38050
rect 31502 37942 31554 37994
rect 35086 37998 35138 38050
rect 35310 37998 35362 38050
rect 20414 37886 20466 37938
rect 35534 37942 35586 37994
rect 35646 37970 35698 38022
rect 35926 37963 35978 38015
rect 36374 37998 36426 38050
rect 36094 37942 36146 37994
rect 36878 37998 36930 38050
rect 37774 37998 37826 38050
rect 41246 37998 41298 38050
rect 41582 37983 41634 38035
rect 42254 37998 42306 38050
rect 42497 37998 42549 38050
rect 43374 37998 43426 38050
rect 43822 37954 43874 38006
rect 44158 37998 44210 38050
rect 44718 37998 44770 38050
rect 44942 37998 44994 38050
rect 46286 37998 46338 38050
rect 49310 37998 49362 38050
rect 45222 37886 45274 37938
rect 17782 37774 17834 37826
rect 31334 37830 31386 37882
rect 32790 37774 32842 37826
rect 33910 37774 33962 37826
rect 34470 37774 34522 37826
rect 37214 37774 37266 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 8598 37438 8650 37490
rect 9606 37438 9658 37490
rect 13582 37438 13634 37490
rect 15822 37438 15874 37490
rect 16774 37438 16826 37490
rect 19126 37438 19178 37490
rect 21086 37438 21138 37490
rect 25734 37438 25786 37490
rect 28310 37438 28362 37490
rect 30998 37438 31050 37490
rect 45110 37438 45162 37490
rect 12910 37326 12962 37378
rect 6246 37270 6298 37322
rect 17502 37326 17554 37378
rect 24222 37326 24274 37378
rect 5966 37214 6018 37266
rect 8430 37214 8482 37266
rect 9774 37214 9826 37266
rect 10222 37214 10274 37266
rect 13246 37214 13298 37266
rect 17745 37270 17797 37322
rect 27134 37326 27186 37378
rect 31894 37326 31946 37378
rect 32398 37326 32450 37378
rect 34414 37326 34466 37378
rect 16158 37214 16210 37266
rect 16942 37214 16994 37266
rect 18622 37214 18674 37266
rect 19854 37214 19906 37266
rect 20190 37214 20242 37266
rect 20526 37214 20578 37266
rect 21422 37214 21474 37266
rect 21534 37214 21586 37266
rect 22318 37214 22370 37266
rect 26014 37214 26066 37266
rect 26890 37214 26942 37266
rect 28590 37214 28642 37266
rect 28926 37229 28978 37281
rect 29262 37214 29314 37266
rect 30158 37214 30210 37266
rect 30830 37214 30882 37266
rect 32062 37214 32114 37266
rect 34170 37270 34222 37322
rect 39118 37326 39170 37378
rect 41694 37382 41746 37434
rect 45950 37438 46002 37490
rect 47070 37382 47122 37434
rect 40406 37326 40458 37378
rect 33294 37214 33346 37266
rect 35758 37214 35810 37266
rect 36430 37214 36482 37266
rect 37214 37214 37266 37266
rect 41022 37214 41074 37266
rect 41246 37241 41298 37293
rect 41582 37214 41634 37266
rect 42366 37214 42418 37266
rect 44270 37241 44322 37293
rect 46790 37270 46842 37322
rect 44942 37214 44994 37266
rect 46286 37214 46338 37266
rect 46622 37214 46674 37266
rect 47182 37214 47234 37266
rect 47742 37214 47794 37266
rect 48078 37214 48130 37266
rect 49310 37214 49362 37266
rect 6414 37102 6466 37154
rect 11006 37102 11058 37154
rect 19518 36990 19570 37042
rect 20078 37046 20130 37098
rect 27750 37102 27802 37154
rect 29038 37102 29090 37154
rect 36150 37102 36202 37154
rect 39734 37102 39786 37154
rect 29598 36990 29650 37042
rect 30494 36990 30546 37042
rect 48190 37046 48242 37098
rect 48974 36990 49026 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 11454 36654 11506 36706
rect 14926 36654 14978 36706
rect 9998 36542 10050 36594
rect 17726 36542 17778 36594
rect 20806 36542 20858 36594
rect 21702 36542 21754 36594
rect 22150 36542 22202 36594
rect 22542 36598 22594 36650
rect 23382 36654 23434 36706
rect 37102 36654 37154 36706
rect 44942 36598 44994 36650
rect 27022 36542 27074 36594
rect 29822 36542 29874 36594
rect 31726 36542 31778 36594
rect 35758 36542 35810 36594
rect 43710 36542 43762 36594
rect 6638 36430 6690 36482
rect 7310 36430 7362 36482
rect 8094 36430 8146 36482
rect 11790 36430 11842 36482
rect 12070 36430 12122 36482
rect 12294 36395 12346 36447
rect 12574 36402 12626 36454
rect 12798 36374 12850 36426
rect 12966 36414 13018 36466
rect 14590 36430 14642 36482
rect 16382 36374 16434 36426
rect 16494 36374 16546 36426
rect 16718 36402 16770 36454
rect 16942 36402 16994 36454
rect 19630 36430 19682 36482
rect 20414 36430 20466 36482
rect 22654 36430 22706 36482
rect 22878 36430 22930 36482
rect 23662 36430 23714 36482
rect 23942 36486 23994 36538
rect 24110 36430 24162 36482
rect 24334 36430 24386 36482
rect 25118 36430 25170 36482
rect 27750 36395 27802 36447
rect 28030 36402 28082 36454
rect 17222 36318 17274 36370
rect 23774 36318 23826 36370
rect 28254 36374 28306 36426
rect 28366 36374 28418 36426
rect 32510 36430 32562 36482
rect 33182 36430 33234 36482
rect 36542 36430 36594 36482
rect 37438 36430 37490 36482
rect 38278 36430 38330 36482
rect 39342 36430 39394 36482
rect 41582 36430 41634 36482
rect 42366 36430 42418 36482
rect 42478 36409 42530 36461
rect 43822 36415 43874 36467
rect 44046 36430 44098 36482
rect 44830 36430 44882 36482
rect 45166 36430 45218 36482
rect 45614 36430 45666 36482
rect 45838 36430 45890 36482
rect 48526 36430 48578 36482
rect 49310 36430 49362 36482
rect 27526 36318 27578 36370
rect 29318 36318 29370 36370
rect 33854 36318 33906 36370
rect 39678 36318 39730 36370
rect 46118 36318 46170 36370
rect 46622 36318 46674 36370
rect 6302 36206 6354 36258
rect 13638 36206 13690 36258
rect 16102 36206 16154 36258
rect 32846 36206 32898 36258
rect 37830 36206 37882 36258
rect 39006 36206 39058 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 8766 35870 8818 35922
rect 18398 35870 18450 35922
rect 19182 35870 19234 35922
rect 24166 35870 24218 35922
rect 25790 35870 25842 35922
rect 31222 35870 31274 35922
rect 31614 35870 31666 35922
rect 35422 35870 35474 35922
rect 39622 35870 39674 35922
rect 42366 35870 42418 35922
rect 7870 35758 7922 35810
rect 16158 35758 16210 35810
rect 5182 35646 5234 35698
rect 5966 35646 6018 35698
rect 9102 35646 9154 35698
rect 9886 35702 9938 35754
rect 9606 35646 9658 35698
rect 10110 35674 10162 35726
rect 10334 35674 10386 35726
rect 10502 35662 10554 35714
rect 12238 35702 12290 35754
rect 12462 35702 12514 35754
rect 12686 35702 12738 35754
rect 21198 35758 21250 35810
rect 30102 35758 30154 35810
rect 40238 35814 40290 35866
rect 41022 35814 41074 35866
rect 12798 35681 12850 35733
rect 13470 35646 13522 35698
rect 14254 35646 14306 35698
rect 17502 35646 17554 35698
rect 17726 35646 17778 35698
rect 18734 35646 18786 35698
rect 18846 35646 18898 35698
rect 20078 35646 20130 35698
rect 20302 35646 20354 35698
rect 20806 35646 20858 35698
rect 21086 35646 21138 35698
rect 10950 35534 11002 35586
rect 16886 35534 16938 35586
rect 21366 35590 21418 35642
rect 21534 35646 21586 35698
rect 22766 35646 22818 35698
rect 23438 35646 23490 35698
rect 25398 35646 25450 35698
rect 26126 35646 26178 35698
rect 27134 35674 27186 35726
rect 27358 35702 27410 35754
rect 27582 35674 27634 35726
rect 27694 35702 27746 35754
rect 29038 35646 29090 35698
rect 29262 35681 29314 35733
rect 29374 35674 29426 35726
rect 29598 35702 29650 35754
rect 29822 35702 29874 35754
rect 31950 35646 32002 35698
rect 32062 35646 32114 35698
rect 33182 35646 33234 35698
rect 33518 35646 33570 35698
rect 34414 35646 34466 35698
rect 37102 35673 37154 35725
rect 37326 35646 37378 35698
rect 38558 35646 38610 35698
rect 39230 35646 39282 35698
rect 39902 35646 39954 35698
rect 40238 35661 40290 35713
rect 41022 35646 41074 35698
rect 41246 35673 41298 35725
rect 42030 35646 42082 35698
rect 22374 35534 22426 35586
rect 11958 35422 12010 35474
rect 17838 35478 17890 35530
rect 20190 35478 20242 35530
rect 23102 35534 23154 35586
rect 24614 35534 24666 35586
rect 26518 35534 26570 35586
rect 28198 35534 28250 35586
rect 30662 35534 30714 35586
rect 41582 35590 41634 35642
rect 42702 35646 42754 35698
rect 43486 35646 43538 35698
rect 45838 35646 45890 35698
rect 46174 35673 46226 35725
rect 46510 35646 46562 35698
rect 46846 35646 46898 35698
rect 47518 35661 47570 35713
rect 47742 35646 47794 35698
rect 48862 35690 48914 35742
rect 49086 35646 49138 35698
rect 37662 35534 37714 35586
rect 45390 35534 45442 35586
rect 45950 35534 46002 35586
rect 47406 35534 47458 35586
rect 48750 35534 48802 35586
rect 26854 35422 26906 35474
rect 28702 35422 28754 35474
rect 33294 35478 33346 35530
rect 32398 35422 32450 35474
rect 34078 35422 34130 35474
rect 38222 35422 38274 35474
rect 38894 35422 38946 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 14422 35086 14474 35138
rect 7422 34974 7474 35026
rect 23438 34974 23490 35026
rect 28478 34974 28530 35026
rect 34078 34974 34130 35026
rect 35646 35030 35698 35082
rect 37774 35030 37826 35082
rect 43598 35086 43650 35138
rect 44886 35086 44938 35138
rect 35982 34974 36034 35026
rect 38782 34974 38834 35026
rect 47182 34974 47234 35026
rect 4846 34862 4898 34914
rect 6190 34862 6242 34914
rect 6638 34834 6690 34886
rect 10110 34862 10162 34914
rect 10894 34862 10946 34914
rect 14646 34827 14698 34879
rect 14926 34834 14978 34886
rect 15150 34834 15202 34886
rect 15822 34862 15874 34914
rect 17502 34862 17554 34914
rect 20078 34862 20130 34914
rect 20862 34862 20914 34914
rect 12798 34750 12850 34802
rect 15262 34806 15314 34858
rect 24222 34862 24274 34914
rect 25790 34862 25842 34914
rect 26574 34862 26626 34914
rect 29038 34862 29090 34914
rect 29822 34862 29874 34914
rect 32734 34862 32786 34914
rect 18174 34750 18226 34802
rect 21534 34750 21586 34802
rect 24446 34806 24498 34858
rect 24558 34806 24610 34858
rect 24782 34806 24834 34858
rect 25006 34806 25058 34858
rect 32958 34862 33010 34914
rect 33742 34918 33794 34970
rect 33406 34862 33458 34914
rect 34302 34862 34354 34914
rect 34918 34862 34970 34914
rect 35198 34862 35250 34914
rect 35534 34862 35586 34914
rect 25286 34750 25338 34802
rect 34078 34806 34130 34858
rect 36094 34847 36146 34899
rect 36430 34862 36482 34914
rect 36934 34815 36986 34867
rect 37662 34862 37714 34914
rect 37998 34862 38050 34914
rect 40686 34862 40738 34914
rect 41694 34862 41746 34914
rect 42254 34862 42306 34914
rect 42590 34862 42642 34914
rect 43262 34862 43314 34914
rect 42030 34806 42082 34858
rect 45166 34862 45218 34914
rect 45278 34862 45330 34914
rect 45614 34862 45666 34914
rect 45446 34806 45498 34858
rect 46286 34806 46338 34858
rect 46398 34862 46450 34914
rect 31726 34750 31778 34802
rect 32454 34750 32506 34802
rect 5854 34638 5906 34690
rect 9382 34638 9434 34690
rect 9942 34638 9994 34690
rect 15654 34638 15706 34690
rect 16214 34638 16266 34690
rect 16774 34638 16826 34690
rect 17334 34638 17386 34690
rect 42142 34694 42194 34746
rect 42758 34694 42810 34746
rect 49086 34750 49138 34802
rect 17670 34638 17722 34690
rect 44326 34638 44378 34690
rect 46118 34638 46170 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 12238 34302 12290 34354
rect 12854 34302 12906 34354
rect 27246 34302 27298 34354
rect 9606 34190 9658 34242
rect 19854 34246 19906 34298
rect 30270 34302 30322 34354
rect 31670 34302 31722 34354
rect 34974 34302 35026 34354
rect 43094 34302 43146 34354
rect 44158 34302 44210 34354
rect 47966 34302 48018 34354
rect 17502 34190 17554 34242
rect 5518 34078 5570 34130
rect 6302 34078 6354 34130
rect 8206 34078 8258 34130
rect 9886 34134 9938 34186
rect 9102 34078 9154 34130
rect 10110 34106 10162 34158
rect 10334 34106 10386 34158
rect 10446 34134 10498 34186
rect 11118 34134 11170 34186
rect 33742 34190 33794 34242
rect 10838 34078 10890 34130
rect 11286 34113 11338 34165
rect 11566 34106 11618 34158
rect 11678 34113 11730 34165
rect 11902 34078 11954 34130
rect 13022 34078 13074 34130
rect 16382 34078 16434 34130
rect 16718 34122 16770 34174
rect 17745 34078 17797 34130
rect 18622 34078 18674 34130
rect 19014 34078 19066 34130
rect 19294 34078 19346 34130
rect 19518 34078 19570 34130
rect 19742 34078 19794 34130
rect 20078 34122 20130 34174
rect 20638 34078 20690 34130
rect 21086 34117 21138 34169
rect 21310 34078 21362 34130
rect 21646 34078 21698 34130
rect 22206 34105 22258 34157
rect 25118 34078 25170 34130
rect 26518 34078 26570 34130
rect 26910 34078 26962 34130
rect 28814 34134 28866 34186
rect 28926 34134 28978 34186
rect 29150 34134 29202 34186
rect 29374 34134 29426 34186
rect 29654 34078 29706 34130
rect 29934 34078 29986 34130
rect 31278 34078 31330 34130
rect 33574 34134 33626 34186
rect 37998 34190 38050 34242
rect 41078 34190 41130 34242
rect 33406 34078 33458 34130
rect 33854 34078 33906 34130
rect 34638 34078 34690 34130
rect 35310 34078 35362 34130
rect 36094 34078 36146 34130
rect 38558 34108 38610 34160
rect 38894 34134 38946 34186
rect 39062 34134 39114 34186
rect 40238 34078 40290 34130
rect 41358 34078 41410 34130
rect 41582 34078 41634 34130
rect 41918 34122 41970 34174
rect 42142 34078 42194 34130
rect 42478 34078 42530 34130
rect 42926 34078 42978 34130
rect 43654 34078 43706 34130
rect 43822 34078 43874 34130
rect 44718 34108 44770 34160
rect 44942 34117 44994 34169
rect 45222 34134 45274 34186
rect 45502 34190 45554 34242
rect 47294 34190 47346 34242
rect 47050 34134 47102 34186
rect 46174 34078 46226 34130
rect 47630 34078 47682 34130
rect 49310 34078 49362 34130
rect 13806 33966 13858 34018
rect 15710 33966 15762 34018
rect 16830 33966 16882 34018
rect 20974 33966 21026 34018
rect 26070 33966 26122 34018
rect 41806 33966 41858 34018
rect 48974 33966 49026 34018
rect 8766 33854 8818 33906
rect 23214 33854 23266 33906
rect 25454 33854 25506 33906
rect 30942 33854 30994 33906
rect 34134 33854 34186 33906
rect 39342 33854 39394 33906
rect 39902 33854 39954 33906
rect 42646 33854 42698 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 10166 33518 10218 33570
rect 15038 33462 15090 33514
rect 22374 33518 22426 33570
rect 38110 33518 38162 33570
rect 41974 33518 42026 33570
rect 7758 33406 7810 33458
rect 11454 33406 11506 33458
rect 12910 33406 12962 33458
rect 16606 33406 16658 33458
rect 18510 33406 18562 33458
rect 23774 33406 23826 33458
rect 25678 33406 25730 33458
rect 30494 33406 30546 33458
rect 32398 33406 32450 33458
rect 33854 33406 33906 33458
rect 35758 33406 35810 33458
rect 46622 33406 46674 33458
rect 6974 33294 7026 33346
rect 9662 33294 9714 33346
rect 10446 33266 10498 33318
rect 10670 33238 10722 33290
rect 10894 33238 10946 33290
rect 11006 33238 11058 33290
rect 11510 33264 11562 33316
rect 11902 33294 11954 33346
rect 12462 33294 12514 33346
rect 12798 33279 12850 33331
rect 13582 33294 13634 33346
rect 14702 33294 14754 33346
rect 15150 33294 15202 33346
rect 15486 33294 15538 33346
rect 15822 33294 15874 33346
rect 19406 33294 19458 33346
rect 13825 33238 13877 33290
rect 19630 33238 19682 33290
rect 19742 33266 19794 33318
rect 19966 33238 20018 33290
rect 20190 33266 20242 33318
rect 22094 33294 22146 33346
rect 22654 33266 22706 33318
rect 22878 33266 22930 33318
rect 23102 33238 23154 33290
rect 23214 33259 23266 33311
rect 26462 33294 26514 33346
rect 29710 33294 29762 33346
rect 33070 33294 33122 33346
rect 39454 33266 39506 33318
rect 39678 33294 39730 33346
rect 19238 33126 19290 33178
rect 20470 33182 20522 33234
rect 26854 33182 26906 33234
rect 40518 33238 40570 33290
rect 40686 33238 40738 33290
rect 40910 33255 40962 33307
rect 41806 33294 41858 33346
rect 42590 33259 42642 33311
rect 42758 33259 42810 33311
rect 42926 33238 42978 33290
rect 43150 33266 43202 33318
rect 44046 33294 44098 33346
rect 45950 33294 46002 33346
rect 48526 33294 48578 33346
rect 49310 33294 49362 33346
rect 41470 33182 41522 33234
rect 43430 33182 43482 33234
rect 45166 33238 45218 33290
rect 45390 33238 45442 33290
rect 45614 33238 45666 33290
rect 45726 33238 45778 33290
rect 21758 33070 21810 33122
rect 36374 33070 36426 33122
rect 40014 33070 40066 33122
rect 43878 33126 43930 33178
rect 44886 33182 44938 33234
rect 46118 33126 46170 33178
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 8766 32734 8818 32786
rect 25342 32734 25394 32786
rect 32566 32622 32618 32674
rect 33126 32622 33178 32674
rect 35142 32622 35194 32674
rect 5070 32510 5122 32562
rect 7086 32510 7138 32562
rect 7422 32525 7474 32577
rect 9102 32510 9154 32562
rect 9998 32510 10050 32562
rect 10782 32510 10834 32562
rect 13246 32525 13298 32577
rect 13582 32510 13634 32562
rect 14366 32537 14418 32589
rect 16270 32510 16322 32562
rect 17390 32510 17442 32562
rect 17726 32510 17778 32562
rect 18286 32510 18338 32562
rect 18510 32510 18562 32562
rect 19182 32510 19234 32562
rect 19406 32549 19458 32601
rect 19854 32510 19906 32562
rect 20190 32510 20242 32562
rect 20302 32510 20354 32562
rect 20862 32510 20914 32562
rect 21758 32510 21810 32562
rect 22542 32510 22594 32562
rect 25678 32510 25730 32562
rect 28702 32510 28754 32562
rect 29150 32510 29202 32562
rect 31054 32537 31106 32589
rect 31614 32510 31666 32562
rect 33350 32566 33402 32618
rect 33630 32538 33682 32590
rect 33854 32566 33906 32618
rect 33966 32566 34018 32618
rect 34302 32545 34354 32597
rect 34414 32566 34466 32618
rect 34638 32538 34690 32590
rect 34862 32566 34914 32618
rect 39006 32622 39058 32674
rect 35534 32510 35586 32562
rect 36318 32510 36370 32562
rect 37102 32510 37154 32562
rect 39454 32545 39506 32597
rect 39566 32538 39618 32590
rect 39846 32545 39898 32597
rect 40014 32566 40066 32618
rect 40294 32510 40346 32562
rect 40798 32510 40850 32562
rect 42030 32510 42082 32562
rect 42254 32510 42306 32562
rect 42702 32510 42754 32562
rect 42814 32510 42866 32562
rect 43000 32548 43052 32600
rect 44270 32510 44322 32562
rect 44606 32510 44658 32562
rect 45054 32510 45106 32562
rect 45278 32510 45330 32562
rect 45838 32537 45890 32589
rect 47966 32510 48018 32562
rect 48638 32510 48690 32562
rect 2382 32398 2434 32450
rect 4286 32398 4338 32450
rect 7534 32398 7586 32450
rect 9718 32398 9770 32450
rect 12686 32398 12738 32450
rect 13134 32398 13186 32450
rect 17278 32398 17330 32450
rect 19518 32398 19570 32450
rect 24446 32398 24498 32450
rect 26014 32398 26066 32450
rect 27918 32398 27970 32450
rect 43374 32398 43426 32450
rect 45166 32398 45218 32450
rect 20582 32286 20634 32338
rect 21198 32286 21250 32338
rect 31950 32286 32002 32338
rect 42254 32342 42306 32394
rect 41134 32286 41186 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 4622 31894 4674 31946
rect 11006 31950 11058 32002
rect 22934 31950 22986 32002
rect 3614 31838 3666 31890
rect 36262 31894 36314 31946
rect 38670 31950 38722 32002
rect 8542 31838 8594 31890
rect 9662 31838 9714 31890
rect 16606 31838 16658 31890
rect 20526 31838 20578 31890
rect 21422 31838 21474 31890
rect 24334 31838 24386 31890
rect 26574 31838 26626 31890
rect 27078 31838 27130 31890
rect 27862 31838 27914 31890
rect 29822 31838 29874 31890
rect 31726 31838 31778 31890
rect 32174 31838 32226 31890
rect 33854 31838 33906 31890
rect 45222 31894 45274 31946
rect 48862 31950 48914 32002
rect 40686 31838 40738 31890
rect 42590 31838 42642 31890
rect 3166 31726 3218 31778
rect 3502 31682 3554 31734
rect 4734 31726 4786 31778
rect 4958 31726 5010 31778
rect 5518 31726 5570 31778
rect 5742 31726 5794 31778
rect 9326 31726 9378 31778
rect 9774 31711 9826 31763
rect 10110 31726 10162 31778
rect 11249 31726 11301 31778
rect 12126 31726 12178 31778
rect 12798 31726 12850 31778
rect 13022 31726 13074 31778
rect 13358 31726 13410 31778
rect 13918 31670 13970 31722
rect 14030 31670 14082 31722
rect 14254 31698 14306 31750
rect 14478 31698 14530 31750
rect 17614 31698 17666 31750
rect 17838 31726 17890 31778
rect 18622 31726 18674 31778
rect 21982 31726 22034 31778
rect 22094 31726 22146 31778
rect 22654 31726 22706 31778
rect 6022 31614 6074 31666
rect 6638 31614 6690 31666
rect 12518 31614 12570 31666
rect 21814 31670 21866 31722
rect 23214 31698 23266 31750
rect 23438 31698 23490 31750
rect 23662 31698 23714 31750
rect 23774 31691 23826 31743
rect 24446 31682 24498 31734
rect 24782 31726 24834 31778
rect 25118 31691 25170 31743
rect 25286 31691 25338 31743
rect 25454 31698 25506 31750
rect 25678 31698 25730 31750
rect 25958 31726 26010 31778
rect 26238 31726 26290 31778
rect 27358 31726 27410 31778
rect 27582 31726 27634 31778
rect 28142 31726 28194 31778
rect 28366 31726 28418 31778
rect 29038 31726 29090 31778
rect 32286 31682 32338 31734
rect 32622 31726 32674 31778
rect 33070 31726 33122 31778
rect 36094 31726 36146 31778
rect 37326 31698 37378 31750
rect 39902 31726 39954 31778
rect 42926 31726 42978 31778
rect 44158 31726 44210 31778
rect 45390 31726 45442 31778
rect 47742 31726 47794 31778
rect 48526 31726 48578 31778
rect 49198 31726 49250 31778
rect 14758 31614 14810 31666
rect 10614 31502 10666 31554
rect 13526 31502 13578 31554
rect 22486 31558 22538 31610
rect 35758 31614 35810 31666
rect 45838 31614 45890 31666
rect 43262 31502 43314 31554
rect 43822 31502 43874 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 10390 31166 10442 31218
rect 11902 31166 11954 31218
rect 16606 31166 16658 31218
rect 5686 31054 5738 31106
rect 7310 31054 7362 31106
rect 12518 31054 12570 31106
rect 19126 31110 19178 31162
rect 30382 31166 30434 31218
rect 40294 31166 40346 31218
rect 46174 31166 46226 31218
rect 46790 31166 46842 31218
rect 47910 31166 47962 31218
rect 48974 31166 49026 31218
rect 28646 31054 28698 31106
rect 31558 31054 31610 31106
rect 1598 30942 1650 30994
rect 4958 30942 5010 30994
rect 5294 30942 5346 30994
rect 5406 30942 5458 30994
rect 5126 30886 5178 30938
rect 6190 30942 6242 30994
rect 7066 30942 7118 30994
rect 11006 30942 11058 30994
rect 12238 30942 12290 30994
rect 12742 30998 12794 31050
rect 13022 30970 13074 31022
rect 13246 30970 13298 31022
rect 13358 30977 13410 31029
rect 15598 30998 15650 31050
rect 15822 30998 15874 31050
rect 16046 30998 16098 31050
rect 13694 30942 13746 30994
rect 14030 30942 14082 30994
rect 14590 30942 14642 30994
rect 14814 30942 14866 30994
rect 16158 30977 16210 31029
rect 16942 30942 16994 30994
rect 18266 30998 18318 31050
rect 17390 30942 17442 30994
rect 18958 30942 19010 30994
rect 19406 30942 19458 30994
rect 19630 30942 19682 30994
rect 20302 30998 20354 31050
rect 20414 30998 20466 31050
rect 20638 30970 20690 31022
rect 20862 30998 20914 31050
rect 21142 30942 21194 30994
rect 22284 30979 22336 31031
rect 22430 30942 22482 30994
rect 22542 30942 22594 30994
rect 22766 30942 22818 30994
rect 22990 30942 23042 30994
rect 24110 30942 24162 30994
rect 24222 30942 24274 30994
rect 24558 30942 24610 30994
rect 25510 30977 25562 31029
rect 25790 30970 25842 31022
rect 25958 30977 26010 31029
rect 26126 30998 26178 31050
rect 26798 30942 26850 30994
rect 28926 30942 28978 30994
rect 29038 30942 29090 30994
rect 30718 30942 30770 30994
rect 31838 30998 31890 31050
rect 32062 30998 32114 31050
rect 31110 30942 31162 30994
rect 32286 30970 32338 31022
rect 32398 30998 32450 31050
rect 33630 30998 33682 31050
rect 34470 31054 34522 31106
rect 33742 30970 33794 31022
rect 34022 30998 34074 31050
rect 34190 30998 34242 31050
rect 38446 31054 38498 31106
rect 39734 31054 39786 31106
rect 34974 30942 35026 30994
rect 35198 30942 35250 30994
rect 38819 30998 38871 31050
rect 35758 30942 35810 30994
rect 36542 30942 36594 30994
rect 39006 30970 39058 31022
rect 39230 30970 39282 31022
rect 39454 30998 39506 31050
rect 42254 31054 42306 31106
rect 40462 30942 40514 30994
rect 40910 30977 40962 31029
rect 41022 30970 41074 31022
rect 41246 30970 41298 31022
rect 41508 30958 41560 31010
rect 42590 30942 42642 30994
rect 42814 30942 42866 30994
rect 43598 30942 43650 30994
rect 45838 30942 45890 30994
rect 47182 30942 47234 30994
rect 47406 30942 47458 30994
rect 47742 30942 47794 30994
rect 48638 30942 48690 30994
rect 2382 30830 2434 30882
rect 4286 30830 4338 30882
rect 15038 30830 15090 30882
rect 26630 30830 26682 30882
rect 27750 30830 27802 30882
rect 33238 30830 33290 30882
rect 45502 30830 45554 30882
rect 11342 30718 11394 30770
rect 15318 30718 15370 30770
rect 18510 30718 18562 30770
rect 19910 30718 19962 30770
rect 21870 30718 21922 30770
rect 23270 30718 23322 30770
rect 23774 30718 23826 30770
rect 25286 30718 25338 30770
rect 27134 30718 27186 30770
rect 35478 30718 35530 30770
rect 41750 30718 41802 30770
rect 47518 30774 47570 30826
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 2494 30382 2546 30434
rect 12406 30382 12458 30434
rect 20302 30326 20354 30378
rect 22150 30382 22202 30434
rect 32118 30382 32170 30434
rect 32734 30382 32786 30434
rect 44102 30382 44154 30434
rect 45670 30382 45722 30434
rect 4958 30270 5010 30322
rect 16382 30270 16434 30322
rect 18174 30270 18226 30322
rect 27918 30270 27970 30322
rect 38166 30270 38218 30322
rect 41918 30270 41970 30322
rect 2830 30158 2882 30210
rect 4062 30158 4114 30210
rect 4398 30158 4450 30210
rect 5070 30158 5122 30210
rect 5630 30158 5682 30210
rect 6302 30158 6354 30210
rect 6862 30158 6914 30210
rect 4734 30102 4786 30154
rect 5910 30102 5962 30154
rect 7198 30114 7250 30166
rect 7534 30158 7586 30210
rect 8318 30158 8370 30210
rect 9102 30158 9154 30210
rect 11006 30158 11058 30210
rect 11454 30158 11506 30210
rect 11678 30158 11730 30210
rect 12238 30158 12290 30210
rect 13918 30158 13970 30210
rect 14758 30123 14810 30175
rect 15038 30130 15090 30182
rect 15262 30102 15314 30154
rect 15374 30102 15426 30154
rect 15710 30158 15762 30210
rect 15822 30158 15874 30210
rect 15988 30158 16040 30210
rect 16942 30158 16994 30210
rect 17278 30131 17330 30183
rect 17614 30158 17666 30210
rect 18286 30114 18338 30166
rect 18622 30158 18674 30210
rect 18846 30158 18898 30210
rect 19070 30158 19122 30210
rect 19350 30158 19402 30210
rect 19910 30158 19962 30210
rect 20414 30158 20466 30210
rect 20750 30158 20802 30210
rect 11958 30046 12010 30098
rect 5742 29990 5794 30042
rect 7086 29990 7138 30042
rect 7870 29934 7922 29986
rect 14086 29990 14138 30042
rect 14534 30046 14586 30098
rect 21310 30102 21362 30154
rect 21422 30130 21474 30182
rect 21702 30123 21754 30175
rect 21926 30123 21978 30175
rect 22766 30158 22818 30210
rect 23550 30158 23602 30210
rect 26014 30158 26066 30210
rect 28702 30158 28754 30210
rect 31726 30158 31778 30210
rect 31838 30158 31890 30210
rect 32398 30158 32450 30210
rect 33070 30158 33122 30210
rect 33294 30158 33346 30210
rect 33574 30158 33626 30210
rect 33966 30158 34018 30210
rect 34638 30158 34690 30210
rect 35198 30158 35250 30210
rect 35870 30158 35922 30210
rect 34302 30102 34354 30154
rect 35534 30102 35586 30154
rect 37326 30123 37378 30175
rect 37438 30130 37490 30182
rect 37662 30102 37714 30154
rect 37886 30130 37938 30182
rect 38670 30158 38722 30210
rect 39006 30158 39058 30210
rect 39230 30158 39282 30210
rect 40014 30158 40066 30210
rect 42254 30158 42306 30210
rect 43262 30102 43314 30154
rect 43374 30102 43426 30154
rect 43598 30130 43650 30182
rect 43822 30130 43874 30182
rect 44830 30102 44882 30154
rect 44942 30102 44994 30154
rect 45166 30130 45218 30182
rect 45390 30130 45442 30182
rect 46398 30158 46450 30210
rect 47182 30158 47234 30210
rect 25454 30046 25506 30098
rect 17726 29990 17778 30042
rect 49086 30046 49138 30098
rect 34190 29990 34242 30042
rect 35310 29990 35362 30042
rect 42590 29934 42642 29986
rect 46230 29934 46282 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 9046 29598 9098 29650
rect 14982 29598 15034 29650
rect 4622 29486 4674 29538
rect 12686 29542 12738 29594
rect 15654 29598 15706 29650
rect 24446 29598 24498 29650
rect 22542 29542 22594 29594
rect 33574 29598 33626 29650
rect 35366 29598 35418 29650
rect 10446 29486 10498 29538
rect 24054 29486 24106 29538
rect 34078 29542 34130 29594
rect 40126 29598 40178 29650
rect 47014 29598 47066 29650
rect 1934 29374 1986 29426
rect 5294 29374 5346 29426
rect 7534 29401 7586 29453
rect 8206 29389 8258 29441
rect 8542 29374 8594 29426
rect 9662 29418 9714 29470
rect 10689 29430 10741 29482
rect 9998 29374 10050 29426
rect 11566 29374 11618 29426
rect 12126 29374 12178 29426
rect 12350 29413 12402 29465
rect 12798 29374 12850 29426
rect 15150 29374 15202 29426
rect 15766 29374 15818 29426
rect 15934 29374 15986 29426
rect 17278 29374 17330 29426
rect 19966 29374 20018 29426
rect 21086 29418 21138 29470
rect 26966 29486 27018 29538
rect 47854 29542 47906 29594
rect 21310 29374 21362 29426
rect 21982 29374 22034 29426
rect 22206 29413 22258 29465
rect 22654 29374 22706 29426
rect 22878 29374 22930 29426
rect 23102 29374 23154 29426
rect 24782 29374 24834 29426
rect 25342 29374 25394 29426
rect 26126 29430 26178 29482
rect 26238 29402 26290 29454
rect 26462 29430 26514 29482
rect 26686 29430 26738 29482
rect 27526 29374 27578 29426
rect 27806 29374 27858 29426
rect 28030 29374 28082 29426
rect 28142 29374 28194 29426
rect 31278 29374 31330 29426
rect 31390 29374 31442 29426
rect 33406 29374 33458 29426
rect 33966 29374 34018 29426
rect 34302 29401 34354 29453
rect 34638 29374 34690 29426
rect 35982 29401 36034 29453
rect 38558 29374 38610 29426
rect 38782 29374 38834 29426
rect 39454 29374 39506 29426
rect 40462 29374 40514 29426
rect 41078 29374 41130 29426
rect 41470 29401 41522 29453
rect 44382 29430 44434 29482
rect 44494 29430 44546 29482
rect 44718 29430 44770 29482
rect 44998 29430 45050 29482
rect 46454 29486 46506 29538
rect 45222 29374 45274 29426
rect 45502 29374 45554 29426
rect 47182 29374 47234 29426
rect 47406 29374 47458 29426
rect 48078 29374 48130 29426
rect 2718 29262 2770 29314
rect 8094 29262 8146 29314
rect 9550 29262 9602 29314
rect 18062 29262 18114 29314
rect 20974 29262 21026 29314
rect 28926 29262 28978 29314
rect 30830 29262 30882 29314
rect 38446 29206 38498 29258
rect 23382 29150 23434 29202
rect 25678 29150 25730 29202
rect 31670 29150 31722 29202
rect 39286 29150 39338 29202
rect 42814 29150 42866 29202
rect 45838 29150 45890 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 11398 28814 11450 28866
rect 16942 28814 16994 28866
rect 18398 28814 18450 28866
rect 19294 28814 19346 28866
rect 22598 28814 22650 28866
rect 24950 28814 25002 28866
rect 30326 28814 30378 28866
rect 33350 28814 33402 28866
rect 35366 28814 35418 28866
rect 3614 28702 3666 28754
rect 5742 28702 5794 28754
rect 7758 28702 7810 28754
rect 12126 28702 12178 28754
rect 25734 28702 25786 28754
rect 31838 28758 31890 28810
rect 43934 28814 43986 28866
rect 28534 28702 28586 28754
rect 32622 28702 32674 28754
rect 36038 28702 36090 28754
rect 37886 28702 37938 28754
rect 42254 28702 42306 28754
rect 44942 28702 44994 28754
rect 46846 28702 46898 28754
rect 2942 28590 2994 28642
rect 3110 28560 3162 28612
rect 3726 28575 3778 28627
rect 3950 28590 4002 28642
rect 4286 28590 4338 28642
rect 5966 28590 6018 28642
rect 5574 28534 5626 28586
rect 6302 28534 6354 28586
rect 6974 28590 7026 28642
rect 11678 28590 11730 28642
rect 11902 28590 11954 28642
rect 12238 28575 12290 28627
rect 12462 28590 12514 28642
rect 13358 28590 13410 28642
rect 13694 28590 13746 28642
rect 14814 28590 14866 28642
rect 15262 28590 15314 28642
rect 15934 28590 15986 28642
rect 14982 28534 15034 28586
rect 16270 28575 16322 28627
rect 17278 28590 17330 28642
rect 17390 28590 17442 28642
rect 18062 28590 18114 28642
rect 19630 28590 19682 28642
rect 9662 28478 9714 28530
rect 2942 28422 2994 28474
rect 15150 28478 15202 28530
rect 21254 28534 21306 28586
rect 21422 28534 21474 28586
rect 21646 28562 21698 28614
rect 21870 28562 21922 28614
rect 22430 28590 22482 28642
rect 25118 28590 25170 28642
rect 15542 28478 15594 28530
rect 26014 28534 26066 28586
rect 26238 28534 26290 28586
rect 26462 28562 26514 28614
rect 26574 28555 26626 28607
rect 26798 28590 26850 28642
rect 27134 28590 27186 28642
rect 27638 28590 27690 28642
rect 27918 28590 27970 28642
rect 28142 28590 28194 28642
rect 29486 28590 29538 28642
rect 29710 28590 29762 28642
rect 30606 28590 30658 28642
rect 30830 28590 30882 28642
rect 31054 28590 31106 28642
rect 31726 28590 31778 28642
rect 32174 28590 32226 28642
rect 32510 28546 32562 28598
rect 32846 28590 32898 28642
rect 33070 28590 33122 28642
rect 34302 28590 34354 28642
rect 34526 28551 34578 28603
rect 34974 28590 35026 28642
rect 35198 28590 35250 28642
rect 36486 28590 36538 28642
rect 37214 28590 37266 28642
rect 37550 28590 37602 28642
rect 37774 28551 37826 28603
rect 38222 28590 38274 28642
rect 38894 28590 38946 28642
rect 40798 28590 40850 28642
rect 41582 28590 41634 28642
rect 41918 28590 41970 28642
rect 42142 28575 42194 28627
rect 42534 28574 42586 28626
rect 42702 28562 42754 28614
rect 42926 28562 42978 28614
rect 43150 28562 43202 28614
rect 44270 28590 44322 28642
rect 47630 28590 47682 28642
rect 22150 28478 22202 28530
rect 29206 28478 29258 28530
rect 43430 28478 43482 28530
rect 16158 28422 16210 28474
rect 34190 28422 34242 28474
rect 17726 28366 17778 28418
rect 49254 28366 49306 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 7254 28030 7306 28082
rect 16886 28030 16938 28082
rect 29374 28030 29426 28082
rect 17614 27974 17666 28026
rect 20414 27974 20466 28026
rect 30046 28030 30098 28082
rect 32398 28030 32450 28082
rect 7870 27918 7922 27970
rect 31054 27974 31106 28026
rect 36150 28030 36202 28082
rect 36598 28030 36650 28082
rect 40238 28030 40290 28082
rect 37774 27974 37826 28026
rect 41078 28030 41130 28082
rect 42646 28030 42698 28082
rect 48974 28030 49026 28082
rect 1934 27806 1986 27858
rect 2158 27850 2210 27902
rect 2718 27806 2770 27858
rect 2961 27806 3013 27858
rect 3838 27806 3890 27858
rect 8113 27862 8165 27914
rect 4062 27806 4114 27858
rect 4846 27806 4898 27858
rect 6750 27806 6802 27858
rect 7086 27806 7138 27858
rect 8990 27806 9042 27858
rect 9494 27862 9546 27914
rect 22766 27918 22818 27970
rect 34246 27918 34298 27970
rect 45502 27918 45554 27970
rect 10222 27862 10274 27914
rect 9886 27806 9938 27858
rect 13246 27806 13298 27858
rect 14030 27806 14082 27858
rect 14814 27806 14866 27858
rect 14926 27806 14978 27858
rect 15072 27844 15124 27896
rect 15822 27806 15874 27858
rect 17838 27862 17890 27914
rect 16046 27806 16098 27858
rect 17502 27806 17554 27858
rect 18062 27806 18114 27858
rect 18902 27835 18954 27887
rect 19182 27806 19234 27858
rect 19630 27850 19682 27902
rect 19966 27806 20018 27858
rect 20526 27806 20578 27858
rect 20862 27833 20914 27885
rect 21198 27806 21250 27858
rect 21646 27839 21698 27891
rect 21982 27842 22034 27894
rect 22430 27842 22482 27894
rect 22586 27846 22638 27898
rect 23214 27806 23266 27858
rect 23438 27806 23490 27858
rect 25678 27833 25730 27885
rect 27918 27806 27970 27858
rect 28814 27806 28866 27858
rect 28926 27806 28978 27858
rect 29710 27806 29762 27858
rect 30382 27806 30434 27858
rect 31166 27806 31218 27858
rect 31838 27806 31890 27858
rect 32062 27806 32114 27858
rect 33406 27806 33458 27858
rect 33630 27806 33682 27858
rect 33742 27806 33794 27858
rect 33966 27806 34018 27858
rect 35086 27806 35138 27858
rect 36766 27806 36818 27858
rect 36990 27806 37042 27858
rect 37886 27806 37938 27858
rect 38110 27845 38162 27897
rect 38446 27806 38498 27858
rect 38894 27806 38946 27858
rect 39006 27806 39058 27858
rect 39152 27844 39204 27896
rect 39902 27806 39954 27858
rect 41358 27806 41410 27858
rect 42814 27806 42866 27858
rect 49310 27806 49362 27858
rect 2270 27694 2322 27746
rect 9662 27694 9714 27746
rect 11342 27694 11394 27746
rect 18734 27694 18786 27746
rect 19518 27694 19570 27746
rect 25398 27694 25450 27746
rect 43598 27694 43650 27746
rect 48246 27694 48298 27746
rect 23326 27638 23378 27690
rect 15486 27582 15538 27634
rect 16326 27582 16378 27634
rect 28534 27582 28586 27634
rect 33126 27582 33178 27634
rect 34750 27582 34802 27634
rect 37270 27582 37322 27634
rect 39566 27582 39618 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 4790 27190 4842 27242
rect 2382 27134 2434 27186
rect 4286 27134 4338 27186
rect 12854 27246 12906 27298
rect 14310 27246 14362 27298
rect 14870 27246 14922 27298
rect 21366 27246 21418 27298
rect 10278 27190 10330 27242
rect 22990 27246 23042 27298
rect 30774 27246 30826 27298
rect 38390 27246 38442 27298
rect 39398 27246 39450 27298
rect 48974 27246 49026 27298
rect 9774 27134 9826 27186
rect 11678 27134 11730 27186
rect 16270 27134 16322 27186
rect 17166 27134 17218 27186
rect 18342 27134 18394 27186
rect 24222 27134 24274 27186
rect 26126 27134 26178 27186
rect 32342 27134 32394 27186
rect 40798 27134 40850 27186
rect 41918 27134 41970 27186
rect 1598 27022 1650 27074
rect 4622 27022 4674 27074
rect 5630 27022 5682 27074
rect 6078 26983 6130 27035
rect 6302 27022 6354 27074
rect 7086 27022 7138 27074
rect 7870 27022 7922 27074
rect 10110 27022 10162 27074
rect 10670 27022 10722 27074
rect 11118 27022 11170 27074
rect 11454 27022 11506 27074
rect 11790 27022 11842 27074
rect 12462 27022 12514 27074
rect 12574 27022 12626 27074
rect 13470 26987 13522 27039
rect 13582 26966 13634 27018
rect 13806 26994 13858 27046
rect 14030 26994 14082 27046
rect 15150 27022 15202 27074
rect 15374 27022 15426 27074
rect 15598 27022 15650 27074
rect 15710 27022 15762 27074
rect 15878 27022 15930 27074
rect 17726 27022 17778 27074
rect 17838 27022 17890 27074
rect 18622 27022 18674 27074
rect 17558 26966 17610 27018
rect 18958 26995 19010 27047
rect 19294 27022 19346 27074
rect 20134 27022 20186 27074
rect 20414 27022 20466 27074
rect 20638 27022 20690 27074
rect 21534 27022 21586 27074
rect 21870 27022 21922 27074
rect 22746 27022 22798 27074
rect 26910 27022 26962 27074
rect 27022 27022 27074 27074
rect 27358 27022 27410 27074
rect 28086 27022 28138 27074
rect 28366 27022 28418 27074
rect 28590 27022 28642 27074
rect 29038 27022 29090 27074
rect 29710 27022 29762 27074
rect 31054 27022 31106 27074
rect 31278 27022 31330 27074
rect 31558 27022 31610 27074
rect 31838 27022 31890 27074
rect 31950 27022 32002 27074
rect 32622 27022 32674 27074
rect 32734 27022 32786 27074
rect 33518 27022 33570 27074
rect 33854 27022 33906 27074
rect 34078 27022 34130 27074
rect 34190 27022 34242 27074
rect 34470 27022 34522 27074
rect 34750 27022 34802 27074
rect 34974 27022 35026 27074
rect 35254 27022 35306 27074
rect 35534 27022 35586 27074
rect 37158 27022 37210 27074
rect 37886 27022 37938 27074
rect 38110 27022 38162 27074
rect 39006 27022 39058 27074
rect 39118 27022 39170 27074
rect 39678 27022 39730 27074
rect 40462 27022 40514 27074
rect 41134 27022 41186 27074
rect 44718 27022 44770 27074
rect 45502 27022 45554 27074
rect 47742 27022 47794 27074
rect 47966 27022 48018 27074
rect 49310 27022 49362 27074
rect 29374 26910 29426 26962
rect 6414 26854 6466 26906
rect 19406 26854 19458 26906
rect 36486 26910 36538 26962
rect 43822 26910 43874 26962
rect 47406 26910 47458 26962
rect 48246 26910 48298 26962
rect 30046 26798 30098 26850
rect 35870 26798 35922 26850
rect 37606 26798 37658 26850
rect 40014 26798 40066 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 10278 26462 10330 26514
rect 11958 26462 12010 26514
rect 13302 26462 13354 26514
rect 17614 26462 17666 26514
rect 27190 26462 27242 26514
rect 38390 26462 38442 26514
rect 42086 26462 42138 26514
rect 43598 26462 43650 26514
rect 44214 26462 44266 26514
rect 5686 26350 5738 26402
rect 2718 26238 2770 26290
rect 3054 26253 3106 26305
rect 5014 26238 5066 26290
rect 5182 26238 5234 26290
rect 5406 26238 5458 26290
rect 5966 26238 6018 26290
rect 6974 26282 7026 26334
rect 7198 26238 7250 26290
rect 8318 26282 8370 26334
rect 8654 26238 8706 26290
rect 9998 26238 10050 26290
rect 10110 26238 10162 26290
rect 10894 26238 10946 26290
rect 11118 26282 11170 26334
rect 13694 26294 13746 26346
rect 21758 26350 21810 26402
rect 26070 26350 26122 26402
rect 11790 26238 11842 26290
rect 12238 26238 12290 26290
rect 13470 26238 13522 26290
rect 13806 26266 13858 26318
rect 14086 26273 14138 26325
rect 14254 26266 14306 26318
rect 14534 26238 14586 26290
rect 14814 26238 14866 26290
rect 17278 26238 17330 26290
rect 17950 26238 18002 26290
rect 19070 26238 19122 26290
rect 22318 26238 22370 26290
rect 23058 26276 23110 26328
rect 24726 26238 24778 26290
rect 25230 26273 25282 26325
rect 25342 26294 25394 26346
rect 25622 26273 25674 26325
rect 25790 26294 25842 26346
rect 30270 26350 30322 26402
rect 32286 26350 32338 26402
rect 34638 26350 34690 26402
rect 26910 26238 26962 26290
rect 27022 26238 27074 26290
rect 27582 26238 27634 26290
rect 28366 26238 28418 26290
rect 31390 26238 31442 26290
rect 31726 26276 31778 26328
rect 35310 26350 35362 26402
rect 3166 26126 3218 26178
rect 6862 26126 6914 26178
rect 8206 26126 8258 26178
rect 11230 26126 11282 26178
rect 15766 26126 15818 26178
rect 16662 26126 16714 26178
rect 19854 26126 19906 26178
rect 24278 26126 24330 26178
rect 6302 26014 6354 26066
rect 9662 26014 9714 26066
rect 12574 26014 12626 26066
rect 15150 26014 15202 26066
rect 22542 26070 22594 26122
rect 31614 26182 31666 26234
rect 32454 26182 32506 26234
rect 33182 26238 33234 26290
rect 33294 26238 33346 26290
rect 34078 26276 34130 26328
rect 37214 26238 37266 26290
rect 37998 26238 38050 26290
rect 39118 26294 39170 26346
rect 40182 26350 40234 26402
rect 46118 26406 46170 26458
rect 39342 26294 39394 26346
rect 39454 26266 39506 26318
rect 39734 26273 39786 26325
rect 39902 26294 39954 26346
rect 33966 26182 34018 26234
rect 34806 26182 34858 26234
rect 41134 26238 41186 26290
rect 43262 26238 43314 26290
rect 45110 26294 45162 26346
rect 44942 26238 44994 26290
rect 45278 26238 45330 26290
rect 45390 26238 45442 26290
rect 46286 26238 46338 26290
rect 47630 26238 47682 26290
rect 47966 26276 48018 26328
rect 49198 26238 49250 26290
rect 30886 26126 30938 26178
rect 42534 26126 42586 26178
rect 47238 26182 47290 26234
rect 47406 26126 47458 26178
rect 18286 26014 18338 26066
rect 26574 26014 26626 26066
rect 31222 26014 31274 26066
rect 33574 26014 33626 26066
rect 38782 26014 38834 26066
rect 41470 26014 41522 26066
rect 45670 26014 45722 26066
rect 48862 26014 48914 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 11510 25678 11562 25730
rect 20302 25678 20354 25730
rect 21702 25678 21754 25730
rect 37438 25678 37490 25730
rect 38950 25678 39002 25730
rect 44886 25678 44938 25730
rect 3726 25566 3778 25618
rect 9102 25566 9154 25618
rect 11006 25566 11058 25618
rect 13918 25566 13970 25618
rect 15822 25566 15874 25618
rect 17726 25566 17778 25618
rect 19630 25566 19682 25618
rect 23438 25566 23490 25618
rect 25342 25566 25394 25618
rect 28254 25566 28306 25618
rect 29822 25566 29874 25618
rect 32790 25566 32842 25618
rect 40014 25566 40066 25618
rect 44326 25566 44378 25618
rect 46062 25566 46114 25618
rect 46622 25566 46674 25618
rect 48526 25566 48578 25618
rect 4510 25454 4562 25506
rect 5854 25454 5906 25506
rect 6190 25427 6242 25479
rect 6414 25454 6466 25506
rect 7982 25454 8034 25506
rect 8318 25454 8370 25506
rect 11790 25426 11842 25478
rect 12014 25398 12066 25450
rect 12238 25426 12290 25478
rect 12350 25398 12402 25450
rect 16606 25454 16658 25506
rect 16942 25454 16994 25506
rect 19966 25454 20018 25506
rect 21870 25454 21922 25506
rect 23102 25454 23154 25506
rect 26126 25454 26178 25506
rect 26350 25454 26402 25506
rect 27806 25426 27858 25478
rect 28030 25454 28082 25506
rect 1822 25342 1874 25394
rect 28422 25398 28474 25450
rect 29038 25454 29090 25506
rect 33854 25454 33906 25506
rect 34190 25416 34242 25468
rect 34526 25454 34578 25506
rect 34750 25454 34802 25506
rect 31726 25342 31778 25394
rect 34918 25398 34970 25450
rect 35086 25454 35138 25506
rect 35310 25454 35362 25506
rect 35590 25454 35642 25506
rect 35870 25454 35922 25506
rect 37774 25454 37826 25506
rect 38110 25419 38162 25471
rect 38222 25398 38274 25450
rect 38502 25419 38554 25471
rect 38670 25426 38722 25478
rect 39230 25454 39282 25506
rect 41918 25454 41970 25506
rect 42590 25454 42642 25506
rect 43466 25454 43518 25506
rect 44718 25454 44770 25506
rect 45838 25454 45890 25506
rect 45614 25398 45666 25450
rect 46230 25398 46282 25450
rect 49310 25454 49362 25506
rect 5966 25286 6018 25338
rect 43710 25342 43762 25394
rect 12854 25230 12906 25282
rect 22766 25230 22818 25282
rect 32342 25230 32394 25282
rect 33350 25230 33402 25282
rect 33686 25230 33738 25282
rect 36206 25230 36258 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 15262 24894 15314 24946
rect 29038 24894 29090 24946
rect 33182 24894 33234 24946
rect 34246 24894 34298 24946
rect 3950 24782 4002 24834
rect 4566 24782 4618 24834
rect 5406 24782 5458 24834
rect 35310 24782 35362 24834
rect 2830 24670 2882 24722
rect 3706 24670 3758 24722
rect 4846 24670 4898 24722
rect 5070 24670 5122 24722
rect 7310 24670 7362 24722
rect 8094 24670 8146 24722
rect 9102 24670 9154 24722
rect 10446 24726 10498 24778
rect 10670 24726 10722 24778
rect 10894 24726 10946 24778
rect 11006 24726 11058 24778
rect 10166 24670 10218 24722
rect 11230 24670 11282 24722
rect 12014 24670 12066 24722
rect 14478 24714 14530 24766
rect 14702 24670 14754 24722
rect 15598 24670 15650 24722
rect 16494 24670 16546 24722
rect 16606 24670 16658 24722
rect 17390 24670 17442 24722
rect 17726 24670 17778 24722
rect 18174 24670 18226 24722
rect 18286 24670 18338 24722
rect 21086 24697 21138 24749
rect 21758 24670 21810 24722
rect 22542 24670 22594 24722
rect 25118 24670 25170 24722
rect 25902 24670 25954 24722
rect 30718 24697 30770 24749
rect 31409 24726 31461 24778
rect 40294 24782 40346 24834
rect 32286 24670 32338 24722
rect 38502 24726 38554 24778
rect 39454 24726 39506 24778
rect 33518 24670 33570 24722
rect 34078 24670 34130 24722
rect 37214 24670 37266 24722
rect 37998 24670 38050 24722
rect 38222 24670 38274 24722
rect 39566 24698 39618 24750
rect 39846 24705 39898 24757
rect 40014 24726 40066 24778
rect 43822 24782 43874 24834
rect 49142 24782 49194 24834
rect 41134 24670 41186 24722
rect 41918 24670 41970 24722
rect 44270 24670 44322 24722
rect 44382 24670 44434 24722
rect 44568 24708 44620 24760
rect 45838 24670 45890 24722
rect 45950 24670 46002 24722
rect 46958 24670 47010 24722
rect 47294 24697 47346 24749
rect 47630 24670 47682 24722
rect 47966 24670 48018 24722
rect 48638 24670 48690 24722
rect 48862 24670 48914 24722
rect 13918 24558 13970 24610
rect 14366 24558 14418 24610
rect 24446 24558 24498 24610
rect 27806 24558 27858 24610
rect 33910 24558 33962 24610
rect 8766 24446 8818 24498
rect 17614 24502 17666 24554
rect 34918 24558 34970 24610
rect 38670 24558 38722 24610
rect 39174 24558 39226 24610
rect 45558 24558 45610 24610
rect 47070 24558 47122 24610
rect 16158 24446 16210 24498
rect 18566 24446 18618 24498
rect 20414 24446 20466 24498
rect 31166 24446 31218 24498
rect 44942 24446 44994 24498
rect 46230 24446 46282 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 12070 24110 12122 24162
rect 16998 24110 17050 24162
rect 23942 24110 23994 24162
rect 26854 24110 26906 24162
rect 28534 24110 28586 24162
rect 34974 24110 35026 24162
rect 35758 24110 35810 24162
rect 37102 24110 37154 24162
rect 37774 24110 37826 24162
rect 5966 23998 6018 24050
rect 8654 23998 8706 24050
rect 10558 23998 10610 24050
rect 13582 23998 13634 24050
rect 14646 23998 14698 24050
rect 15094 23998 15146 24050
rect 15542 23998 15594 24050
rect 15990 23998 16042 24050
rect 25734 23998 25786 24050
rect 34078 23998 34130 24050
rect 34582 23998 34634 24050
rect 40238 23998 40290 24050
rect 45502 23998 45554 24050
rect 1598 23886 1650 23938
rect 2382 23886 2434 23938
rect 5630 23886 5682 23938
rect 6078 23847 6130 23899
rect 6302 23886 6354 23938
rect 6638 23886 6690 23938
rect 7870 23886 7922 23938
rect 12350 23858 12402 23910
rect 12574 23858 12626 23910
rect 12798 23858 12850 23910
rect 4286 23774 4338 23826
rect 11734 23774 11786 23826
rect 12910 23830 12962 23882
rect 13918 23886 13970 23938
rect 16718 23886 16770 23938
rect 17278 23886 17330 23938
rect 17726 23886 17778 23938
rect 16382 23774 16434 23826
rect 17558 23830 17610 23882
rect 17950 23886 18002 23938
rect 18734 23886 18786 23938
rect 21758 23886 21810 23938
rect 22430 23886 22482 23938
rect 22673 23886 22725 23938
rect 23550 23886 23602 23938
rect 24222 23886 24274 23938
rect 24446 23886 24498 23938
rect 25958 23870 26010 23922
rect 17390 23774 17442 23826
rect 26126 23830 26178 23882
rect 26350 23830 26402 23882
rect 26574 23858 26626 23910
rect 27134 23886 27186 23938
rect 27358 23886 27410 23938
rect 28142 23886 28194 23938
rect 28254 23886 28306 23938
rect 29038 23886 29090 23938
rect 29822 23886 29874 23938
rect 32622 23886 32674 23938
rect 33294 23886 33346 23938
rect 33630 23886 33682 23938
rect 33910 23856 33962 23908
rect 35310 23886 35362 23938
rect 35422 23886 35474 23938
rect 37438 23886 37490 23938
rect 38110 23886 38162 23938
rect 20638 23774 20690 23826
rect 27638 23774 27690 23826
rect 31726 23774 31778 23826
rect 38334 23830 38386 23882
rect 38446 23858 38498 23910
rect 38670 23858 38722 23910
rect 39454 23886 39506 23938
rect 38894 23830 38946 23882
rect 42478 23886 42530 23938
rect 42702 23886 42754 23938
rect 42982 23886 43034 23938
rect 44046 23886 44098 23938
rect 44830 23886 44882 23938
rect 44942 23886 44994 23938
rect 45108 23886 45160 23938
rect 46734 23886 46786 23938
rect 46958 23886 47010 23938
rect 47630 23886 47682 23938
rect 39174 23774 39226 23826
rect 47406 23830 47458 23882
rect 48078 23886 48130 23938
rect 48302 23886 48354 23938
rect 48582 23886 48634 23938
rect 42142 23774 42194 23826
rect 21422 23662 21474 23714
rect 32286 23662 32338 23714
rect 32958 23662 33010 23714
rect 36374 23662 36426 23714
rect 43542 23662 43594 23714
rect 44214 23718 44266 23770
rect 47742 23718 47794 23770
rect 46398 23662 46450 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 2382 23326 2434 23378
rect 7870 23326 7922 23378
rect 3614 23270 3666 23322
rect 9662 23326 9714 23378
rect 13190 23326 13242 23378
rect 18790 23326 18842 23378
rect 19294 23326 19346 23378
rect 5350 23214 5402 23266
rect 11398 23214 11450 23266
rect 2718 23102 2770 23154
rect 3502 23102 3554 23154
rect 3838 23129 3890 23181
rect 4174 23102 4226 23154
rect 4846 23102 4898 23154
rect 5070 23102 5122 23154
rect 5742 23102 5794 23154
rect 6078 23117 6130 23169
rect 6862 23129 6914 23181
rect 9998 23102 10050 23154
rect 10838 23102 10890 23154
rect 11958 23137 12010 23189
rect 12238 23130 12290 23182
rect 12462 23130 12514 23182
rect 12574 23158 12626 23210
rect 13358 23102 13410 23154
rect 14590 23102 14642 23154
rect 15262 23102 15314 23154
rect 16494 23102 16546 23154
rect 17614 23158 17666 23210
rect 18174 23214 18226 23266
rect 20918 23270 20970 23322
rect 25398 23326 25450 23378
rect 34470 23326 34522 23378
rect 34918 23326 34970 23378
rect 38334 23326 38386 23378
rect 40406 23326 40458 23378
rect 44718 23214 44770 23266
rect 18342 23158 18394 23210
rect 18958 23102 19010 23154
rect 6190 22990 6242 23042
rect 10390 22990 10442 23042
rect 15094 22990 15146 23042
rect 17502 23046 17554 23098
rect 19910 23102 19962 23154
rect 21086 23102 21138 23154
rect 24782 23102 24834 23154
rect 25734 23102 25786 23154
rect 26014 23130 26066 23182
rect 26238 23158 26290 23210
rect 26406 23137 26458 23189
rect 26649 23158 26701 23210
rect 26798 23102 26850 23154
rect 27022 23102 27074 23154
rect 27806 23102 27858 23154
rect 28142 23146 28194 23198
rect 28702 23102 28754 23154
rect 29038 23102 29090 23154
rect 29598 23158 29650 23210
rect 29822 23158 29874 23210
rect 30046 23158 30098 23210
rect 30158 23158 30210 23210
rect 29318 23102 29370 23154
rect 31166 23102 31218 23154
rect 31278 23102 31330 23154
rect 31670 23102 31722 23154
rect 31950 23130 32002 23182
rect 32174 23158 32226 23210
rect 32398 23158 32450 23210
rect 32585 23158 32637 23210
rect 32958 23102 33010 23154
rect 33910 23102 33962 23154
rect 37998 23102 38050 23154
rect 38670 23102 38722 23154
rect 39006 23102 39058 23154
rect 41246 23129 41298 23181
rect 44550 23158 44602 23210
rect 48078 23214 48130 23266
rect 44046 23102 44098 23154
rect 44942 23102 44994 23154
rect 45390 23102 45442 23154
rect 48638 23102 48690 23154
rect 16886 22990 16938 23042
rect 21926 22990 21978 23042
rect 28254 22990 28306 23042
rect 35310 22990 35362 23042
rect 37214 22990 37266 23042
rect 39958 22990 40010 23042
rect 46174 22990 46226 23042
rect 48974 22990 49026 23042
rect 11734 22878 11786 22930
rect 13694 22878 13746 22930
rect 14254 22878 14306 22930
rect 15598 22878 15650 22930
rect 16158 22878 16210 22930
rect 24446 22878 24498 22930
rect 27302 22878 27354 22930
rect 30886 22878 30938 22930
rect 33294 22878 33346 22930
rect 39342 22878 39394 22930
rect 41918 22878 41970 22930
rect 43804 22878 43856 22930
rect 45110 22878 45162 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 3446 22542 3498 22594
rect 13526 22542 13578 22594
rect 37214 22542 37266 22594
rect 45950 22542 46002 22594
rect 4286 22430 4338 22482
rect 6638 22430 6690 22482
rect 15710 22430 15762 22482
rect 23998 22430 24050 22482
rect 25902 22430 25954 22482
rect 26854 22430 26906 22482
rect 29318 22430 29370 22482
rect 31166 22430 31218 22482
rect 33070 22430 33122 22482
rect 39006 22430 39058 22482
rect 40910 22430 40962 22482
rect 2270 22318 2322 22370
rect 2382 22318 2434 22370
rect 3054 22318 3106 22370
rect 3166 22318 3218 22370
rect 3950 22318 4002 22370
rect 4174 22274 4226 22326
rect 4958 22318 5010 22370
rect 5182 22318 5234 22370
rect 5854 22318 5906 22370
rect 8878 22318 8930 22370
rect 9662 22318 9714 22370
rect 11566 22318 11618 22370
rect 12350 22290 12402 22342
rect 2662 22206 2714 22258
rect 4678 22206 4730 22258
rect 8542 22206 8594 22258
rect 12574 22262 12626 22314
rect 12798 22290 12850 22342
rect 12910 22283 12962 22335
rect 13806 22262 13858 22314
rect 14030 22262 14082 22314
rect 14254 22290 14306 22342
rect 14366 22262 14418 22314
rect 14926 22318 14978 22370
rect 18510 22318 18562 22370
rect 18734 22318 18786 22370
rect 19014 22318 19066 22370
rect 19294 22318 19346 22370
rect 20862 22318 20914 22370
rect 21422 22318 21474 22370
rect 23214 22318 23266 22370
rect 27918 22290 27970 22342
rect 12070 22206 12122 22258
rect 17614 22206 17666 22258
rect 28142 22262 28194 22314
rect 28366 22262 28418 22314
rect 28478 22283 28530 22335
rect 29486 22318 29538 22370
rect 29710 22318 29762 22370
rect 33854 22318 33906 22370
rect 34414 22262 34466 22314
rect 34638 22290 34690 22342
rect 34862 22290 34914 22342
rect 34974 22283 35026 22335
rect 35254 22302 35306 22354
rect 35422 22290 35474 22342
rect 35646 22290 35698 22342
rect 36150 22318 36202 22370
rect 35870 22262 35922 22314
rect 36878 22318 36930 22370
rect 37550 22318 37602 22370
rect 38222 22318 38274 22370
rect 41470 22318 41522 22370
rect 42254 22318 42306 22370
rect 44830 22318 44882 22370
rect 45706 22287 45758 22339
rect 46734 22290 46786 22342
rect 48974 22318 49026 22370
rect 27638 22206 27690 22258
rect 29990 22206 30042 22258
rect 34134 22206 34186 22258
rect 44158 22206 44210 22258
rect 18230 22094 18282 22146
rect 19630 22094 19682 22146
rect 20526 22094 20578 22146
rect 21758 22094 21810 22146
rect 22486 22094 22538 22146
rect 30550 22094 30602 22146
rect 37886 22094 37938 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 9886 21758 9938 21810
rect 11398 21758 11450 21810
rect 37214 21758 37266 21810
rect 38558 21758 38610 21810
rect 39230 21758 39282 21810
rect 43262 21758 43314 21810
rect 44438 21758 44490 21810
rect 6414 21646 6466 21698
rect 15150 21646 15202 21698
rect 16550 21646 16602 21698
rect 1598 21534 1650 21586
rect 5294 21534 5346 21586
rect 5518 21534 5570 21586
rect 6657 21534 6709 21586
rect 7534 21534 7586 21586
rect 10222 21534 10274 21586
rect 15635 21590 15687 21642
rect 15822 21590 15874 21642
rect 16046 21590 16098 21642
rect 16270 21590 16322 21642
rect 46622 21702 46674 21754
rect 33406 21646 33458 21698
rect 10894 21534 10946 21586
rect 12014 21534 12066 21586
rect 12462 21534 12514 21586
rect 13246 21534 13298 21586
rect 17278 21534 17330 21586
rect 19854 21534 19906 21586
rect 20638 21534 20690 21586
rect 22878 21534 22930 21586
rect 23662 21534 23714 21586
rect 23998 21578 24050 21630
rect 24334 21534 24386 21586
rect 25678 21534 25730 21586
rect 26574 21534 26626 21586
rect 26966 21534 27018 21586
rect 31278 21590 31330 21642
rect 27806 21534 27858 21586
rect 30942 21534 30994 21586
rect 31614 21534 31666 21586
rect 36094 21534 36146 21586
rect 36206 21534 36258 21586
rect 37550 21534 37602 21586
rect 38222 21534 38274 21586
rect 38894 21534 38946 21586
rect 39566 21534 39618 21586
rect 39678 21534 39730 21586
rect 41134 21534 41186 21586
rect 41918 21534 41970 21586
rect 42366 21578 42418 21630
rect 42702 21534 42754 21586
rect 43598 21534 43650 21586
rect 44886 21534 44938 21586
rect 45278 21534 45330 21586
rect 45502 21578 45554 21630
rect 46174 21534 46226 21586
rect 46398 21573 46450 21625
rect 46846 21534 46898 21586
rect 47742 21549 47794 21601
rect 48078 21534 48130 21586
rect 48638 21534 48690 21586
rect 48862 21534 48914 21586
rect 2382 21422 2434 21474
rect 4286 21422 4338 21474
rect 11846 21422 11898 21474
rect 17950 21422 18002 21474
rect 20974 21422 21026 21474
rect 23886 21422 23938 21474
rect 28590 21422 28642 21474
rect 30494 21422 30546 21474
rect 31278 21422 31330 21474
rect 32566 21422 32618 21474
rect 35310 21422 35362 21474
rect 37886 21422 37938 21474
rect 42254 21422 42306 21474
rect 43990 21422 44042 21474
rect 45614 21422 45666 21474
rect 47350 21422 47402 21474
rect 47630 21422 47682 21474
rect 5798 21310 5850 21362
rect 10558 21310 10610 21362
rect 12182 21310 12234 21362
rect 17446 21310 17498 21362
rect 25342 21310 25394 21362
rect 26238 21310 26290 21362
rect 36542 21310 36594 21362
rect 40014 21310 40066 21362
rect 41302 21366 41354 21418
rect 41750 21310 41802 21362
rect 49142 21310 49194 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 2046 20974 2098 21026
rect 7086 20974 7138 21026
rect 7702 20974 7754 21026
rect 19518 20974 19570 21026
rect 14702 20918 14754 20970
rect 21366 20974 21418 21026
rect 22766 20974 22818 21026
rect 24110 20974 24162 21026
rect 24782 20974 24834 21026
rect 28366 20974 28418 21026
rect 2606 20862 2658 20914
rect 10110 20862 10162 20914
rect 20358 20862 20410 20914
rect 25902 20862 25954 20914
rect 27806 20862 27858 20914
rect 30550 20862 30602 20914
rect 32958 20918 33010 20970
rect 34302 20974 34354 21026
rect 34750 20862 34802 20914
rect 38782 20862 38834 20914
rect 43150 20862 43202 20914
rect 45054 20862 45106 20914
rect 2382 20750 2434 20802
rect 2718 20735 2770 20787
rect 3054 20750 3106 20802
rect 3390 20750 3442 20802
rect 3726 20723 3778 20775
rect 4062 20750 4114 20802
rect 4958 20750 5010 20802
rect 5182 20750 5234 20802
rect 6190 20750 6242 20802
rect 6470 20806 6522 20858
rect 6638 20750 6690 20802
rect 7422 20750 7474 20802
rect 7870 20750 7922 20802
rect 9326 20750 9378 20802
rect 12350 20750 12402 20802
rect 12574 20750 12626 20802
rect 13358 20750 13410 20802
rect 14590 20750 14642 20802
rect 15330 20712 15382 20764
rect 15934 20722 15986 20774
rect 17614 20750 17666 20802
rect 18398 20750 18450 20802
rect 19274 20750 19326 20802
rect 20862 20750 20914 20802
rect 21590 20715 21642 20767
rect 21870 20722 21922 20774
rect 22094 20722 22146 20774
rect 4678 20638 4730 20690
rect 5910 20638 5962 20690
rect 3502 20582 3554 20634
rect 6302 20638 6354 20690
rect 22206 20694 22258 20746
rect 22430 20750 22482 20802
rect 23102 20750 23154 20802
rect 23774 20750 23826 20802
rect 24446 20750 24498 20802
rect 25118 20750 25170 20802
rect 28702 20750 28754 20802
rect 29206 20750 29258 20802
rect 29486 20722 29538 20774
rect 29710 20722 29762 20774
rect 29934 20722 29986 20774
rect 33070 20750 33122 20802
rect 12014 20638 12066 20690
rect 12854 20638 12906 20690
rect 30046 20694 30098 20746
rect 31390 20694 31442 20746
rect 32062 20694 32114 20746
rect 32398 20694 32450 20746
rect 33746 20712 33798 20764
rect 33966 20750 34018 20802
rect 34862 20735 34914 20787
rect 35198 20750 35250 20802
rect 35422 20750 35474 20802
rect 37438 20750 37490 20802
rect 37998 20750 38050 20802
rect 41246 20711 41298 20763
rect 20694 20526 20746 20578
rect 23438 20526 23490 20578
rect 32622 20582 32674 20634
rect 40686 20638 40738 20690
rect 41750 20694 41802 20746
rect 42030 20694 42082 20746
rect 42254 20694 42306 20746
rect 42366 20715 42418 20767
rect 43393 20750 43445 20802
rect 44270 20750 44322 20802
rect 46958 20750 47010 20802
rect 47742 20750 47794 20802
rect 47966 20750 48018 20802
rect 48638 20750 48690 20802
rect 48302 20694 48354 20746
rect 35758 20526 35810 20578
rect 36374 20526 36426 20578
rect 37102 20526 37154 20578
rect 48078 20582 48130 20634
rect 37830 20526 37882 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 8822 20190 8874 20242
rect 5294 20134 5346 20186
rect 7198 20134 7250 20186
rect 23494 20190 23546 20242
rect 46062 20190 46114 20242
rect 20246 20078 20298 20130
rect 1598 19966 1650 20018
rect 4734 19966 4786 20018
rect 5070 19993 5122 20045
rect 6974 20022 7026 20074
rect 5406 19966 5458 20018
rect 5854 19966 5906 20018
rect 6638 19966 6690 20018
rect 7310 19966 7362 20018
rect 7758 20004 7810 20056
rect 8094 19966 8146 20018
rect 8486 19966 8538 20018
rect 8990 19966 9042 20018
rect 11510 19995 11562 20047
rect 12070 20022 12122 20074
rect 12294 20022 12346 20074
rect 12574 20022 12626 20074
rect 24054 20078 24106 20130
rect 11790 19966 11842 20018
rect 13470 19993 13522 20045
rect 16718 19966 16770 20018
rect 16830 19966 16882 20018
rect 17390 19966 17442 20018
rect 17726 19993 17778 20045
rect 18062 19966 18114 20018
rect 18734 19966 18786 20018
rect 18958 19966 19010 20018
rect 19294 19966 19346 20018
rect 21030 19966 21082 20018
rect 21870 19966 21922 20018
rect 22206 19966 22258 20018
rect 22542 19966 22594 20018
rect 24782 19966 24834 20018
rect 25230 19993 25282 20045
rect 27470 19966 27522 20018
rect 28366 19994 28418 20046
rect 28590 19994 28642 20046
rect 28814 20022 28866 20074
rect 28926 20022 28978 20074
rect 29486 20078 29538 20130
rect 33238 20078 33290 20130
rect 40014 20134 40066 20186
rect 30158 20022 30210 20074
rect 31502 20022 31554 20074
rect 34358 20078 34410 20130
rect 33518 20022 33570 20074
rect 33630 20022 33682 20074
rect 45334 20078 45386 20130
rect 29150 19966 29202 20018
rect 30382 19966 30434 20018
rect 2382 19854 2434 19906
rect 4286 19854 4338 19906
rect 6022 19798 6074 19850
rect 8318 19854 8370 19906
rect 11342 19854 11394 19906
rect 17614 19854 17666 19906
rect 13022 19742 13074 19794
rect 18622 19798 18674 19850
rect 21478 19854 21530 19906
rect 30606 19854 30658 19906
rect 30774 19910 30826 19962
rect 31278 19966 31330 20018
rect 31950 19966 32002 20018
rect 33854 19994 33906 20046
rect 34078 19994 34130 20046
rect 34638 19966 34690 20018
rect 34862 19966 34914 20018
rect 35142 19966 35194 20018
rect 35982 19993 36034 20045
rect 38558 19981 38610 20033
rect 38894 19966 38946 20018
rect 39566 19966 39618 20018
rect 39902 20005 39954 20057
rect 41190 20022 41242 20074
rect 40126 19966 40178 20018
rect 40910 19966 40962 20018
rect 41918 19966 41970 20018
rect 42254 19966 42306 20018
rect 42922 20004 42974 20056
rect 43598 19966 43650 20018
rect 44046 19966 44098 20018
rect 44158 19966 44210 20018
rect 44324 19966 44376 20018
rect 46398 19966 46450 20018
rect 46734 20010 46786 20062
rect 47070 19966 47122 20018
rect 47294 19966 47346 20018
rect 48638 19966 48690 20018
rect 48862 19966 48914 20018
rect 14478 19742 14530 19794
rect 16438 19742 16490 19794
rect 21870 19798 21922 19850
rect 31614 19854 31666 19906
rect 32454 19854 32506 19906
rect 38446 19854 38498 19906
rect 41358 19854 41410 19906
rect 42646 19854 42698 19906
rect 46622 19854 46674 19906
rect 19630 19742 19682 19794
rect 22878 19742 22930 19794
rect 24446 19742 24498 19794
rect 28086 19742 28138 19794
rect 36990 19742 37042 19794
rect 43710 19798 43762 19850
rect 44718 19742 44770 19794
rect 49142 19742 49194 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 2046 19406 2098 19458
rect 16998 19406 17050 19458
rect 24558 19406 24610 19458
rect 4062 19294 4114 19346
rect 5630 19294 5682 19346
rect 9326 19294 9378 19346
rect 10446 19294 10498 19346
rect 12350 19294 12402 19346
rect 12966 19294 13018 19346
rect 14590 19294 14642 19346
rect 31054 19350 31106 19402
rect 2382 19182 2434 19234
rect 4958 19154 5010 19206
rect 5742 19138 5794 19190
rect 5966 19182 6018 19234
rect 6638 19182 6690 19234
rect 7422 19182 7474 19234
rect 9662 19182 9714 19234
rect 13358 19182 13410 19234
rect 13918 19182 13970 19234
rect 14030 19182 14082 19234
rect 14196 19182 14248 19234
rect 15094 19182 15146 19234
rect 15318 19126 15370 19178
rect 15598 19126 15650 19178
rect 15822 19126 15874 19178
rect 15934 19126 15986 19178
rect 16270 19182 16322 19234
rect 16438 19238 16490 19290
rect 17782 19294 17834 19346
rect 20078 19294 20130 19346
rect 27582 19294 27634 19346
rect 28478 19294 28530 19346
rect 35758 19294 35810 19346
rect 37886 19294 37938 19346
rect 39790 19294 39842 19346
rect 45446 19294 45498 19346
rect 45894 19294 45946 19346
rect 49086 19294 49138 19346
rect 16718 19182 16770 19234
rect 20862 19182 20914 19234
rect 21198 19182 21250 19234
rect 21982 19182 22034 19234
rect 24222 19182 24274 19234
rect 24894 19182 24946 19234
rect 25678 19182 25730 19234
rect 28142 19182 28194 19234
rect 28310 19152 28362 19204
rect 29150 19147 29202 19199
rect 29262 19154 29314 19206
rect 29486 19154 29538 19206
rect 29710 19154 29762 19206
rect 30490 19144 30542 19196
rect 31166 19182 31218 19234
rect 36542 19182 36594 19234
rect 16606 19070 16658 19122
rect 18174 19070 18226 19122
rect 23886 19070 23938 19122
rect 31726 19126 31778 19178
rect 32174 19126 32226 19178
rect 32846 19126 32898 19178
rect 37102 19182 37154 19234
rect 40294 19182 40346 19234
rect 40574 19182 40626 19234
rect 40686 19182 40738 19234
rect 41022 19182 41074 19234
rect 41470 19182 41522 19234
rect 42254 19182 42306 19234
rect 46398 19182 46450 19234
rect 47182 19182 47234 19234
rect 29990 19070 30042 19122
rect 33854 19070 33906 19122
rect 32734 19014 32786 19066
rect 44158 19070 44210 19122
rect 13526 18958 13578 19010
rect 41190 18958 41242 19010
rect 44998 18958 45050 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 8094 18622 8146 18674
rect 4286 18566 4338 18618
rect 7422 18566 7474 18618
rect 19798 18622 19850 18674
rect 24054 18622 24106 18674
rect 26014 18622 26066 18674
rect 27302 18622 27354 18674
rect 43430 18622 43482 18674
rect 11678 18510 11730 18562
rect 17782 18510 17834 18562
rect 2046 18398 2098 18450
rect 3054 18398 3106 18450
rect 3502 18398 3554 18450
rect 3726 18442 3778 18494
rect 4734 18454 4786 18506
rect 4398 18398 4450 18450
rect 4958 18398 5010 18450
rect 5742 18398 5794 18450
rect 5854 18398 5906 18450
rect 6078 18398 6130 18450
rect 6638 18398 6690 18450
rect 7086 18437 7138 18489
rect 7310 18398 7362 18450
rect 7758 18398 7810 18450
rect 11921 18398 11973 18450
rect 12798 18398 12850 18450
rect 13358 18398 13410 18450
rect 13470 18398 13522 18450
rect 13750 18398 13802 18450
rect 14030 18398 14082 18450
rect 17278 18398 17330 18450
rect 17502 18398 17554 18450
rect 18398 18433 18450 18485
rect 18566 18454 18618 18506
rect 18790 18454 18842 18506
rect 19238 18510 19290 18562
rect 44046 18566 44098 18618
rect 47070 18622 47122 18674
rect 18958 18426 19010 18478
rect 20246 18398 20298 18450
rect 20750 18398 20802 18450
rect 21534 18398 21586 18450
rect 22274 18436 22326 18488
rect 22542 18398 22594 18450
rect 23214 18398 23266 18450
rect 24222 18398 24274 18450
rect 26350 18398 26402 18450
rect 28030 18398 28082 18450
rect 28142 18398 28194 18450
rect 30830 18398 30882 18450
rect 31614 18398 31666 18450
rect 31950 18425 32002 18477
rect 32286 18398 32338 18450
rect 33070 18454 33122 18506
rect 33238 18433 33290 18485
rect 33462 18454 33514 18506
rect 33630 18426 33682 18478
rect 33910 18398 33962 18450
rect 34526 18398 34578 18450
rect 36430 18398 36482 18450
rect 37214 18398 37266 18450
rect 37662 18398 37714 18450
rect 39902 18425 39954 18477
rect 41022 18398 41074 18450
rect 41246 18413 41298 18465
rect 41582 18398 41634 18450
rect 41806 18398 41858 18450
rect 42366 18398 42418 18450
rect 42590 18398 42642 18450
rect 43822 18398 43874 18450
rect 44046 18413 44098 18465
rect 44494 18398 44546 18450
rect 45370 18398 45422 18450
rect 45950 18398 46002 18450
rect 46174 18398 46226 18450
rect 46454 18398 46506 18450
rect 47406 18398 47458 18450
rect 47518 18398 47570 18450
rect 48806 18398 48858 18450
rect 49086 18398 49138 18450
rect 49198 18398 49250 18450
rect 3838 18286 3890 18338
rect 14814 18286 14866 18338
rect 16718 18286 16770 18338
rect 6246 18230 6298 18282
rect 2718 18174 2770 18226
rect 5462 18174 5514 18226
rect 24558 18286 24610 18338
rect 20918 18230 20970 18282
rect 21758 18230 21810 18282
rect 23326 18230 23378 18282
rect 27694 18286 27746 18338
rect 28926 18286 28978 18338
rect 31726 18286 31778 18338
rect 40406 18286 40458 18338
rect 41358 18286 41410 18338
rect 42086 18174 42138 18226
rect 42870 18174 42922 18226
rect 45614 18174 45666 18226
rect 47854 18174 47906 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 4846 17838 4898 17890
rect 7646 17838 7698 17890
rect 35030 17838 35082 17890
rect 42814 17838 42866 17890
rect 2382 17726 2434 17778
rect 7086 17726 7138 17778
rect 8990 17726 9042 17778
rect 11566 17726 11618 17778
rect 15822 17726 15874 17778
rect 19350 17726 19402 17778
rect 1598 17614 1650 17666
rect 4286 17614 4338 17666
rect 5182 17614 5234 17666
rect 6190 17614 6242 17666
rect 6302 17614 6354 17666
rect 6638 17614 6690 17666
rect 6974 17570 7026 17622
rect 7310 17614 7362 17666
rect 8318 17599 8370 17651
rect 8654 17614 8706 17666
rect 9102 17570 9154 17622
rect 9326 17614 9378 17666
rect 9942 17614 9994 17666
rect 11230 17614 11282 17666
rect 11454 17599 11506 17651
rect 11902 17614 11954 17666
rect 12238 17587 12290 17639
rect 12574 17614 12626 17666
rect 13358 17614 13410 17666
rect 15542 17670 15594 17722
rect 45502 17782 45554 17834
rect 26238 17726 26290 17778
rect 41022 17726 41074 17778
rect 43934 17726 43986 17778
rect 48526 17726 48578 17778
rect 13582 17614 13634 17666
rect 13862 17614 13914 17666
rect 15150 17614 15202 17666
rect 14814 17558 14866 17610
rect 15934 17570 15986 17622
rect 16158 17614 16210 17666
rect 16494 17614 16546 17666
rect 16718 17614 16770 17666
rect 17950 17614 18002 17666
rect 18398 17614 18450 17666
rect 5910 17502 5962 17554
rect 21310 17558 21362 17610
rect 15374 17502 15426 17554
rect 16998 17502 17050 17554
rect 21422 17558 21474 17610
rect 21982 17502 22034 17554
rect 22150 17558 22202 17610
rect 23102 17614 23154 17666
rect 23326 17614 23378 17666
rect 23774 17614 23826 17666
rect 24782 17614 24834 17666
rect 23494 17558 23546 17610
rect 25230 17586 25282 17638
rect 25454 17614 25506 17666
rect 25846 17614 25898 17666
rect 26798 17614 26850 17666
rect 26910 17614 26962 17666
rect 8430 17446 8482 17498
rect 12014 17446 12066 17498
rect 23662 17502 23714 17554
rect 24054 17502 24106 17554
rect 26632 17558 26684 17610
rect 27694 17614 27746 17666
rect 28086 17614 28138 17666
rect 31166 17614 31218 17666
rect 31950 17614 32002 17666
rect 32174 17586 32226 17638
rect 35310 17614 35362 17666
rect 35422 17614 35474 17666
rect 35646 17614 35698 17666
rect 36878 17614 36930 17666
rect 38222 17614 38274 17666
rect 38334 17614 38386 17666
rect 39118 17614 39170 17666
rect 41470 17614 41522 17666
rect 42142 17614 42194 17666
rect 25678 17502 25730 17554
rect 41750 17558 41802 17610
rect 43150 17614 43202 17666
rect 43486 17614 43538 17666
rect 43822 17599 43874 17651
rect 45278 17614 45330 17666
rect 45502 17614 45554 17666
rect 46622 17614 46674 17666
rect 49310 17614 49362 17666
rect 29262 17502 29314 17554
rect 17614 17390 17666 17442
rect 18734 17390 18786 17442
rect 22766 17390 22818 17442
rect 24614 17390 24666 17442
rect 27358 17390 27410 17442
rect 35982 17390 36034 17442
rect 41582 17446 41634 17498
rect 37886 17390 37938 17442
rect 46118 17390 46170 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 6134 17054 6186 17106
rect 5294 16998 5346 17050
rect 28590 17054 28642 17106
rect 36710 17054 36762 17106
rect 37158 17054 37210 17106
rect 37886 17054 37938 17106
rect 40126 17054 40178 17106
rect 48974 17054 49026 17106
rect 4286 16942 4338 16994
rect 8710 16942 8762 16994
rect 12798 16942 12850 16994
rect 1598 16830 1650 16882
rect 4846 16830 4898 16882
rect 5070 16857 5122 16909
rect 6862 16886 6914 16938
rect 13358 16942 13410 16994
rect 23438 16942 23490 16994
rect 5406 16830 5458 16882
rect 6414 16830 6466 16882
rect 7086 16830 7138 16882
rect 7422 16830 7474 16882
rect 8206 16830 8258 16882
rect 8430 16830 8482 16882
rect 9438 16830 9490 16882
rect 10110 16830 10162 16882
rect 16046 16830 16098 16882
rect 16382 16874 16434 16926
rect 16606 16830 16658 16882
rect 17838 16868 17890 16920
rect 33238 16942 33290 16994
rect 18174 16830 18226 16882
rect 2382 16718 2434 16770
rect 6750 16718 6802 16770
rect 10894 16718 10946 16770
rect 15262 16718 15314 16770
rect 16270 16718 16322 16770
rect 18398 16718 18450 16770
rect 18566 16774 18618 16826
rect 18846 16830 18898 16882
rect 18958 16830 19010 16882
rect 19104 16868 19156 16920
rect 20078 16830 20130 16882
rect 22766 16830 22818 16882
rect 24110 16886 24162 16938
rect 24726 16886 24778 16938
rect 26350 16886 26402 16938
rect 41078 16942 41130 16994
rect 46342 16942 46394 16994
rect 23102 16830 23154 16882
rect 24334 16830 24386 16882
rect 26574 16830 26626 16882
rect 26798 16830 26850 16882
rect 26966 16830 27018 16882
rect 27246 16830 27298 16882
rect 27358 16830 27410 16882
rect 27544 16868 27596 16920
rect 28926 16830 28978 16882
rect 29598 16830 29650 16882
rect 30382 16857 30434 16909
rect 33406 16830 33458 16882
rect 37550 16830 37602 16882
rect 38558 16845 38610 16897
rect 38894 16830 38946 16882
rect 39230 16830 39282 16882
rect 39342 16830 39394 16882
rect 40462 16830 40514 16882
rect 42366 16830 42418 16882
rect 42478 16830 42530 16882
rect 42702 16830 42754 16882
rect 42926 16830 42978 16882
rect 44046 16830 44098 16882
rect 44270 16830 44322 16882
rect 44550 16830 44602 16882
rect 45166 16830 45218 16882
rect 45278 16830 45330 16882
rect 45558 16830 45610 16882
rect 45950 16830 46002 16882
rect 46902 16859 46954 16911
rect 47070 16830 47122 16882
rect 49310 16830 49362 16882
rect 19518 16718 19570 16770
rect 20862 16718 20914 16770
rect 24558 16718 24610 16770
rect 27918 16718 27970 16770
rect 34190 16718 34242 16770
rect 36094 16718 36146 16770
rect 38446 16718 38498 16770
rect 41750 16718 41802 16770
rect 46062 16774 46114 16826
rect 46734 16718 46786 16770
rect 9774 16606 9826 16658
rect 29262 16606 29314 16658
rect 31054 16606 31106 16658
rect 39622 16606 39674 16658
rect 42086 16606 42138 16658
rect 43206 16606 43258 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 2494 16270 2546 16322
rect 5014 16270 5066 16322
rect 6134 16270 6186 16322
rect 11678 16270 11730 16322
rect 15038 16270 15090 16322
rect 16662 16270 16714 16322
rect 20134 16214 20186 16266
rect 20694 16270 20746 16322
rect 21534 16270 21586 16322
rect 3502 16158 3554 16210
rect 4286 16158 4338 16210
rect 8542 16158 8594 16210
rect 10446 16158 10498 16210
rect 19070 16158 19122 16210
rect 23326 16214 23378 16266
rect 25510 16270 25562 16322
rect 30158 16214 30210 16266
rect 27918 16158 27970 16210
rect 29598 16158 29650 16210
rect 36486 16158 36538 16210
rect 39566 16158 39618 16210
rect 41134 16158 41186 16210
rect 44214 16158 44266 16210
rect 44942 16158 44994 16210
rect 46846 16158 46898 16210
rect 49254 16158 49306 16210
rect 2830 16046 2882 16098
rect 3166 16046 3218 16098
rect 3390 16031 3442 16083
rect 3950 16046 4002 16098
rect 4118 16016 4170 16068
rect 4622 16046 4674 16098
rect 4734 16046 4786 16098
rect 5742 16046 5794 16098
rect 5854 16046 5906 16098
rect 6526 16046 6578 16098
rect 6694 16102 6746 16154
rect 6974 16046 7026 16098
rect 11230 16046 11282 16098
rect 12014 16046 12066 16098
rect 13918 16046 13970 16098
rect 14794 16046 14846 16098
rect 16494 16046 16546 16098
rect 17166 16046 17218 16098
rect 19854 16046 19906 16098
rect 19966 16025 20018 16077
rect 20862 16046 20914 16098
rect 22094 16046 22146 16098
rect 22206 16046 22258 16098
rect 22990 16046 23042 16098
rect 23214 16046 23266 16098
rect 23550 16046 23602 16098
rect 6862 15934 6914 15986
rect 21928 15990 21980 16042
rect 24222 16046 24274 16098
rect 24446 16046 24498 16098
rect 25342 16046 25394 16098
rect 28702 16046 28754 16098
rect 29262 16046 29314 16098
rect 29486 16002 29538 16054
rect 30046 16046 30098 16098
rect 30786 16008 30838 16060
rect 30942 16046 30994 16098
rect 31726 16046 31778 16098
rect 34526 16046 34578 16098
rect 35086 16046 35138 16098
rect 35758 16046 35810 16098
rect 7254 15934 7306 15986
rect 24726 15934 24778 15986
rect 26014 15934 26066 15986
rect 35534 15990 35586 16042
rect 36878 16046 36930 16098
rect 37662 16046 37714 16098
rect 39902 16046 39954 16098
rect 40238 16046 40290 16098
rect 43038 16046 43090 16098
rect 43822 16046 43874 16098
rect 47630 16046 47682 16098
rect 47742 16046 47794 16098
rect 33630 15934 33682 15986
rect 13638 15822 13690 15874
rect 23886 15822 23938 15874
rect 35646 15878 35698 15930
rect 34190 15822 34242 15874
rect 48078 15822 48130 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 9718 15486 9770 15538
rect 4622 15430 4674 15482
rect 20022 15486 20074 15538
rect 24502 15486 24554 15538
rect 23774 15430 23826 15482
rect 26406 15486 26458 15538
rect 16494 15374 16546 15426
rect 4790 15318 4842 15370
rect 2830 15262 2882 15314
rect 4510 15262 4562 15314
rect 5182 15262 5234 15314
rect 5966 15262 6018 15314
rect 6302 15306 6354 15358
rect 6974 15262 7026 15314
rect 7198 15262 7250 15314
rect 8038 15262 8090 15314
rect 9886 15282 9938 15334
rect 9998 15262 10050 15314
rect 11006 15289 11058 15341
rect 12238 15262 12290 15314
rect 17614 15318 17666 15370
rect 18230 15318 18282 15370
rect 30494 15374 30546 15426
rect 31390 15430 31442 15482
rect 37494 15486 37546 15538
rect 44718 15486 44770 15538
rect 39118 15430 39170 15482
rect 33126 15374 33178 15426
rect 36822 15374 36874 15426
rect 13806 15262 13858 15314
rect 17838 15262 17890 15314
rect 19220 15300 19272 15352
rect 19406 15262 19458 15314
rect 19518 15262 19570 15314
rect 20302 15289 20354 15341
rect 22542 15262 22594 15314
rect 23214 15262 23266 15314
rect 23662 15301 23714 15353
rect 23886 15262 23938 15314
rect 24334 15262 24386 15314
rect 25118 15262 25170 15314
rect 26238 15262 26290 15314
rect 27806 15262 27858 15314
rect 28590 15262 28642 15314
rect 31054 15262 31106 15314
rect 31502 15301 31554 15353
rect 31726 15262 31778 15314
rect 33406 15262 33458 15314
rect 33630 15262 33682 15314
rect 33966 15262 34018 15314
rect 34190 15262 34242 15314
rect 34918 15262 34970 15314
rect 35198 15262 35250 15314
rect 35422 15262 35474 15314
rect 35758 15277 35810 15329
rect 36094 15262 36146 15314
rect 36318 15262 36370 15314
rect 38782 15318 38834 15370
rect 36542 15262 36594 15314
rect 38334 15262 38386 15314
rect 39006 15262 39058 15314
rect 39566 15262 39618 15314
rect 39678 15262 39730 15314
rect 41918 15262 41970 15314
rect 42254 15277 42306 15329
rect 42814 15262 42866 15314
rect 43038 15262 43090 15314
rect 45726 15289 45778 15341
rect 46398 15262 46450 15314
rect 46734 15262 46786 15314
rect 47350 15262 47402 15314
rect 47742 15277 47794 15329
rect 48078 15262 48130 15314
rect 48638 15262 48690 15314
rect 6414 15150 6466 15202
rect 14590 15150 14642 15202
rect 18062 15150 18114 15202
rect 18846 15150 18898 15202
rect 35646 15150 35698 15202
rect 41638 15150 41690 15202
rect 42366 15150 42418 15202
rect 42702 15094 42754 15146
rect 2494 15038 2546 15090
rect 7478 15038 7530 15090
rect 25454 15038 25506 15090
rect 34470 15038 34522 15090
rect 39958 15038 40010 15090
rect 47630 15150 47682 15202
rect 46846 15094 46898 15146
rect 48974 15038 49026 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 30886 14702 30938 14754
rect 32622 14702 32674 14754
rect 42758 14702 42810 14754
rect 2382 14590 2434 14642
rect 4286 14590 4338 14642
rect 6414 14590 6466 14642
rect 7422 14590 7474 14642
rect 8542 14590 8594 14642
rect 10446 14590 10498 14642
rect 20078 14590 20130 14642
rect 24894 14590 24946 14642
rect 26798 14590 26850 14642
rect 31614 14590 31666 14642
rect 34190 14590 34242 14642
rect 36990 14590 37042 14642
rect 39790 14590 39842 14642
rect 47182 14590 47234 14642
rect 49086 14590 49138 14642
rect 1598 14478 1650 14530
rect 7590 14534 7642 14586
rect 5182 14478 5234 14530
rect 5966 14478 6018 14530
rect 6302 14463 6354 14515
rect 6974 14450 7026 14502
rect 7198 14478 7250 14530
rect 7758 14478 7810 14530
rect 11790 14478 11842 14530
rect 12126 14463 12178 14515
rect 12462 14478 12514 14530
rect 13470 14478 13522 14530
rect 14254 14478 14306 14530
rect 16606 14478 16658 14530
rect 17278 14478 17330 14530
rect 16942 14422 16994 14474
rect 18398 14478 18450 14530
rect 18622 14478 18674 14530
rect 19070 14450 19122 14502
rect 19294 14478 19346 14530
rect 19686 14478 19738 14530
rect 20472 14478 20524 14530
rect 20638 14478 20690 14530
rect 20750 14478 20802 14530
rect 21646 14450 21698 14502
rect 27582 14478 27634 14530
rect 29374 14478 29426 14530
rect 29710 14439 29762 14491
rect 29934 14478 29986 14530
rect 30494 14478 30546 14530
rect 30606 14478 30658 14530
rect 31726 14463 31778 14515
rect 31950 14478 32002 14530
rect 32286 14478 32338 14530
rect 33854 14478 33906 14530
rect 34078 14463 34130 14515
rect 35198 14478 35250 14530
rect 35646 14439 35698 14491
rect 35870 14478 35922 14530
rect 37102 14463 37154 14515
rect 37326 14478 37378 14530
rect 37662 14478 37714 14530
rect 38670 14478 38722 14530
rect 39230 14478 39282 14530
rect 41694 14478 41746 14530
rect 42478 14478 42530 14530
rect 39062 14422 39114 14474
rect 43038 14478 43090 14530
rect 43262 14478 43314 14530
rect 43374 14478 43426 14530
rect 46062 14478 46114 14530
rect 4846 14254 4898 14306
rect 11454 14254 11506 14306
rect 12126 14310 12178 14362
rect 16158 14366 16210 14418
rect 18118 14366 18170 14418
rect 19518 14366 19570 14418
rect 17390 14310 17442 14362
rect 45185 14422 45237 14474
rect 46398 14478 46450 14530
rect 44942 14366 44994 14418
rect 29822 14310 29874 14362
rect 35982 14310 36034 14362
rect 39230 14310 39282 14362
rect 37998 14254 38050 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 8038 13918 8090 13970
rect 7422 13862 7474 13914
rect 19070 13918 19122 13970
rect 9662 13862 9714 13914
rect 40238 13918 40290 13970
rect 13806 13806 13858 13858
rect 33742 13862 33794 13914
rect 41974 13918 42026 13970
rect 2606 13694 2658 13746
rect 5294 13694 5346 13746
rect 6078 13738 6130 13790
rect 7198 13750 7250 13802
rect 6414 13694 6466 13746
rect 6974 13694 7026 13746
rect 7534 13694 7586 13746
rect 7870 13694 7922 13746
rect 9102 13694 9154 13746
rect 9550 13694 9602 13746
rect 9886 13721 9938 13773
rect 10222 13694 10274 13746
rect 16494 13750 16546 13802
rect 22430 13806 22482 13858
rect 47406 13862 47458 13914
rect 35310 13806 35362 13858
rect 11118 13694 11170 13746
rect 11902 13694 11954 13746
rect 16606 13694 16658 13746
rect 17838 13694 17890 13746
rect 17950 13694 18002 13746
rect 18118 13694 18170 13746
rect 19406 13694 19458 13746
rect 19742 13694 19794 13746
rect 20526 13694 20578 13746
rect 22878 13727 22930 13779
rect 23214 13750 23266 13802
rect 23774 13750 23826 13802
rect 23972 13734 24024 13786
rect 25230 13694 25282 13746
rect 25342 13694 25394 13746
rect 25528 13732 25580 13784
rect 26798 13694 26850 13746
rect 34078 13750 34130 13802
rect 32622 13694 32674 13746
rect 33630 13694 33682 13746
rect 34302 13694 34354 13746
rect 37214 13694 37266 13746
rect 37998 13694 38050 13746
rect 38782 13694 38834 13746
rect 38894 13694 38946 13746
rect 39342 13738 39394 13790
rect 39678 13694 39730 13746
rect 39902 13694 39954 13746
rect 42142 13694 42194 13746
rect 42926 13694 42978 13746
rect 45950 13694 46002 13746
rect 46174 13694 46226 13746
rect 47182 13694 47234 13746
rect 47518 13721 47570 13773
rect 47854 13694 47906 13746
rect 48638 13694 48690 13746
rect 48862 13694 48914 13746
rect 3390 13582 3442 13634
rect 5966 13582 6018 13634
rect 23998 13582 24050 13634
rect 27582 13582 27634 13634
rect 29486 13582 29538 13634
rect 39230 13582 39282 13634
rect 43710 13582 43762 13634
rect 45614 13582 45666 13634
rect 49142 13582 49194 13634
rect 8766 13470 8818 13522
rect 16326 13470 16378 13522
rect 16774 13526 16826 13578
rect 18510 13470 18562 13522
rect 25902 13470 25954 13522
rect 32286 13470 32338 13522
rect 38502 13470 38554 13522
rect 42478 13470 42530 13522
rect 46454 13470 46506 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 3390 13134 3442 13186
rect 7814 13134 7866 13186
rect 21422 13134 21474 13186
rect 7310 13078 7362 13130
rect 23102 13134 23154 13186
rect 27918 13134 27970 13186
rect 2550 13022 2602 13074
rect 4622 13022 4674 13074
rect 9214 13022 9266 13074
rect 16382 13022 16434 13074
rect 18062 13022 18114 13074
rect 2718 12910 2770 12962
rect 3726 12910 3778 12962
rect 4398 12910 4450 12962
rect 5070 12910 5122 12962
rect 5630 12910 5682 12962
rect 4790 12854 4842 12906
rect 5966 12883 6018 12935
rect 6302 12910 6354 12962
rect 6974 12910 7026 12962
rect 7198 12910 7250 12962
rect 8094 12910 8146 12962
rect 8318 12910 8370 12962
rect 8430 12910 8482 12962
rect 11902 12910 11954 12962
rect 12126 12883 12178 12935
rect 12462 12910 12514 12962
rect 18230 12966 18282 13018
rect 19182 13022 19234 13074
rect 26742 13022 26794 13074
rect 30382 13022 30434 13074
rect 31838 13022 31890 13074
rect 33742 13022 33794 13074
rect 37774 13022 37826 13074
rect 39398 13022 39450 13074
rect 39902 13022 39954 13074
rect 43822 13022 43874 13074
rect 13694 12910 13746 12962
rect 14478 12910 14530 12962
rect 17502 12872 17554 12924
rect 17838 12910 17890 12962
rect 18510 12910 18562 12962
rect 18622 12910 18674 12962
rect 19966 12910 20018 12962
rect 18790 12854 18842 12906
rect 20302 12910 20354 12962
rect 21758 12910 21810 12962
rect 22430 12910 22482 12962
rect 22766 12910 22818 12962
rect 23438 12910 23490 12962
rect 24222 12910 24274 12962
rect 28254 12910 28306 12962
rect 28366 12910 28418 12962
rect 29374 12910 29426 12962
rect 29710 12883 29762 12935
rect 30046 12910 30098 12962
rect 30494 12895 30546 12947
rect 30718 12910 30770 12962
rect 31054 12910 31106 12962
rect 34190 12910 34242 12962
rect 34862 12910 34914 12962
rect 11118 12798 11170 12850
rect 5742 12742 5794 12794
rect 34470 12854 34522 12906
rect 35982 12910 36034 12962
rect 37326 12910 37378 12962
rect 37662 12866 37714 12918
rect 38334 12910 38386 12962
rect 38558 12910 38610 12962
rect 39566 12910 39618 12962
rect 41358 12910 41410 12962
rect 41694 12910 41746 12962
rect 41918 12895 41970 12947
rect 42254 12910 42306 12962
rect 42478 12910 42530 12962
rect 43598 12910 43650 12962
rect 43934 12895 43986 12947
rect 44270 12910 44322 12962
rect 45278 12910 45330 12962
rect 45502 12910 45554 12962
rect 45670 12966 45722 13018
rect 48526 12910 48578 12962
rect 49310 12910 49362 12962
rect 44942 12854 44994 12906
rect 26126 12798 26178 12850
rect 38838 12798 38890 12850
rect 12014 12742 12066 12794
rect 42758 12798 42810 12850
rect 46622 12798 46674 12850
rect 4062 12686 4114 12738
rect 29262 12742 29314 12794
rect 34302 12742 34354 12794
rect 22094 12686 22146 12738
rect 36318 12686 36370 12738
rect 40518 12686 40570 12738
rect 41022 12686 41074 12738
rect 41918 12742 41970 12794
rect 43262 12686 43314 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 6414 12350 6466 12402
rect 9718 12350 9770 12402
rect 26742 12350 26794 12402
rect 10222 12294 10274 12346
rect 32566 12350 32618 12402
rect 48974 12350 49026 12402
rect 13190 12238 13242 12290
rect 1598 12126 1650 12178
rect 4286 12126 4338 12178
rect 4958 12153 5010 12205
rect 7534 12126 7586 12178
rect 7646 12126 7698 12178
rect 8654 12126 8706 12178
rect 8878 12170 8930 12222
rect 10446 12126 10498 12178
rect 11006 12126 11058 12178
rect 11566 12126 11618 12178
rect 11902 12153 11954 12205
rect 12238 12126 12290 12178
rect 12798 12126 12850 12178
rect 12910 12126 12962 12178
rect 14030 12126 14082 12178
rect 17502 12182 17554 12234
rect 18062 12238 18114 12290
rect 21926 12238 21978 12290
rect 24446 12238 24498 12290
rect 18230 12182 18282 12234
rect 17838 12126 17890 12178
rect 18510 12126 18562 12178
rect 18622 12126 18674 12178
rect 18808 12163 18860 12215
rect 19574 12126 19626 12178
rect 20190 12154 20242 12206
rect 21310 12126 21362 12178
rect 2382 12014 2434 12066
rect 7926 12014 7978 12066
rect 8990 12014 9042 12066
rect 11678 12014 11730 12066
rect 14814 12014 14866 12066
rect 16718 12014 16770 12066
rect 19182 12014 19234 12066
rect 20414 12070 20466 12122
rect 21422 12126 21474 12178
rect 22934 12182 22986 12234
rect 23774 12182 23826 12234
rect 23998 12182 24050 12234
rect 27582 12238 27634 12290
rect 47854 12294 47906 12346
rect 45838 12238 45890 12290
rect 21646 12126 21698 12178
rect 23102 12126 23154 12178
rect 19742 12014 19794 12066
rect 23326 12014 23378 12066
rect 23494 12070 23546 12122
rect 24614 12070 24666 12122
rect 25454 12126 25506 12178
rect 25790 12126 25842 12178
rect 26126 12126 26178 12178
rect 26574 12126 26626 12178
rect 27246 12126 27298 12178
rect 28142 12126 28194 12178
rect 28366 12170 28418 12222
rect 29150 12153 29202 12205
rect 31502 12126 31554 12178
rect 31726 12126 31778 12178
rect 32006 12126 32058 12178
rect 32958 12126 33010 12178
rect 35982 12126 36034 12178
rect 36766 12126 36818 12178
rect 39006 12126 39058 12178
rect 39230 12126 39282 12178
rect 39790 12126 39842 12178
rect 42030 12126 42082 12178
rect 42142 12126 42194 12178
rect 42590 12170 42642 12222
rect 42814 12126 42866 12178
rect 43150 12126 43202 12178
rect 43934 12126 43986 12178
rect 46286 12126 46338 12178
rect 46622 12141 46674 12193
rect 47182 12126 47234 12178
rect 47406 12153 47458 12205
rect 47742 12126 47794 12178
rect 48638 12126 48690 12178
rect 28478 12014 28530 12066
rect 33742 12014 33794 12066
rect 35646 12014 35698 12066
rect 38670 12014 38722 12066
rect 41414 12014 41466 12066
rect 42478 12014 42530 12066
rect 46734 12014 46786 12066
rect 20974 11902 21026 11954
rect 26294 11902 26346 11954
rect 29822 11902 29874 11954
rect 39510 11902 39562 11954
rect 40126 11902 40178 11954
rect 41750 11902 41802 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 2382 11566 2434 11618
rect 18118 11566 18170 11618
rect 19742 11566 19794 11618
rect 21702 11566 21754 11618
rect 32622 11566 32674 11618
rect 34694 11566 34746 11618
rect 48246 11566 48298 11618
rect 7198 11510 7250 11562
rect 3502 11454 3554 11506
rect 5742 11454 5794 11506
rect 14254 11454 14306 11506
rect 15878 11454 15930 11506
rect 16326 11454 16378 11506
rect 18622 11454 18674 11506
rect 23550 11454 23602 11506
rect 25454 11454 25506 11506
rect 31726 11454 31778 11506
rect 40126 11454 40178 11506
rect 2718 11342 2770 11394
rect 3166 11342 3218 11394
rect 3390 11298 3442 11350
rect 4062 11342 4114 11394
rect 4286 11303 4338 11355
rect 4622 11342 4674 11394
rect 5630 11342 5682 11394
rect 6302 11342 6354 11394
rect 5966 11286 6018 11338
rect 6638 11342 6690 11394
rect 7310 11342 7362 11394
rect 7534 11342 7586 11394
rect 7870 11342 7922 11394
rect 8542 11342 8594 11394
rect 9326 11342 9378 11394
rect 11902 11342 11954 11394
rect 12350 11303 12402 11355
rect 12574 11342 12626 11394
rect 13806 11342 13858 11394
rect 13918 11342 13970 11394
rect 14366 11327 14418 11379
rect 14590 11342 14642 11394
rect 16830 11342 16882 11394
rect 16942 11342 16994 11394
rect 17614 11342 17666 11394
rect 17838 11342 17890 11394
rect 19016 11342 19068 11394
rect 19182 11342 19234 11394
rect 19294 11342 19346 11394
rect 20078 11342 20130 11394
rect 20414 11342 20466 11394
rect 20750 11342 20802 11394
rect 21982 11342 22034 11394
rect 22094 11342 22146 11394
rect 22766 11342 22818 11394
rect 25790 11342 25842 11394
rect 26574 11342 26626 11394
rect 29374 11342 29426 11394
rect 8206 11230 8258 11282
rect 3950 11174 4002 11226
rect 29598 11303 29650 11355
rect 30046 11342 30098 11394
rect 30494 11342 30546 11394
rect 30942 11303 30994 11355
rect 31166 11342 31218 11394
rect 31838 11327 31890 11379
rect 32174 11342 32226 11394
rect 32958 11342 33010 11394
rect 33630 11298 33682 11350
rect 33966 11342 34018 11394
rect 34302 11342 34354 11394
rect 34414 11342 34466 11394
rect 36318 11342 36370 11394
rect 36542 11342 36594 11394
rect 36878 11342 36930 11394
rect 40910 11342 40962 11394
rect 41022 11342 41074 11394
rect 41806 11342 41858 11394
rect 44718 11342 44770 11394
rect 45502 11342 45554 11394
rect 47854 11342 47906 11394
rect 47966 11342 48018 11394
rect 48526 11342 48578 11394
rect 11230 11230 11282 11282
rect 13526 11230 13578 11282
rect 28478 11230 28530 11282
rect 36038 11230 36090 11282
rect 38222 11230 38274 11282
rect 12014 11174 12066 11226
rect 16662 11118 16714 11170
rect 29262 11174 29314 11226
rect 31278 11174 31330 11226
rect 33854 11174 33906 11226
rect 43710 11230 43762 11282
rect 47406 11230 47458 11282
rect 17278 11118 17330 11170
rect 35254 11118 35306 11170
rect 35702 11118 35754 11170
rect 44326 11118 44378 11170
rect 48862 11118 48914 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 8094 10782 8146 10834
rect 8878 10782 8930 10834
rect 21142 10782 21194 10834
rect 9662 10726 9714 10778
rect 27806 10782 27858 10834
rect 4286 10670 4338 10722
rect 25342 10726 25394 10778
rect 34358 10782 34410 10834
rect 36766 10782 36818 10834
rect 39566 10726 39618 10778
rect 11230 10670 11282 10722
rect 1598 10558 1650 10610
rect 4790 10558 4842 10610
rect 5070 10558 5122 10610
rect 5294 10558 5346 10610
rect 5854 10558 5906 10610
rect 5966 10558 6018 10610
rect 6190 10558 6242 10610
rect 6414 10558 6466 10610
rect 7534 10558 7586 10610
rect 8430 10558 8482 10610
rect 8542 10558 8594 10610
rect 9774 10558 9826 10610
rect 10110 10585 10162 10637
rect 10446 10558 10498 10610
rect 13918 10558 13970 10610
rect 14030 10558 14082 10610
rect 17558 10614 17610 10666
rect 29094 10670 29146 10722
rect 33462 10670 33514 10722
rect 43038 10670 43090 10722
rect 18286 10614 18338 10666
rect 17950 10558 18002 10610
rect 18734 10558 18786 10610
rect 18846 10558 18898 10610
rect 19004 10608 19056 10660
rect 20340 10596 20392 10648
rect 20526 10558 20578 10610
rect 20638 10558 20690 10610
rect 21422 10558 21474 10610
rect 21534 10558 21586 10610
rect 21680 10596 21732 10648
rect 22486 10558 22538 10610
rect 22878 10558 22930 10610
rect 23102 10586 23154 10638
rect 24176 10608 24228 10660
rect 24334 10558 24386 10610
rect 24446 10558 24498 10610
rect 25678 10614 25730 10666
rect 25454 10558 25506 10610
rect 26126 10558 26178 10610
rect 26350 10558 26402 10610
rect 28142 10558 28194 10610
rect 28590 10558 28642 10610
rect 28814 10558 28866 10610
rect 29374 10558 29426 10610
rect 32062 10558 32114 10610
rect 32958 10558 33010 10610
rect 33182 10558 33234 10610
rect 34638 10558 34690 10610
rect 34974 10573 35026 10625
rect 35310 10558 35362 10610
rect 38446 10585 38498 10637
rect 39006 10558 39058 10610
rect 39342 10585 39394 10637
rect 39678 10558 39730 10610
rect 39902 10558 39954 10610
rect 41022 10573 41074 10625
rect 41246 10558 41298 10610
rect 42124 10558 42176 10610
rect 42366 10558 42418 10610
rect 2382 10446 2434 10498
rect 13134 10446 13186 10498
rect 14814 10446 14866 10498
rect 16718 10446 16770 10498
rect 17726 10446 17778 10498
rect 22094 10446 22146 10498
rect 22654 10446 22706 10498
rect 42870 10502 42922 10554
rect 43374 10558 43426 10610
rect 43934 10558 43986 10610
rect 44606 10602 44658 10654
rect 44942 10558 44994 10610
rect 47406 10585 47458 10637
rect 48246 10558 48298 10610
rect 48638 10558 48690 10610
rect 23774 10446 23826 10498
rect 30158 10446 30210 10498
rect 35086 10446 35138 10498
rect 40910 10446 40962 10498
rect 41582 10446 41634 10498
rect 41806 10446 41858 10498
rect 44494 10446 44546 10498
rect 5574 10334 5626 10386
rect 6694 10334 6746 10386
rect 7198 10334 7250 10386
rect 19406 10334 19458 10386
rect 19966 10334 20018 10386
rect 26518 10390 26570 10442
rect 35478 10334 35530 10386
rect 44158 10390 44210 10442
rect 40238 10334 40290 10386
rect 46062 10334 46114 10386
rect 48974 10334 49026 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 2382 9998 2434 10050
rect 30494 9998 30546 10050
rect 34862 9998 34914 10050
rect 36262 9998 36314 10050
rect 41470 9998 41522 10050
rect 12350 9886 12402 9938
rect 2718 9774 2770 9826
rect 3726 9774 3778 9826
rect 3950 9735 4002 9787
rect 4286 9774 4338 9826
rect 5630 9774 5682 9826
rect 6302 9774 6354 9826
rect 19686 9830 19738 9882
rect 21422 9886 21474 9938
rect 23662 9886 23714 9938
rect 25566 9886 25618 9938
rect 28142 9886 28194 9938
rect 37158 9886 37210 9938
rect 38334 9886 38386 9938
rect 40294 9886 40346 9938
rect 45502 9886 45554 9938
rect 47406 9886 47458 9938
rect 48638 9886 48690 9938
rect 6078 9718 6130 9770
rect 7310 9741 7362 9793
rect 7758 9718 7810 9770
rect 8094 9718 8146 9770
rect 8404 9741 8456 9793
rect 10782 9774 10834 9826
rect 11342 9774 11394 9826
rect 11902 9774 11954 9826
rect 12238 9759 12290 9811
rect 13582 9774 13634 9826
rect 14366 9774 14418 9826
rect 15150 9774 15202 9826
rect 17726 9774 17778 9826
rect 18286 9774 18338 9826
rect 8542 9662 8594 9714
rect 3614 9606 3666 9658
rect 6414 9606 6466 9658
rect 18062 9718 18114 9770
rect 18958 9736 19010 9788
rect 19294 9774 19346 9826
rect 20190 9746 20242 9798
rect 20414 9774 20466 9826
rect 20806 9774 20858 9826
rect 21814 9774 21866 9826
rect 21982 9774 22034 9826
rect 22094 9774 22146 9826
rect 22318 9774 22370 9826
rect 22878 9774 22930 9826
rect 27582 9774 27634 9826
rect 28254 9759 28306 9811
rect 28590 9774 28642 9826
rect 30830 9774 30882 9826
rect 31614 9774 31666 9826
rect 32490 9774 32542 9826
rect 17054 9662 17106 9714
rect 11566 9606 11618 9658
rect 19518 9662 19570 9714
rect 17838 9606 17890 9658
rect 20638 9662 20690 9714
rect 32734 9662 32786 9714
rect 33126 9718 33178 9770
rect 33294 9718 33346 9770
rect 33518 9735 33570 9787
rect 35254 9774 35306 9826
rect 35422 9774 35474 9826
rect 35534 9774 35586 9826
rect 35870 9774 35922 9826
rect 35982 9774 36034 9826
rect 37662 9774 37714 9826
rect 37998 9774 38050 9826
rect 38222 9735 38274 9787
rect 38670 9774 38722 9826
rect 39006 9774 39058 9826
rect 39342 9747 39394 9799
rect 39678 9774 39730 9826
rect 40574 9774 40626 9826
rect 41022 9774 41074 9826
rect 34078 9662 34130 9714
rect 40854 9718 40906 9770
rect 41806 9774 41858 9826
rect 41918 9774 41970 9826
rect 43318 9774 43370 9826
rect 43598 9774 43650 9826
rect 43822 9774 43874 9826
rect 48190 9774 48242 9826
rect 48302 9774 48354 9826
rect 40686 9662 40738 9714
rect 39118 9606 39170 9658
rect 27246 9550 27298 9602
rect 42254 9550 42306 9602
rect 42870 9550 42922 9602
rect 44214 9550 44266 9602
rect 44998 9550 45050 9602
rect 49142 9550 49194 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4902 9158 4954 9210
rect 6582 9214 6634 9266
rect 7086 9214 7138 9266
rect 10894 9102 10946 9154
rect 19406 9102 19458 9154
rect 19910 9158 19962 9210
rect 24726 9214 24778 9266
rect 1598 8990 1650 9042
rect 4286 8990 4338 9042
rect 4734 8990 4786 9042
rect 5820 9028 5872 9080
rect 5966 8990 6018 9042
rect 6078 8990 6130 9042
rect 7422 8990 7474 9042
rect 8206 8990 8258 9042
rect 8318 8990 8370 9042
rect 9998 8990 10050 9042
rect 12798 8990 12850 9042
rect 13582 8990 13634 9042
rect 18958 9046 19010 9098
rect 19574 9046 19626 9098
rect 28702 9102 28754 9154
rect 33406 9102 33458 9154
rect 38894 9102 38946 9154
rect 39510 9102 39562 9154
rect 43486 9102 43538 9154
rect 48134 9158 48186 9210
rect 14030 8990 14082 9042
rect 14814 8990 14866 9042
rect 17278 8990 17330 9042
rect 17950 8990 18002 9042
rect 19182 8990 19234 9042
rect 19742 8990 19794 9042
rect 20526 8990 20578 9042
rect 21310 8990 21362 9042
rect 24110 8990 24162 9042
rect 25118 8990 25170 9042
rect 26014 8990 26066 9042
rect 26798 8990 26850 9042
rect 29038 8990 29090 9042
rect 29262 8990 29314 9042
rect 30830 8990 30882 9042
rect 31502 9005 31554 9057
rect 31838 8990 31890 9042
rect 35310 8990 35362 9042
rect 36094 8990 36146 9042
rect 36206 8990 36258 9042
rect 39790 8990 39842 9042
rect 39902 8990 39954 9042
rect 40070 8990 40122 9042
rect 40238 8990 40290 9042
rect 44270 9046 44322 9098
rect 40798 8990 40850 9042
rect 41582 8990 41634 9042
rect 43990 8990 44042 9042
rect 44494 9018 44546 9070
rect 44718 9018 44770 9070
rect 44830 9025 44882 9077
rect 45614 9017 45666 9069
rect 48638 8990 48690 9042
rect 2382 8878 2434 8930
rect 16718 8878 16770 8930
rect 23214 8878 23266 8930
rect 31390 8878 31442 8930
rect 36990 8878 37042 8930
rect 5406 8766 5458 8818
rect 7870 8766 7922 8818
rect 8654 8766 8706 8818
rect 9662 8766 9714 8818
rect 17614 8766 17666 8818
rect 18118 8766 18170 8818
rect 23774 8766 23826 8818
rect 25454 8766 25506 8818
rect 29542 8766 29594 8818
rect 30494 8766 30546 8818
rect 48974 8766 49026 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 21926 8430 21978 8482
rect 23326 8430 23378 8482
rect 37214 8430 37266 8482
rect 39286 8430 39338 8482
rect 4958 8318 5010 8370
rect 5126 8262 5178 8314
rect 7254 8318 7306 8370
rect 12798 8318 12850 8370
rect 30046 8318 30098 8370
rect 36318 8318 36370 8370
rect 41134 8318 41186 8370
rect 43038 8318 43090 8370
rect 44326 8318 44378 8370
rect 3390 8178 3442 8230
rect 3614 8206 3666 8258
rect 3838 8094 3890 8146
rect 4006 8150 4058 8202
rect 4398 8168 4450 8220
rect 4734 8206 4786 8258
rect 5630 8206 5682 8258
rect 6302 8206 6354 8258
rect 6078 8150 6130 8202
rect 7422 8206 7474 8258
rect 8206 8206 8258 8258
rect 10558 8206 10610 8258
rect 11230 8206 11282 8258
rect 12350 8206 12402 8258
rect 12462 8206 12514 8258
rect 13918 8206 13970 8258
rect 10894 8150 10946 8202
rect 16158 8178 16210 8230
rect 18622 8178 18674 8230
rect 19854 8206 19906 8258
rect 20078 8206 20130 8258
rect 20190 8206 20242 8258
rect 21590 8206 21642 8258
rect 22094 8206 22146 8258
rect 22318 8178 22370 8230
rect 25006 8206 25058 8258
rect 25230 8206 25282 8258
rect 26574 8206 26626 8258
rect 26966 8206 27018 8258
rect 27470 8206 27522 8258
rect 28030 8206 28082 8258
rect 29262 8206 29314 8258
rect 27806 8150 27858 8202
rect 32398 8206 32450 8258
rect 33274 8206 33326 8258
rect 33854 8206 33906 8258
rect 34918 8206 34970 8258
rect 35646 8206 35698 8258
rect 35870 8206 35922 8258
rect 36150 8176 36202 8228
rect 37550 8206 37602 8258
rect 37774 8206 37826 8258
rect 38110 8206 38162 8258
rect 38222 8206 38274 8258
rect 10110 8094 10162 8146
rect 19574 8094 19626 8146
rect 25510 8094 25562 8146
rect 31950 8094 32002 8146
rect 6190 8038 6242 8090
rect 10670 8038 10722 8090
rect 12182 7982 12234 8034
rect 17614 7982 17666 8034
rect 20526 7982 20578 8034
rect 27918 8038 27970 8090
rect 37942 8150 37994 8202
rect 38502 8206 38554 8258
rect 38894 8206 38946 8258
rect 39006 8206 39058 8258
rect 39566 8206 39618 8258
rect 39790 8206 39842 8258
rect 40350 8206 40402 8258
rect 43374 8206 43426 8258
rect 45166 8150 45218 8202
rect 45278 8178 45330 8230
rect 48526 8206 48578 8258
rect 49310 8206 49362 8258
rect 45502 8150 45554 8202
rect 45749 8150 45801 8202
rect 33518 8094 33570 8146
rect 40070 8094 40122 8146
rect 46006 8094 46058 8146
rect 46622 8094 46674 8146
rect 26238 7982 26290 8034
rect 34190 7982 34242 8034
rect 35310 7982 35362 8034
rect 43710 7982 43762 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 5854 7646 5906 7698
rect 7590 7646 7642 7698
rect 48974 7646 49026 7698
rect 11006 7590 11058 7642
rect 1598 7422 1650 7474
rect 7198 7449 7250 7501
rect 7982 7478 8034 7530
rect 8654 7534 8706 7586
rect 7758 7422 7810 7474
rect 11846 7534 11898 7586
rect 12294 7534 12346 7586
rect 20302 7534 20354 7586
rect 8094 7460 8146 7512
rect 9662 7422 9714 7474
rect 9998 7437 10050 7489
rect 10446 7422 10498 7474
rect 10782 7449 10834 7501
rect 11118 7422 11170 7474
rect 8822 7366 8874 7418
rect 13450 7478 13502 7530
rect 24446 7534 24498 7586
rect 31166 7590 31218 7642
rect 29262 7534 29314 7586
rect 38558 7534 38610 7586
rect 12574 7422 12626 7474
rect 14030 7422 14082 7474
rect 14814 7422 14866 7474
rect 17614 7422 17666 7474
rect 18398 7422 18450 7474
rect 20862 7437 20914 7489
rect 21086 7422 21138 7474
rect 21758 7422 21810 7474
rect 25118 7422 25170 7474
rect 25902 7422 25954 7474
rect 27806 7422 27858 7474
rect 28142 7422 28194 7474
rect 28366 7422 28418 7474
rect 28926 7422 28978 7474
rect 30718 7422 30770 7474
rect 31054 7449 31106 7501
rect 31278 7422 31330 7474
rect 31782 7422 31834 7474
rect 32062 7422 32114 7474
rect 32174 7422 32226 7474
rect 34862 7422 34914 7474
rect 34974 7422 35026 7474
rect 35198 7422 35250 7474
rect 35422 7422 35474 7474
rect 35702 7422 35754 7474
rect 36206 7422 36258 7474
rect 36542 7422 36594 7474
rect 37438 7422 37490 7474
rect 38314 7422 38366 7474
rect 39454 7422 39506 7474
rect 41134 7422 41186 7474
rect 43038 7449 43090 7501
rect 43598 7422 43650 7474
rect 44774 7457 44826 7509
rect 45054 7450 45106 7502
rect 45278 7478 45330 7530
rect 45465 7478 45517 7530
rect 45726 7449 45778 7501
rect 48638 7422 48690 7474
rect 2382 7310 2434 7362
rect 4286 7310 4338 7362
rect 10110 7310 10162 7362
rect 16718 7310 16770 7362
rect 20750 7310 20802 7362
rect 22542 7310 22594 7362
rect 33238 7310 33290 7362
rect 33686 7310 33738 7362
rect 34246 7310 34298 7362
rect 36094 7254 36146 7306
rect 37046 7310 37098 7362
rect 39174 7310 39226 7362
rect 13694 7198 13746 7250
rect 28646 7198 28698 7250
rect 34582 7198 34634 7250
rect 43934 7198 43986 7250
rect 44550 7198 44602 7250
rect 47070 7198 47122 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 2494 6862 2546 6914
rect 23102 6862 23154 6914
rect 37158 6862 37210 6914
rect 37942 6862 37994 6914
rect 5070 6750 5122 6802
rect 7758 6750 7810 6802
rect 9774 6750 9826 6802
rect 12238 6750 12290 6802
rect 14142 6750 14194 6802
rect 25454 6750 25506 6802
rect 27470 6750 27522 6802
rect 30270 6750 30322 6802
rect 33182 6750 33234 6802
rect 40462 6750 40514 6802
rect 2830 6638 2882 6690
rect 3726 6638 3778 6690
rect 4622 6638 4674 6690
rect 4958 6623 5010 6675
rect 5630 6638 5682 6690
rect 6302 6638 6354 6690
rect 7086 6638 7138 6690
rect 7422 6638 7474 6690
rect 8094 6638 8146 6690
rect 5966 6582 6018 6634
rect 7758 6582 7810 6634
rect 8654 6605 8706 6657
rect 8990 6582 9042 6634
rect 9438 6582 9490 6634
rect 9748 6598 9800 6650
rect 13022 6638 13074 6690
rect 13358 6638 13410 6690
rect 16606 6638 16658 6690
rect 17166 6638 17218 6690
rect 5742 6470 5794 6522
rect 6918 6470 6970 6522
rect 10334 6526 10386 6578
rect 16942 6582 16994 6634
rect 17614 6638 17666 6690
rect 17838 6638 17890 6690
rect 18398 6638 18450 6690
rect 19070 6638 19122 6690
rect 19406 6599 19458 6651
rect 19630 6638 19682 6690
rect 20078 6638 20130 6690
rect 20302 6638 20354 6690
rect 21198 6638 21250 6690
rect 22430 6638 22482 6690
rect 23438 6638 23490 6690
rect 23998 6638 24050 6690
rect 24334 6611 24386 6663
rect 24558 6638 24610 6690
rect 25006 6638 25058 6690
rect 25342 6623 25394 6675
rect 25958 6638 26010 6690
rect 26462 6638 26514 6690
rect 26798 6611 26850 6663
rect 27134 6638 27186 6690
rect 27582 6623 27634 6675
rect 27918 6638 27970 6690
rect 29598 6638 29650 6690
rect 29934 6638 29986 6690
rect 30158 6594 30210 6646
rect 30494 6638 30546 6690
rect 30718 6638 30770 6690
rect 31838 6638 31890 6690
rect 32342 6638 32394 6690
rect 32622 6638 32674 6690
rect 32846 6638 32898 6690
rect 35086 6638 35138 6690
rect 35870 6638 35922 6690
rect 36542 6638 36594 6690
rect 37326 6638 37378 6690
rect 37550 6638 37602 6690
rect 37662 6638 37714 6690
rect 38558 6638 38610 6690
rect 41246 6638 41298 6690
rect 41358 6638 41410 6690
rect 41694 6638 41746 6690
rect 42590 6638 42642 6690
rect 43150 6610 43202 6662
rect 43374 6582 43426 6634
rect 43598 6582 43650 6634
rect 43710 6582 43762 6634
rect 16046 6526 16098 6578
rect 18118 6526 18170 6578
rect 20582 6526 20634 6578
rect 30998 6526 31050 6578
rect 42870 6526 42922 6578
rect 17278 6470 17330 6522
rect 18566 6470 18618 6522
rect 19518 6470 19570 6522
rect 21534 6414 21586 6466
rect 23886 6470 23938 6522
rect 26350 6470 26402 6522
rect 44886 6526 44938 6578
rect 45110 6582 45162 6634
rect 45390 6582 45442 6634
rect 45558 6603 45610 6655
rect 48526 6638 48578 6690
rect 49310 6638 49362 6690
rect 45726 6582 45778 6634
rect 46622 6526 46674 6578
rect 22094 6414 22146 6466
rect 29262 6414 29314 6466
rect 31502 6414 31554 6466
rect 36206 6414 36258 6466
rect 42254 6414 42306 6466
rect 44214 6414 44266 6466
rect 46118 6414 46170 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 11454 6078 11506 6130
rect 5070 6022 5122 6074
rect 18342 6078 18394 6130
rect 18734 6078 18786 6130
rect 25398 6078 25450 6130
rect 25846 6078 25898 6130
rect 26518 6078 26570 6130
rect 6582 5966 6634 6018
rect 8430 5966 8482 6018
rect 5238 5910 5290 5962
rect 4734 5854 4786 5906
rect 4958 5854 5010 5906
rect 5630 5854 5682 5906
rect 6078 5854 6130 5906
rect 6302 5854 6354 5906
rect 6974 5854 7026 5906
rect 7310 5854 7362 5906
rect 7422 5854 7474 5906
rect 7142 5798 7194 5850
rect 8262 5910 8314 5962
rect 8822 5966 8874 6018
rect 30382 6022 30434 6074
rect 31726 6022 31778 6074
rect 29822 5966 29874 6018
rect 8094 5854 8146 5906
rect 8542 5854 8594 5906
rect 9998 5854 10050 5906
rect 10334 5854 10386 5906
rect 11118 5854 11170 5906
rect 15374 5854 15426 5906
rect 15710 5854 15762 5906
rect 15934 5869 15986 5921
rect 16382 5854 16434 5906
rect 16494 5854 16546 5906
rect 17502 5869 17554 5921
rect 17726 5854 17778 5906
rect 19070 5854 19122 5906
rect 19294 5881 19346 5933
rect 22188 5854 22240 5906
rect 22934 5910 22986 5962
rect 22430 5854 22482 5906
rect 23102 5854 23154 5906
rect 24446 5854 24498 5906
rect 24558 5854 24610 5906
rect 30550 5910 30602 5962
rect 27134 5854 27186 5906
rect 27918 5854 27970 5906
rect 30270 5854 30322 5906
rect 30942 5854 30994 5906
rect 31614 5854 31666 5906
rect 32062 5893 32114 5945
rect 32286 5854 32338 5906
rect 33126 5854 33178 5906
rect 33406 5854 33458 5906
rect 33518 5854 33570 5906
rect 33854 5854 33906 5906
rect 34190 5869 34242 5921
rect 34750 5854 34802 5906
rect 34974 5898 35026 5950
rect 35646 5854 35698 5906
rect 37886 5881 37938 5933
rect 38558 5910 38610 5962
rect 39118 5966 39170 6018
rect 43598 5966 43650 6018
rect 44102 5966 44154 6018
rect 44382 5910 44434 5962
rect 44606 5910 44658 5962
rect 38894 5854 38946 5906
rect 39678 5854 39730 5906
rect 39902 5854 39954 5906
rect 40910 5854 40962 5906
rect 44830 5882 44882 5934
rect 44942 5889 44994 5941
rect 47518 5854 47570 5906
rect 48302 5854 48354 5906
rect 48638 5854 48690 5906
rect 39286 5798 39338 5850
rect 16046 5742 16098 5794
rect 17390 5742 17442 5794
rect 23606 5742 23658 5794
rect 34302 5742 34354 5794
rect 35086 5742 35138 5794
rect 4398 5630 4450 5682
rect 10110 5686 10162 5738
rect 41694 5742 41746 5794
rect 45614 5742 45666 5794
rect 7702 5630 7754 5682
rect 39566 5686 39618 5738
rect 15038 5630 15090 5682
rect 16774 5630 16826 5682
rect 20302 5630 20354 5682
rect 24166 5630 24218 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 6190 5294 6242 5346
rect 6862 5294 6914 5346
rect 9718 5294 9770 5346
rect 10334 5294 10386 5346
rect 3054 5182 3106 5234
rect 4958 5182 5010 5234
rect 7982 5182 8034 5234
rect 8318 5182 8370 5234
rect 14814 5182 14866 5234
rect 16718 5182 16770 5234
rect 18510 5182 18562 5234
rect 20750 5182 20802 5234
rect 2270 5070 2322 5122
rect 5854 5070 5906 5122
rect 6526 5070 6578 5122
rect 7534 5070 7586 5122
rect 7870 5055 7922 5107
rect 8430 5055 8482 5107
rect 8654 5070 8706 5122
rect 9214 5070 9266 5122
rect 9438 5070 9490 5122
rect 9998 5070 10050 5122
rect 14030 5070 14082 5122
rect 17502 5042 17554 5094
rect 20302 5070 20354 5122
rect 20638 5055 20690 5107
rect 21198 5070 21250 5122
rect 22430 5070 22482 5122
rect 22934 5126 22986 5178
rect 29318 5182 29370 5234
rect 33182 5182 33234 5234
rect 36318 5182 36370 5234
rect 37158 5182 37210 5234
rect 39342 5182 39394 5234
rect 44942 5182 44994 5234
rect 23102 5070 23154 5122
rect 23662 5070 23714 5122
rect 25566 5070 25618 5122
rect 26350 5070 26402 5122
rect 27022 5070 27074 5122
rect 27918 5070 27970 5122
rect 28198 5070 28250 5122
rect 28478 5070 28530 5122
rect 28702 5070 28754 5122
rect 29486 5070 29538 5122
rect 30494 5070 30546 5122
rect 31278 5070 31330 5122
rect 33630 5070 33682 5122
rect 34414 5070 34466 5122
rect 37438 5070 37490 5122
rect 38110 5070 38162 5122
rect 37886 5014 37938 5066
rect 38558 5070 38610 5122
rect 41246 5070 41298 5122
rect 41694 5042 41746 5094
rect 46846 5070 46898 5122
rect 47630 5070 47682 5122
rect 47854 5035 47906 5087
rect 47966 5042 48018 5094
rect 48190 5042 48242 5094
rect 48414 5042 48466 5094
rect 22188 4958 22240 5010
rect 48694 4958 48746 5010
rect 21534 4846 21586 4898
rect 26686 4846 26738 4898
rect 38222 4902 38274 4954
rect 27582 4846 27634 4898
rect 43038 4846 43090 4898
rect 49142 4846 49194 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 15374 4510 15426 4562
rect 24558 4510 24610 4562
rect 16046 4454 16098 4506
rect 18510 4454 18562 4506
rect 8878 4398 8930 4450
rect 22318 4398 22370 4450
rect 6190 4286 6242 4338
rect 6974 4286 7026 4338
rect 14366 4286 14418 4338
rect 15038 4286 15090 4338
rect 16214 4342 16266 4394
rect 15710 4286 15762 4338
rect 16046 4286 16098 4338
rect 16606 4286 16658 4338
rect 17726 4286 17778 4338
rect 17950 4286 18002 4338
rect 18734 4342 18786 4394
rect 22860 4398 22912 4450
rect 23774 4398 23826 4450
rect 23606 4342 23658 4394
rect 25230 4398 25282 4450
rect 26144 4398 26196 4450
rect 26630 4454 26682 4506
rect 31166 4510 31218 4562
rect 18398 4286 18450 4338
rect 18958 4286 19010 4338
rect 19630 4286 19682 4338
rect 20414 4286 20466 4338
rect 23102 4286 23154 4338
rect 25398 4342 25450 4394
rect 29598 4398 29650 4450
rect 38670 4398 38722 4450
rect 40966 4454 41018 4506
rect 47742 4510 47794 4562
rect 48974 4510 49026 4562
rect 44046 4398 44098 4450
rect 44606 4398 44658 4450
rect 24222 4286 24274 4338
rect 25902 4286 25954 4338
rect 26910 4286 26962 4338
rect 27694 4286 27746 4338
rect 32510 4313 32562 4365
rect 33182 4286 33234 4338
rect 35086 4286 35138 4338
rect 35870 4286 35922 4338
rect 35982 4286 36034 4338
rect 36766 4286 36818 4338
rect 39230 4330 39282 4382
rect 39454 4286 39506 4338
rect 39790 4286 39842 4338
rect 40126 4286 40178 4338
rect 41358 4286 41410 4338
rect 42142 4286 42194 4338
rect 47294 4286 47346 4338
rect 47406 4286 47458 4338
rect 48638 4286 48690 4338
rect 17446 4174 17498 4226
rect 39118 4174 39170 4226
rect 46510 4174 46562 4226
rect 14030 4062 14082 4114
rect 14702 4062 14754 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 31054 3726 31106 3778
rect 38838 3726 38890 3778
rect 42702 3726 42754 3778
rect 34974 3670 35026 3722
rect 48302 3726 48354 3778
rect 48974 3726 49026 3778
rect 17726 3614 17778 3666
rect 19630 3614 19682 3666
rect 22094 3614 22146 3666
rect 24782 3614 24834 3666
rect 26686 3614 26738 3666
rect 30606 3614 30658 3666
rect 36990 3614 37042 3666
rect 47630 3614 47682 3666
rect 14030 3474 14082 3526
rect 16942 3502 16994 3554
rect 21422 3474 21474 3526
rect 27470 3502 27522 3554
rect 29150 3502 29202 3554
rect 29486 3475 29538 3527
rect 29710 3502 29762 3554
rect 30158 3502 30210 3554
rect 30494 3487 30546 3539
rect 31390 3502 31442 3554
rect 32398 3502 32450 3554
rect 34638 3474 34690 3526
rect 35086 3502 35138 3554
rect 35422 3502 35474 3554
rect 36206 3474 36258 3526
rect 39118 3502 39170 3554
rect 39342 3502 39394 3554
rect 42030 3474 42082 3526
rect 43038 3502 43090 3554
rect 43766 3502 43818 3554
rect 44046 3474 44098 3526
rect 44270 3446 44322 3498
rect 44494 3474 44546 3526
rect 44606 3467 44658 3519
rect 45558 3467 45610 3519
rect 45838 3474 45890 3526
rect 46062 3446 46114 3498
rect 46230 3486 46282 3538
rect 46958 3502 47010 3554
rect 47294 3502 47346 3554
rect 47966 3502 48018 3554
rect 48638 3502 48690 3554
rect 1766 3278 1818 3330
rect 3222 3278 3274 3330
rect 5574 3334 5626 3386
rect 6806 3278 6858 3330
rect 8598 3278 8650 3330
rect 10390 3278 10442 3330
rect 12182 3278 12234 3330
rect 13526 3278 13578 3330
rect 15598 3278 15650 3330
rect 20134 3334 20186 3386
rect 40574 3390 40626 3442
rect 45334 3390 45386 3442
rect 23942 3278 23994 3330
rect 27750 3334 27802 3386
rect 29038 3334 29090 3386
rect 28422 3278 28474 3330
rect 46622 3278 46674 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 23942 2718 23994 2770
rect 24446 2718 24498 2770
<< metal2 >>
rect 6272 50200 6384 51000
rect 19040 50200 19152 51000
rect 31808 50200 31920 51000
rect 44576 50200 44688 51000
rect 5740 48356 5796 48366
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 5516 41748 5572 41758
rect 5516 41746 5684 41748
rect 5516 41694 5518 41746
rect 5570 41694 5684 41746
rect 5516 41692 5684 41694
rect 5516 41682 5572 41692
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 5628 41300 5684 41692
rect 5628 41234 5684 41244
rect 5516 41186 5572 41198
rect 5516 41134 5518 41186
rect 5570 41134 5572 41186
rect 5404 40516 5460 40526
rect 5516 40516 5572 41134
rect 5460 40460 5572 40516
rect 5404 40402 5460 40460
rect 5404 40350 5406 40402
rect 5458 40350 5460 40402
rect 5404 40338 5460 40350
rect 5740 40068 5796 48300
rect 6300 48356 6356 50200
rect 6300 48290 6356 48300
rect 14700 47740 14980 47796
rect 14364 47684 14420 47694
rect 14700 47684 14756 47740
rect 14364 47682 14756 47684
rect 14364 47630 14366 47682
rect 14418 47630 14756 47682
rect 14364 47628 14756 47630
rect 14364 47618 14420 47628
rect 14812 47570 14868 47582
rect 14812 47518 14814 47570
rect 14866 47518 14868 47570
rect 11788 47458 11844 47470
rect 11788 47406 11790 47458
rect 11842 47406 11844 47458
rect 11452 47236 11508 47246
rect 11004 47234 11508 47236
rect 11004 47182 11454 47234
rect 11506 47182 11508 47234
rect 11004 47180 11508 47182
rect 10220 46674 10276 46686
rect 10220 46622 10222 46674
rect 10274 46622 10276 46674
rect 9548 45892 9604 45902
rect 10220 45892 10276 46622
rect 11004 46674 11060 47180
rect 11452 47170 11508 47180
rect 11788 46900 11844 47406
rect 13244 47458 13300 47470
rect 13244 47406 13246 47458
rect 13298 47406 13300 47458
rect 13244 46900 13300 47406
rect 14120 47402 14176 47414
rect 14120 47350 14122 47402
rect 14174 47350 14176 47402
rect 14120 46900 14176 47350
rect 11788 46844 12180 46900
rect 13244 46844 13636 46900
rect 11004 46622 11006 46674
rect 11058 46622 11060 46674
rect 11004 46610 11060 46622
rect 9548 45890 10276 45892
rect 9548 45838 9550 45890
rect 9602 45838 10276 45890
rect 9548 45836 10276 45838
rect 11116 46004 11172 46014
rect 11116 45890 11172 45948
rect 11116 45838 11118 45890
rect 11170 45838 11172 45890
rect 11452 46002 11508 46014
rect 11452 45950 11454 46002
rect 11506 45950 11508 46002
rect 11452 45892 11508 45950
rect 9436 45108 9492 45118
rect 9548 45108 9604 45836
rect 11116 45826 11172 45838
rect 11340 45846 11396 45858
rect 11340 45794 11342 45846
rect 11394 45794 11396 45846
rect 11452 45826 11508 45836
rect 12012 45892 12068 45902
rect 12012 45798 12068 45836
rect 11340 45780 11396 45794
rect 11340 45714 11396 45724
rect 11676 45780 11732 45790
rect 9436 45106 9604 45108
rect 9436 45054 9438 45106
rect 9490 45054 9604 45106
rect 9436 45052 9604 45054
rect 9436 45042 9492 45052
rect 9100 44548 9156 44558
rect 9100 44454 9156 44492
rect 7420 44434 7476 44446
rect 7420 44382 7422 44434
rect 7474 44382 7476 44434
rect 7420 43988 7476 44382
rect 7868 44322 7924 44334
rect 7196 43932 7476 43988
rect 7532 44278 7588 44290
rect 7532 44226 7534 44278
rect 7586 44226 7588 44278
rect 6188 43538 6244 43550
rect 6188 43486 6190 43538
rect 6242 43486 6244 43538
rect 5852 41970 5908 41982
rect 6188 41972 6244 43486
rect 6972 43540 7028 43550
rect 7196 43540 7252 43932
rect 7532 43764 7588 44226
rect 7868 44270 7870 44322
rect 7922 44270 7924 44322
rect 7868 44100 7924 44270
rect 7868 44034 7924 44044
rect 8764 44324 8820 44334
rect 7532 43698 7588 43708
rect 6972 43538 7252 43540
rect 6972 43486 6974 43538
rect 7026 43486 7252 43538
rect 6972 43484 7252 43486
rect 6972 43474 7028 43484
rect 7196 43316 7252 43326
rect 7196 42978 7252 43260
rect 7196 42926 7198 42978
rect 7250 42926 7252 42978
rect 7196 42914 7252 42926
rect 7439 43092 7495 43102
rect 7439 42756 7495 43036
rect 7196 42754 7495 42756
rect 7196 42702 7441 42754
rect 7493 42702 7495 42754
rect 7196 42700 7495 42702
rect 5852 41918 5854 41970
rect 5906 41918 5908 41970
rect 5852 40292 5908 41918
rect 5964 41916 6244 41972
rect 6412 41972 6468 41982
rect 5964 40516 6020 41916
rect 6412 41878 6468 41916
rect 6636 41970 6692 41982
rect 6636 41918 6638 41970
rect 6690 41918 6692 41970
rect 6636 41860 6692 41918
rect 6916 41972 6972 41982
rect 6916 41878 6972 41916
rect 7196 41970 7252 42700
rect 7439 42690 7495 42700
rect 8316 42754 8372 42766
rect 8316 42702 8318 42754
rect 8370 42702 8372 42754
rect 7756 41985 7812 41997
rect 7196 41918 7198 41970
rect 7250 41918 7252 41970
rect 7196 41906 7252 41918
rect 7420 41970 7476 41982
rect 7420 41918 7422 41970
rect 7474 41918 7476 41970
rect 6636 41794 6692 41804
rect 6132 41746 6188 41758
rect 6132 41694 6134 41746
rect 6186 41694 6188 41746
rect 6132 41636 6188 41694
rect 7420 41748 7476 41918
rect 7756 41972 7758 41985
rect 7810 41972 7812 41985
rect 7756 41893 7812 41916
rect 8092 41972 8148 41982
rect 8316 41972 8372 42702
rect 8764 42754 8820 44268
rect 9436 44322 9492 44334
rect 9436 44270 9438 44322
rect 9490 44270 9492 44322
rect 9436 44212 9492 44270
rect 9548 44324 9604 45052
rect 10220 44994 10276 45006
rect 10220 44942 10222 44994
rect 10274 44942 10276 44994
rect 10220 44548 10276 44942
rect 10220 44482 10276 44492
rect 9548 44258 9604 44268
rect 9884 44324 9940 44334
rect 9884 44230 9940 44268
rect 9436 44146 9492 44156
rect 11340 44212 11396 44222
rect 11116 44100 11172 44110
rect 10780 43582 10836 43594
rect 9996 43538 10052 43550
rect 9996 43486 9998 43538
rect 10050 43486 10052 43538
rect 8876 43426 8932 43438
rect 8876 43374 8878 43426
rect 8930 43374 8932 43426
rect 8876 43316 8932 43374
rect 8876 43250 8932 43260
rect 9660 43314 9716 43326
rect 9660 43262 9662 43314
rect 9714 43262 9716 43314
rect 8764 42702 8766 42754
rect 8818 42702 8820 42754
rect 8764 42690 8820 42702
rect 9548 42754 9604 42766
rect 9548 42702 9550 42754
rect 9602 42702 9604 42754
rect 9548 42196 9604 42702
rect 9548 42130 9604 42140
rect 8092 41970 8260 41972
rect 8092 41918 8094 41970
rect 8146 41918 8260 41970
rect 8092 41916 8260 41918
rect 8092 41906 8148 41916
rect 7420 41682 7476 41692
rect 7644 41858 7700 41870
rect 7644 41806 7646 41858
rect 7698 41806 7700 41858
rect 6132 41580 6468 41636
rect 6300 41300 6356 41310
rect 6300 41206 6356 41244
rect 5964 40450 6020 40460
rect 6188 40516 6244 40526
rect 5852 40226 5908 40236
rect 4476 40012 4740 40022
rect 5740 40012 6132 40068
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 5628 39732 5684 39742
rect 5404 39730 5684 39732
rect 5404 39678 5630 39730
rect 5682 39678 5684 39730
rect 5404 39676 5684 39678
rect 5404 38834 5460 39676
rect 5628 39666 5684 39676
rect 5964 39620 6020 39630
rect 5740 39574 5796 39586
rect 5740 39522 5742 39574
rect 5794 39522 5796 39574
rect 5740 38948 5796 39522
rect 5740 38882 5796 38892
rect 5404 38782 5406 38834
rect 5458 38782 5460 38834
rect 5404 38770 5460 38782
rect 5516 38836 5572 38846
rect 3500 38724 3556 38762
rect 3500 38658 3556 38668
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 5516 38050 5572 38780
rect 5516 37998 5518 38050
rect 5570 37998 5572 38050
rect 5516 37986 5572 37998
rect 5964 37266 6020 39564
rect 5964 37214 5966 37266
rect 6018 37214 6020 37266
rect 5964 37202 6020 37214
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 6076 36372 6132 40012
rect 6188 38836 6244 40460
rect 6412 39732 6468 41580
rect 6748 40628 6804 40638
rect 6636 40429 6692 40441
rect 6636 40404 6638 40429
rect 6690 40404 6692 40429
rect 6636 40337 6692 40348
rect 6412 39666 6468 39676
rect 6524 40292 6580 40302
rect 6188 38742 6244 38780
rect 6300 39508 6356 39518
rect 6300 38276 6356 39452
rect 6524 39450 6580 40236
rect 6748 40180 6804 40572
rect 7644 40628 7700 41806
rect 8204 41860 8260 41916
rect 8204 41076 8260 41804
rect 8316 41748 8372 41916
rect 8876 41970 8932 41982
rect 8876 41918 8878 41970
rect 8930 41918 8932 41970
rect 8316 41682 8372 41692
rect 8596 41748 8652 41758
rect 8596 41654 8652 41692
rect 8540 41188 8596 41198
rect 8204 40982 8260 41020
rect 8428 41186 8596 41188
rect 8428 41134 8542 41186
rect 8594 41134 8596 41186
rect 8428 41132 8596 41134
rect 7644 40562 7700 40572
rect 8316 40516 8372 40526
rect 6636 40124 6804 40180
rect 8204 40404 8260 40414
rect 6636 39618 6692 40124
rect 7308 39844 7364 39854
rect 6636 39566 6638 39618
rect 6690 39566 6692 39618
rect 6636 39554 6692 39566
rect 6860 39732 6916 39742
rect 6860 39579 6916 39676
rect 6860 39527 6862 39579
rect 6914 39527 6916 39579
rect 7308 39618 7364 39788
rect 7308 39566 7310 39618
rect 7362 39566 7364 39618
rect 7756 39732 7812 39742
rect 7756 39580 7812 39676
rect 7308 39554 7364 39566
rect 7644 39562 7700 39574
rect 6860 39508 6916 39527
rect 6524 39398 6526 39450
rect 6578 39398 6580 39450
rect 6524 39386 6580 39398
rect 6767 39452 6916 39508
rect 7644 39510 7646 39562
rect 7698 39510 7700 39562
rect 7756 39528 7758 39580
rect 7810 39528 7812 39580
rect 7756 39516 7812 39528
rect 6524 38948 6580 38958
rect 6524 38854 6580 38892
rect 6767 38890 6823 39452
rect 6767 38838 6769 38890
rect 6821 38838 6823 38890
rect 6767 38826 6823 38838
rect 7644 38836 7700 39510
rect 7644 38770 7700 38780
rect 8204 38744 8260 40348
rect 8316 40402 8372 40460
rect 8316 40350 8318 40402
rect 8370 40350 8372 40402
rect 8316 40338 8372 40350
rect 8428 39640 8484 41132
rect 8540 41122 8596 41132
rect 8764 41186 8820 41198
rect 8764 41134 8766 41186
rect 8818 41134 8820 41186
rect 8652 41076 8708 41086
rect 8428 39618 8540 39640
rect 8428 39566 8486 39618
rect 8538 39566 8540 39618
rect 8428 39554 8540 39566
rect 8652 39618 8708 41020
rect 8764 39956 8820 41134
rect 8876 40628 8932 41918
rect 9100 41972 9156 41982
rect 9660 41972 9716 43262
rect 9996 43316 10052 43486
rect 10556 43540 10612 43550
rect 10556 43538 10724 43540
rect 10556 43486 10558 43538
rect 10610 43486 10724 43538
rect 10556 43484 10724 43486
rect 10556 43474 10612 43484
rect 9996 43250 10052 43260
rect 9996 42196 10052 42206
rect 9996 42102 10052 42140
rect 10332 42196 10388 42206
rect 9100 41970 9604 41972
rect 9100 41918 9102 41970
rect 9154 41918 9604 41970
rect 9100 41916 9604 41918
rect 9100 41906 9156 41916
rect 9044 41076 9100 41086
rect 9044 40982 9100 41020
rect 8876 40562 8932 40572
rect 9548 40404 9604 41916
rect 9660 41188 9716 41916
rect 10332 41970 10388 42140
rect 10332 41918 10334 41970
rect 10386 41918 10388 41970
rect 10332 41906 10388 41918
rect 10668 41870 10724 43484
rect 10780 43530 10782 43582
rect 10834 43530 10836 43582
rect 10780 42532 10836 43530
rect 10892 43540 10948 43550
rect 10892 43426 10948 43484
rect 10892 43374 10894 43426
rect 10946 43374 10948 43426
rect 10892 43362 10948 43374
rect 10780 42466 10836 42476
rect 10892 41972 10948 41982
rect 11116 41972 11172 44044
rect 11340 43706 11396 44156
rect 11340 43654 11342 43706
rect 11394 43654 11396 43706
rect 11340 43642 11396 43654
rect 11452 43764 11508 43774
rect 11340 43540 11396 43550
rect 11452 43540 11508 43708
rect 11228 43538 11508 43540
rect 11228 43486 11342 43538
rect 11394 43486 11508 43538
rect 11228 43484 11508 43486
rect 11676 43594 11732 45724
rect 12124 45722 12180 46844
rect 13356 46674 13412 46686
rect 13356 46622 13358 46674
rect 13410 46622 13412 46674
rect 12908 46564 12964 46574
rect 13356 46564 13412 46622
rect 12908 46562 13412 46564
rect 12908 46510 12910 46562
rect 12962 46510 13412 46562
rect 12908 46508 13412 46510
rect 12908 46498 12964 46508
rect 12348 46452 12404 46462
rect 12348 45863 12404 46396
rect 13356 46004 13412 46508
rect 13356 45938 13412 45948
rect 13468 46674 13524 46686
rect 13468 46622 13470 46674
rect 13522 46622 13524 46674
rect 12572 45892 12628 45902
rect 12348 45811 12350 45863
rect 12402 45811 12404 45863
rect 12348 45799 12404 45811
rect 12460 45890 12628 45892
rect 12460 45838 12574 45890
rect 12626 45838 12628 45890
rect 12460 45836 12628 45838
rect 12124 45670 12126 45722
rect 12178 45670 12180 45722
rect 12124 45658 12180 45670
rect 12460 45444 12516 45836
rect 12572 45826 12628 45836
rect 12012 45388 12516 45444
rect 13468 45780 13524 46622
rect 13580 46564 13636 46844
rect 13580 46228 13636 46508
rect 13916 46844 14176 46900
rect 13748 46452 13804 46462
rect 13916 46452 13972 46844
rect 13804 46396 13972 46452
rect 14028 46674 14084 46686
rect 14028 46622 14030 46674
rect 14082 46622 14084 46674
rect 14028 46452 14084 46622
rect 14812 46674 14868 47518
rect 14924 47443 14980 47740
rect 19068 47582 19124 50200
rect 30660 48018 30716 48030
rect 30660 47966 30662 48018
rect 30714 47966 30716 48018
rect 20972 47740 21252 47796
rect 20972 47684 21028 47740
rect 19012 47570 19124 47582
rect 19012 47518 19014 47570
rect 19066 47518 19124 47570
rect 19012 47506 19124 47518
rect 14924 47391 14926 47443
rect 14978 47391 14980 47443
rect 14924 47379 14980 47391
rect 15148 47458 15204 47470
rect 15148 47406 15150 47458
rect 15202 47406 15204 47458
rect 15148 46900 15204 47406
rect 19068 47460 19124 47506
rect 20636 47628 21028 47684
rect 19180 47460 19236 47470
rect 19068 47458 19236 47460
rect 19068 47406 19182 47458
rect 19234 47406 19236 47458
rect 19068 47404 19236 47406
rect 19180 47394 19236 47404
rect 19516 47236 19572 47246
rect 14812 46622 14814 46674
rect 14866 46622 14868 46674
rect 14812 46610 14868 46622
rect 15036 46844 15204 46900
rect 18508 47234 19572 47236
rect 18508 47182 19518 47234
rect 19570 47182 19572 47234
rect 18508 47180 19572 47182
rect 14028 46396 14980 46452
rect 13748 46358 13804 46396
rect 13580 46172 14084 46228
rect 13692 46004 13748 46014
rect 12012 43764 12068 45388
rect 12124 45220 12180 45230
rect 12124 45218 12964 45220
rect 12124 45166 12126 45218
rect 12178 45166 12964 45218
rect 12124 45164 12964 45166
rect 12124 45154 12180 45164
rect 12740 44996 12796 45006
rect 12684 44994 12796 44996
rect 12684 44942 12742 44994
rect 12794 44942 12796 44994
rect 12684 44930 12796 44942
rect 12460 44434 12516 44446
rect 12460 44382 12462 44434
rect 12514 44382 12516 44434
rect 12124 44294 12180 44306
rect 12124 44242 12126 44294
rect 12178 44242 12180 44294
rect 12124 44212 12180 44242
rect 12124 44146 12180 44156
rect 12012 43698 12068 43708
rect 11676 43542 11678 43594
rect 11730 43542 11732 43594
rect 11228 42420 11284 43484
rect 11340 43474 11396 43484
rect 11564 43428 11620 43438
rect 11452 42644 11508 42654
rect 11228 42354 11284 42364
rect 11340 42642 11508 42644
rect 11340 42590 11454 42642
rect 11506 42590 11508 42642
rect 11340 42588 11508 42590
rect 11228 42196 11284 42206
rect 11228 42138 11284 42140
rect 11228 42086 11230 42138
rect 11282 42086 11284 42138
rect 11228 42074 11284 42086
rect 11228 41972 11284 41982
rect 10892 41970 11060 41972
rect 10892 41918 10894 41970
rect 10946 41918 11060 41970
rect 10892 41916 11060 41918
rect 11116 41970 11284 41972
rect 11116 41918 11230 41970
rect 11282 41918 11284 41970
rect 11116 41916 11284 41918
rect 10892 41906 10948 41916
rect 10668 41860 10780 41870
rect 10668 41804 10724 41860
rect 10724 41802 10780 41804
rect 10332 41748 10388 41758
rect 10724 41750 10726 41802
rect 10778 41750 10780 41802
rect 10724 41738 10780 41750
rect 10108 41412 10164 41422
rect 9884 41188 9940 41198
rect 9660 41132 9884 41188
rect 9884 41094 9940 41132
rect 10108 41186 10164 41356
rect 10108 41134 10110 41186
rect 10162 41134 10164 41186
rect 10108 41122 10164 41134
rect 10220 41354 10276 41366
rect 10220 41302 10222 41354
rect 10274 41302 10276 41354
rect 10220 40740 10276 41302
rect 10220 40674 10276 40684
rect 9212 40402 9604 40404
rect 9212 40350 9550 40402
rect 9602 40350 9604 40402
rect 9212 40348 9604 40350
rect 8764 39900 9044 39956
rect 8820 39786 8876 39798
rect 8820 39734 8822 39786
rect 8874 39734 8876 39786
rect 8820 39732 8876 39734
rect 8820 39666 8876 39676
rect 8652 39566 8654 39618
rect 8706 39566 8708 39618
rect 8652 39554 8708 39566
rect 8316 39508 8372 39518
rect 8316 39414 8372 39452
rect 8204 38722 8316 38744
rect 8204 38670 8262 38722
rect 8314 38670 8316 38722
rect 8204 38668 8316 38670
rect 8204 38612 8372 38668
rect 6188 38220 6356 38276
rect 6188 37380 6244 38220
rect 8204 38164 8260 38174
rect 8204 38070 8260 38108
rect 6300 38052 6356 38062
rect 6300 38050 6468 38052
rect 6300 37998 6302 38050
rect 6354 37998 6468 38050
rect 6300 37996 6468 37998
rect 6300 37986 6356 37996
rect 6188 37324 6300 37380
rect 6244 37322 6300 37324
rect 6244 37270 6246 37322
rect 6298 37270 6300 37322
rect 6244 37258 6300 37270
rect 6412 37154 6468 37996
rect 6412 37102 6414 37154
rect 6466 37102 6468 37154
rect 6412 37090 6468 37102
rect 7868 36932 7924 36942
rect 6636 36484 6692 36494
rect 6636 36390 6692 36428
rect 7308 36482 7364 36494
rect 7308 36430 7310 36482
rect 7362 36430 7364 36482
rect 5852 36316 6132 36372
rect 5180 35698 5236 35710
rect 5180 35646 5182 35698
rect 5234 35646 5236 35698
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4844 34916 4900 34926
rect 4844 34822 4900 34860
rect 5180 34916 5236 35646
rect 5180 34850 5236 34860
rect 5516 34916 5572 34926
rect 5852 34916 5908 36316
rect 6300 36260 6356 36270
rect 6188 36258 6356 36260
rect 6188 36206 6302 36258
rect 6354 36206 6356 36258
rect 6188 36204 6356 36206
rect 6188 35924 6244 36204
rect 6300 36194 6356 36204
rect 5964 35868 6244 35924
rect 5964 35698 6020 35868
rect 5964 35646 5966 35698
rect 6018 35646 6020 35698
rect 5964 35634 6020 35646
rect 7308 35028 7364 36430
rect 7868 35812 7924 36876
rect 8092 36482 8148 36494
rect 8092 36430 8094 36482
rect 8146 36430 8148 36482
rect 8092 35924 8148 36430
rect 8092 35858 8148 35868
rect 7868 35718 7924 35756
rect 7420 35028 7476 35038
rect 7308 35026 7476 35028
rect 7308 34974 7422 35026
rect 7474 34974 7476 35026
rect 7308 34972 7476 34974
rect 5852 34860 6020 34916
rect 5516 34130 5572 34860
rect 5516 34078 5518 34130
rect 5570 34078 5572 34130
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 5516 33684 5572 34078
rect 5852 34690 5908 34702
rect 5852 34638 5854 34690
rect 5906 34638 5908 34690
rect 5852 34132 5908 34638
rect 5852 34066 5908 34076
rect 5068 32564 5124 32574
rect 5516 32564 5572 33628
rect 5068 32562 5572 32564
rect 5068 32510 5070 32562
rect 5122 32510 5572 32562
rect 5068 32508 5572 32510
rect 5068 32498 5124 32508
rect 2380 32450 2436 32462
rect 2380 32398 2382 32450
rect 2434 32398 2436 32450
rect 2044 31780 2100 31790
rect 1596 30994 1652 31006
rect 1596 30942 1598 30994
rect 1650 30942 1652 30994
rect 1596 29540 1652 30942
rect 1596 29484 1988 29540
rect 1596 28644 1652 29484
rect 1932 29426 1988 29484
rect 1932 29374 1934 29426
rect 1986 29374 1988 29426
rect 1932 29362 1988 29374
rect 1596 27074 1652 28588
rect 1596 27022 1598 27074
rect 1650 27022 1652 27074
rect 1596 27010 1652 27022
rect 1932 27860 1988 27870
rect 2044 27860 2100 31724
rect 2380 31220 2436 32398
rect 4284 32450 4340 32462
rect 4284 32398 4286 32450
rect 4338 32398 4340 32450
rect 4284 31948 4340 32398
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4620 31948 4676 31958
rect 5964 31948 6020 34860
rect 6188 34914 6244 34926
rect 6188 34862 6190 34914
rect 6242 34862 6244 34914
rect 7420 34916 7476 34972
rect 6188 34468 6244 34862
rect 6636 34886 6692 34898
rect 6636 34834 6638 34886
rect 6690 34834 6692 34886
rect 6636 34692 6692 34834
rect 6636 34626 6692 34636
rect 6188 34402 6244 34412
rect 6300 34132 6356 34142
rect 6300 34038 6356 34076
rect 6972 33684 7028 33694
rect 6972 33346 7028 33628
rect 7420 33684 7476 34860
rect 8316 34692 8372 38612
rect 8428 38612 8484 39554
rect 8988 38948 9044 39900
rect 9212 39732 9268 40348
rect 9548 40338 9604 40348
rect 9660 40628 9716 40638
rect 9660 39732 9716 40572
rect 9884 40628 9940 40638
rect 9212 39583 9268 39676
rect 9436 39676 9716 39732
rect 9772 40404 9828 40414
rect 9436 39620 9492 39676
rect 9212 39531 9214 39583
rect 9266 39531 9268 39583
rect 9212 39519 9268 39531
rect 9380 39583 9492 39620
rect 9380 39531 9382 39583
rect 9434 39531 9492 39583
rect 9772 39590 9828 40348
rect 9884 40402 9940 40572
rect 10332 40628 10388 41692
rect 10612 41412 10668 41422
rect 10612 41318 10668 41356
rect 10332 40562 10388 40572
rect 10444 41186 10500 41198
rect 10444 41134 10446 41186
rect 10498 41134 10500 41186
rect 9884 40350 9886 40402
rect 9938 40350 9940 40402
rect 9884 40338 9940 40350
rect 10220 40516 10276 40526
rect 10108 40292 10164 40302
rect 10108 40198 10164 40236
rect 10220 40068 10276 40460
rect 10444 40402 10500 41134
rect 10892 41188 10948 41198
rect 11004 41188 11060 41916
rect 11116 41188 11172 41198
rect 11004 41132 11116 41188
rect 10892 41094 10948 41132
rect 11116 41122 11172 41132
rect 11060 40964 11116 40974
rect 10780 40962 11116 40964
rect 10780 40910 11062 40962
rect 11114 40910 11116 40962
rect 10780 40908 11116 40910
rect 10780 40516 10836 40908
rect 11060 40898 11116 40908
rect 10444 40350 10446 40402
rect 10498 40350 10500 40402
rect 10220 40012 10388 40068
rect 9380 39519 9492 39531
rect 9436 39060 9492 39519
rect 9548 39562 9604 39574
rect 9548 39510 9550 39562
rect 9602 39510 9604 39562
rect 9772 39538 9774 39590
rect 9826 39538 9828 39590
rect 9772 39526 9828 39538
rect 9548 39284 9604 39510
rect 9548 39218 9604 39228
rect 10052 39506 10108 39518
rect 10052 39454 10054 39506
rect 10106 39454 10108 39506
rect 8596 38836 8652 38846
rect 8596 38742 8652 38780
rect 8876 38834 8932 38846
rect 8876 38782 8878 38834
rect 8930 38782 8932 38834
rect 8428 38164 8484 38556
rect 8876 38276 8932 38782
rect 8876 38210 8932 38220
rect 8484 38108 8708 38164
rect 8428 38098 8484 38108
rect 8652 38050 8708 38108
rect 8988 38052 9044 38892
rect 9324 39004 9492 39060
rect 9100 38834 9156 38846
rect 9100 38782 9102 38834
rect 9154 38782 9156 38834
rect 9100 38668 9156 38782
rect 9100 38612 9268 38668
rect 9212 38162 9268 38612
rect 9324 38500 9380 39004
rect 9660 38948 9716 38958
rect 9492 38890 9548 38902
rect 9492 38838 9494 38890
rect 9546 38838 9548 38890
rect 9492 38612 9548 38838
rect 9660 38890 9716 38892
rect 9660 38838 9662 38890
rect 9714 38838 9716 38890
rect 10052 38948 10108 39454
rect 9660 38826 9716 38838
rect 9884 38873 9940 38885
rect 10052 38882 10108 38892
rect 9884 38821 9886 38873
rect 9938 38821 9940 38873
rect 9492 38546 9548 38556
rect 9772 38724 9828 38734
rect 9324 38434 9380 38444
rect 9212 38110 9214 38162
rect 9266 38110 9268 38162
rect 9212 38098 9268 38110
rect 9772 38164 9828 38668
rect 9884 38276 9940 38821
rect 10332 38612 10388 40012
rect 10444 39284 10500 40350
rect 10668 40460 10836 40516
rect 11116 40740 11172 40750
rect 10668 40404 10724 40460
rect 10668 40310 10724 40348
rect 11116 40402 11172 40684
rect 11116 40350 11118 40402
rect 11170 40350 11172 40402
rect 11116 40338 11172 40350
rect 10780 40292 10836 40302
rect 10780 39618 10836 40236
rect 10780 39566 10782 39618
rect 10834 39566 10836 39618
rect 10780 39554 10836 39566
rect 10892 39956 10948 39966
rect 10892 39618 10948 39900
rect 10892 39566 10894 39618
rect 10946 39566 10948 39618
rect 11228 39620 11284 41916
rect 11340 41188 11396 42588
rect 11452 42578 11508 42588
rect 11340 41122 11396 41132
rect 11452 42420 11508 42430
rect 11452 40964 11508 42364
rect 11564 42026 11620 43372
rect 11676 42644 11732 43542
rect 11900 43540 11956 43550
rect 12460 43540 12516 44382
rect 11900 43538 12516 43540
rect 11900 43486 11902 43538
rect 11954 43486 12516 43538
rect 11900 43484 12516 43486
rect 12572 44278 12628 44290
rect 12572 44226 12574 44278
rect 12626 44226 12628 44278
rect 12572 43540 12628 44226
rect 12684 44212 12740 44930
rect 12908 44324 12964 45164
rect 13468 45106 13524 45724
rect 13580 45778 13636 45790
rect 13580 45726 13582 45778
rect 13634 45726 13636 45778
rect 13580 45220 13636 45726
rect 13580 45154 13636 45164
rect 13468 45054 13470 45106
rect 13522 45054 13524 45106
rect 13468 45042 13524 45054
rect 13692 45145 13748 45948
rect 13823 45834 13879 45846
rect 13823 45782 13825 45834
rect 13877 45782 13879 45834
rect 13823 45332 13879 45782
rect 13692 45093 13694 45145
rect 13746 45093 13748 45145
rect 13356 44324 13412 44334
rect 12908 44322 13412 44324
rect 12908 44270 12910 44322
rect 12962 44270 13358 44322
rect 13410 44270 13412 44322
rect 12908 44268 13412 44270
rect 13692 44324 13748 45093
rect 13804 45276 13879 45332
rect 13804 44996 13860 45276
rect 14028 45106 14084 46172
rect 14700 45890 14756 45902
rect 14700 45838 14702 45890
rect 14754 45838 14756 45890
rect 14700 45444 14756 45838
rect 14028 45054 14030 45106
rect 14082 45054 14084 45106
rect 14028 45042 14084 45054
rect 14252 45164 14644 45220
rect 13916 44996 13972 45006
rect 13804 44994 13972 44996
rect 13804 44942 13918 44994
rect 13970 44942 13972 44994
rect 13804 44940 13972 44942
rect 13916 44884 13972 44940
rect 14252 44884 14308 45164
rect 14588 45150 14644 45164
rect 14588 45098 14590 45150
rect 14642 45098 14644 45150
rect 14588 45086 14644 45098
rect 14700 45108 14756 45388
rect 14924 45890 14980 46396
rect 15036 46340 15092 46844
rect 17612 46674 17668 46686
rect 17612 46622 17614 46674
rect 17666 46622 17668 46674
rect 16716 46564 16772 46574
rect 16716 46470 16772 46508
rect 17444 46452 17500 46462
rect 17444 46358 17500 46396
rect 15036 46284 15204 46340
rect 14924 45838 14926 45890
rect 14978 45838 14980 45890
rect 14812 45108 14868 45118
rect 14700 45106 14868 45108
rect 14700 45054 14814 45106
rect 14866 45054 14868 45106
rect 14700 45052 14868 45054
rect 14812 45042 14868 45052
rect 14476 44996 14532 45006
rect 13916 44828 14308 44884
rect 14364 44994 14532 44996
rect 14364 44942 14478 44994
rect 14530 44942 14532 44994
rect 14364 44940 14532 44942
rect 13804 44324 13860 44334
rect 13692 44322 13860 44324
rect 13692 44270 13806 44322
rect 13858 44270 13860 44322
rect 13692 44268 13860 44270
rect 12908 44258 12964 44268
rect 12684 44146 12740 44156
rect 13020 43652 13076 43662
rect 11900 43474 11956 43484
rect 12572 43474 12628 43484
rect 12796 43538 12852 43550
rect 12796 43486 12798 43538
rect 12850 43486 12852 43538
rect 12516 43316 12572 43326
rect 11676 42578 11732 42588
rect 11788 43314 12572 43316
rect 11788 43262 12518 43314
rect 12570 43262 12572 43314
rect 11788 43260 12572 43262
rect 11564 41974 11566 42026
rect 11618 41974 11620 42026
rect 11564 41962 11620 41974
rect 11788 41970 11844 43260
rect 12516 43250 12572 43260
rect 12572 42980 12628 42990
rect 12236 42756 12292 42766
rect 12236 42662 12292 42700
rect 12572 42698 12628 42924
rect 12124 42644 12180 42654
rect 12124 42586 12180 42588
rect 12124 42534 12126 42586
rect 12178 42534 12180 42586
rect 12124 42522 12180 42534
rect 12572 42646 12574 42698
rect 12626 42646 12628 42698
rect 12796 42756 12852 43486
rect 12908 43538 12964 43550
rect 12908 43486 12910 43538
rect 12962 43486 12964 43538
rect 12908 42980 12964 43486
rect 12908 42914 12964 42924
rect 12796 42690 12852 42700
rect 12908 42756 12964 42766
rect 13020 42756 13076 43596
rect 12908 42754 13020 42756
rect 12908 42702 12910 42754
rect 12962 42702 13020 42754
rect 12908 42700 13020 42702
rect 12908 42690 12964 42700
rect 13020 42662 13076 42700
rect 11788 41918 11790 41970
rect 11842 41918 11844 41970
rect 11788 41906 11844 41918
rect 12344 42008 12400 42020
rect 12344 41972 12346 42008
rect 12398 41972 12400 42008
rect 12344 41524 12400 41916
rect 12572 41860 12628 42646
rect 13020 41972 13076 41982
rect 13132 41972 13188 44268
rect 13356 44258 13412 44268
rect 13804 44258 13860 44268
rect 13524 44098 13580 44110
rect 13972 44100 14028 44110
rect 13524 44046 13526 44098
rect 13578 44046 13580 44098
rect 13524 43652 13580 44046
rect 13916 44098 14028 44100
rect 13916 44046 13974 44098
rect 14026 44046 14028 44098
rect 13916 44034 14028 44046
rect 13524 43586 13580 43596
rect 13692 43764 13748 43774
rect 13244 43540 13300 43550
rect 13244 42756 13300 43484
rect 13692 43538 13748 43708
rect 13692 43486 13694 43538
rect 13746 43486 13748 43538
rect 13692 43474 13748 43486
rect 13804 43538 13860 43550
rect 13804 43486 13806 43538
rect 13858 43486 13860 43538
rect 13804 43428 13860 43486
rect 13804 43362 13860 43372
rect 13412 43314 13468 43326
rect 13412 43262 13414 43314
rect 13466 43262 13468 43314
rect 13412 43092 13468 43262
rect 13916 43204 13972 44034
rect 14364 43764 14420 44940
rect 14476 44930 14532 44940
rect 14812 44436 14868 44446
rect 14028 43540 14084 43550
rect 14028 43446 14084 43484
rect 13916 43148 14196 43204
rect 13412 43026 13468 43036
rect 13244 42700 13412 42756
rect 13020 41970 13188 41972
rect 13020 41918 13022 41970
rect 13074 41918 13188 41970
rect 13020 41916 13188 41918
rect 13020 41906 13076 41916
rect 12572 41794 12628 41804
rect 12796 41802 12852 41814
rect 12796 41750 12798 41802
rect 12850 41750 12852 41802
rect 12344 41468 12404 41524
rect 11676 41188 11732 41198
rect 11676 41094 11732 41132
rect 11452 40908 11732 40964
rect 11452 40628 11508 40638
rect 11452 40516 11508 40572
rect 10892 39554 10948 39566
rect 11058 39562 11114 39574
rect 10444 39218 10500 39228
rect 11058 39510 11060 39562
rect 11112 39510 11114 39562
rect 11058 39172 11114 39510
rect 11228 39172 11284 39564
rect 11058 39116 11172 39172
rect 10444 39060 10500 39070
rect 10444 38946 10500 39004
rect 10444 38894 10446 38946
rect 10498 38894 10500 38946
rect 10444 38882 10500 38894
rect 11004 38836 11060 38846
rect 11004 38742 11060 38780
rect 10220 38556 10388 38612
rect 11116 38666 11172 39116
rect 11228 39106 11284 39116
rect 11340 40460 11508 40516
rect 11340 38834 11396 40460
rect 11452 40458 11508 40460
rect 11452 40406 11454 40458
rect 11506 40406 11508 40458
rect 11452 40394 11508 40406
rect 11452 40292 11508 40302
rect 11452 40198 11508 40236
rect 11676 39844 11732 40908
rect 12348 40852 12404 41468
rect 12796 41300 12852 41750
rect 12684 41244 12852 41300
rect 12552 41188 12608 41208
rect 12552 41130 12608 41132
rect 12552 41078 12554 41130
rect 12606 41078 12608 41130
rect 12552 40852 12608 41078
rect 11900 40796 12404 40852
rect 12460 40796 12608 40852
rect 11452 39732 11508 39742
rect 11452 39638 11508 39676
rect 11340 38782 11342 38834
rect 11394 38782 11396 38834
rect 11340 38770 11396 38782
rect 11116 38614 11118 38666
rect 11170 38614 11172 38666
rect 11116 38602 11172 38614
rect 9884 38210 9940 38220
rect 9996 38500 10052 38510
rect 8652 37998 8654 38050
rect 8706 37998 8708 38050
rect 8652 37986 8708 37998
rect 8764 38050 9044 38052
rect 8764 37998 8990 38050
rect 9042 37998 9044 38050
rect 8764 37996 9044 37998
rect 8764 37828 8820 37996
rect 8988 37986 9044 37996
rect 9548 38052 9604 38062
rect 8596 37772 8820 37828
rect 8596 37490 8652 37772
rect 8596 37438 8598 37490
rect 8650 37438 8652 37490
rect 8596 37426 8652 37438
rect 9212 37716 9268 37726
rect 8428 37266 8484 37278
rect 8428 37214 8430 37266
rect 8482 37214 8484 37266
rect 8428 36932 8484 37214
rect 8428 36866 8484 36876
rect 9212 36260 9268 37660
rect 9548 37502 9604 37996
rect 9772 38050 9828 38108
rect 9772 37998 9774 38050
rect 9826 37998 9828 38050
rect 9772 37986 9828 37998
rect 9548 37490 9660 37502
rect 9548 37438 9606 37490
rect 9658 37438 9660 37490
rect 9548 37436 9660 37438
rect 9604 37426 9660 37436
rect 8988 36204 9268 36260
rect 9772 37266 9828 37278
rect 9772 37214 9774 37266
rect 9826 37214 9828 37266
rect 8764 35924 8820 35934
rect 8764 35830 8820 35868
rect 8316 34626 8372 34636
rect 8204 34132 8260 34142
rect 8204 34038 8260 34076
rect 7420 33618 7476 33628
rect 7756 33908 7812 33918
rect 7756 33458 7812 33852
rect 8764 33908 8820 33918
rect 8764 33814 8820 33852
rect 7756 33406 7758 33458
rect 7810 33406 7812 33458
rect 7756 33394 7812 33406
rect 6972 33294 6974 33346
rect 7026 33294 7028 33346
rect 6972 33282 7028 33294
rect 8988 33348 9044 36204
rect 9100 35700 9156 35710
rect 9604 35700 9660 35710
rect 9100 35698 9660 35700
rect 9100 35646 9102 35698
rect 9154 35646 9606 35698
rect 9658 35646 9660 35698
rect 9100 35644 9660 35646
rect 9100 35634 9156 35644
rect 9604 35634 9660 35644
rect 9212 34692 9268 34702
rect 9100 34130 9156 34142
rect 9100 34078 9102 34130
rect 9154 34078 9156 34130
rect 9100 33572 9156 34078
rect 9100 33506 9156 33516
rect 8988 33282 9044 33292
rect 8764 32788 8820 32798
rect 8764 32694 8820 32732
rect 7420 32577 7476 32589
rect 7084 32562 7140 32574
rect 7084 32510 7086 32562
rect 7138 32510 7140 32562
rect 3612 31892 4340 31948
rect 4396 31946 4676 31948
rect 4396 31894 4622 31946
rect 4674 31894 4676 31946
rect 4396 31892 4676 31894
rect 5404 31892 5796 31948
rect 5964 31892 6244 31948
rect 3612 31890 3668 31892
rect 3612 31838 3614 31890
rect 3666 31838 3668 31890
rect 3612 31826 3668 31838
rect 3164 31780 3220 31790
rect 3164 31686 3220 31724
rect 3500 31734 3556 31746
rect 3500 31682 3502 31734
rect 3554 31682 3556 31734
rect 3500 31668 3556 31682
rect 4396 31668 4452 31892
rect 4620 31882 4676 31892
rect 5292 31836 5460 31892
rect 3500 31612 4452 31668
rect 4732 31778 4788 31790
rect 4956 31780 5012 31790
rect 4732 31726 4734 31778
rect 4786 31726 4788 31778
rect 2380 31154 2436 31164
rect 4172 31220 4228 31230
rect 4060 30996 4116 31006
rect 2380 30882 2436 30894
rect 2380 30830 2382 30882
rect 2434 30830 2436 30882
rect 2380 30436 2436 30830
rect 2492 30436 2548 30446
rect 2380 30434 2548 30436
rect 2380 30382 2494 30434
rect 2546 30382 2548 30434
rect 2380 30380 2548 30382
rect 2492 30370 2548 30380
rect 2940 30324 2996 30334
rect 2828 30212 2884 30222
rect 2828 30118 2884 30156
rect 2716 29314 2772 29326
rect 2716 29262 2718 29314
rect 2770 29262 2772 29314
rect 2716 28532 2772 29262
rect 2940 29092 2996 30268
rect 4060 30210 4116 30940
rect 4060 30158 4062 30210
rect 4114 30158 4116 30210
rect 4060 30146 4116 30158
rect 4172 30212 4228 31164
rect 4732 31108 4788 31726
rect 4732 31042 4788 31052
rect 4844 31778 5012 31780
rect 4844 31726 4958 31778
rect 5010 31726 5012 31778
rect 4844 31724 5012 31726
rect 4284 30884 4340 30894
rect 4284 30790 4340 30828
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4844 30324 4900 31724
rect 4956 31714 5012 31724
rect 4956 31220 5012 31230
rect 4956 30994 5012 31164
rect 4956 30942 4958 30994
rect 5010 30942 5012 30994
rect 5292 30994 5348 31836
rect 5516 31778 5572 31790
rect 5516 31726 5518 31778
rect 5570 31726 5572 31778
rect 4956 30930 5012 30942
rect 5124 30938 5180 30950
rect 5124 30886 5126 30938
rect 5178 30886 5180 30938
rect 5124 30884 5180 30886
rect 5124 30772 5180 30828
rect 5068 30716 5180 30772
rect 5292 30942 5294 30994
rect 5346 30942 5348 30994
rect 4956 30324 5012 30334
rect 4844 30268 4956 30324
rect 4956 30230 5012 30268
rect 4396 30212 4452 30222
rect 4172 30210 4452 30212
rect 4172 30158 4398 30210
rect 4450 30158 4452 30210
rect 5068 30210 5124 30716
rect 4172 30156 4452 30158
rect 4396 30146 4452 30156
rect 4732 30154 4788 30166
rect 3948 30100 4004 30110
rect 3836 29652 3892 29662
rect 2940 29036 3108 29092
rect 2940 28868 2996 28878
rect 2940 28642 2996 28812
rect 2940 28590 2942 28642
rect 2994 28590 2996 28642
rect 2940 28578 2996 28590
rect 3052 28644 3108 29036
rect 3612 28754 3668 28766
rect 3612 28702 3614 28754
rect 3666 28702 3668 28754
rect 3052 28612 3164 28644
rect 3052 28588 3110 28612
rect 3108 28560 3110 28588
rect 3162 28560 3164 28612
rect 3108 28548 3164 28560
rect 3612 28532 3668 28702
rect 3836 28644 3892 29596
rect 3724 28627 3892 28644
rect 3724 28575 3726 28627
rect 3778 28588 3892 28627
rect 3948 28642 4004 30044
rect 4732 30102 4734 30154
rect 4786 30102 4788 30154
rect 4732 29988 4788 30102
rect 4620 29540 4676 29550
rect 4732 29540 4788 29932
rect 5068 30158 5070 30210
rect 5122 30158 5124 30210
rect 5068 29876 5124 30158
rect 5068 29810 5124 29820
rect 5292 30100 5348 30942
rect 5404 31220 5460 31230
rect 5404 30996 5460 31164
rect 5404 30902 5460 30940
rect 5516 30884 5572 31726
rect 5740 31778 5796 31892
rect 5740 31726 5742 31778
rect 5794 31726 5796 31778
rect 5740 31714 5796 31726
rect 6020 31668 6076 31678
rect 5852 31666 6076 31668
rect 5852 31614 6022 31666
rect 6074 31614 6076 31666
rect 5852 31612 6076 31614
rect 5684 31108 5740 31118
rect 5684 31014 5740 31052
rect 5516 30818 5572 30828
rect 5852 30996 5908 31612
rect 6020 31602 6076 31612
rect 6188 31220 6244 31892
rect 7084 31780 7140 32510
rect 7084 31714 7140 31724
rect 7420 32525 7422 32577
rect 7474 32525 7476 32577
rect 6636 31666 6692 31678
rect 6636 31614 6638 31666
rect 6690 31614 6692 31666
rect 6636 31332 6692 31614
rect 5292 29764 5348 30044
rect 5292 29698 5348 29708
rect 5628 30210 5684 30222
rect 5628 30158 5630 30210
rect 5682 30158 5684 30210
rect 5628 29652 5684 30158
rect 5740 30212 5796 30222
rect 5852 30212 5908 30940
rect 5964 31164 6244 31220
rect 6300 31276 6692 31332
rect 6300 31220 6356 31276
rect 5964 30660 6020 31164
rect 6188 30996 6244 31006
rect 6300 30996 6356 31164
rect 7308 31108 7364 31118
rect 7420 31108 7476 32525
rect 9100 32562 9156 32574
rect 9100 32510 9102 32562
rect 9154 32510 9156 32562
rect 7532 32450 7588 32462
rect 7532 32398 7534 32450
rect 7586 32398 7588 32450
rect 7532 32116 7588 32398
rect 7532 32050 7588 32060
rect 9100 32116 9156 32510
rect 9100 32050 9156 32060
rect 8540 31892 8596 31902
rect 8540 31798 8596 31836
rect 7308 31106 7476 31108
rect 7308 31054 7310 31106
rect 7362 31054 7476 31106
rect 7308 31052 7476 31054
rect 7308 31042 7364 31052
rect 6188 30994 6356 30996
rect 6188 30942 6190 30994
rect 6242 30942 6356 30994
rect 6188 30940 6356 30942
rect 7064 30996 7120 31006
rect 6188 30930 6244 30940
rect 7064 30902 7120 30940
rect 5964 30604 6132 30660
rect 5852 30156 5964 30212
rect 5740 30042 5796 30156
rect 5908 30154 5964 30156
rect 5908 30102 5910 30154
rect 5962 30102 5964 30154
rect 5908 30090 5964 30102
rect 5740 29990 5742 30042
rect 5794 29990 5796 30042
rect 5740 29978 5796 29990
rect 5628 29586 5684 29596
rect 4620 29538 4788 29540
rect 4620 29486 4622 29538
rect 4674 29486 4788 29538
rect 4620 29484 4788 29486
rect 4620 29474 4676 29484
rect 5292 29426 5348 29438
rect 5292 29374 5294 29426
rect 5346 29374 5348 29426
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4844 28756 4900 28766
rect 3948 28590 3950 28642
rect 4002 28590 4004 28642
rect 3778 28575 3780 28588
rect 3948 28578 4004 28590
rect 4060 28644 4116 28654
rect 4284 28644 4340 28654
rect 4116 28642 4340 28644
rect 4116 28590 4286 28642
rect 4338 28590 4340 28642
rect 4116 28588 4340 28590
rect 3724 28563 3780 28575
rect 2716 28466 2772 28476
rect 2940 28474 2996 28486
rect 2940 28422 2942 28474
rect 2994 28422 2996 28474
rect 3612 28466 3668 28476
rect 1932 27858 2100 27860
rect 1932 27806 1934 27858
rect 1986 27806 2100 27858
rect 2156 27916 2772 27972
rect 2156 27902 2212 27916
rect 2156 27850 2158 27902
rect 2210 27850 2212 27902
rect 2156 27838 2212 27850
rect 2716 27858 2772 27916
rect 1932 27804 2100 27806
rect 2716 27806 2718 27858
rect 2770 27806 2772 27858
rect 1932 26180 1988 27804
rect 2716 27794 2772 27806
rect 2940 27870 2996 28422
rect 2940 27858 3015 27870
rect 2940 27806 2961 27858
rect 3013 27806 3015 27858
rect 2940 27804 3015 27806
rect 2268 27746 2324 27758
rect 2268 27694 2270 27746
rect 2322 27694 2324 27746
rect 2268 27188 2324 27694
rect 2959 27636 3015 27804
rect 3836 27860 3892 27898
rect 3836 27794 3892 27804
rect 4060 27858 4116 28588
rect 4284 28578 4340 28588
rect 4060 27806 4062 27858
rect 4114 27806 4116 27858
rect 4060 27794 4116 27806
rect 4284 27860 4340 27870
rect 2604 27580 3015 27636
rect 2380 27188 2436 27198
rect 2268 27186 2436 27188
rect 2268 27134 2382 27186
rect 2434 27134 2436 27186
rect 2268 27132 2436 27134
rect 2380 27122 2436 27132
rect 2604 26852 2660 27580
rect 4284 27188 4340 27804
rect 4844 27858 4900 28700
rect 5292 28644 5348 29374
rect 5964 28868 6020 28878
rect 5740 28756 5796 28766
rect 5740 28662 5796 28700
rect 5964 28642 6020 28812
rect 5292 28578 5348 28588
rect 5572 28586 5628 28598
rect 5572 28534 5574 28586
rect 5626 28534 5628 28586
rect 5572 28084 5628 28534
rect 5964 28590 5966 28642
rect 6018 28590 6020 28642
rect 5964 28308 6020 28590
rect 5964 28242 6020 28252
rect 5572 28028 6020 28084
rect 4844 27806 4846 27858
rect 4898 27806 4900 27858
rect 4844 27794 4900 27806
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4788 27242 4844 27254
rect 4788 27190 4790 27242
rect 4842 27190 4844 27242
rect 4284 27186 4676 27188
rect 4284 27134 4286 27186
rect 4338 27134 4676 27186
rect 4284 27132 4676 27134
rect 4284 27122 4340 27132
rect 4620 27074 4676 27132
rect 4620 27022 4622 27074
rect 4674 27022 4676 27074
rect 4620 27010 4676 27022
rect 4788 27076 4844 27190
rect 5964 27188 6020 28028
rect 6076 27748 6132 30604
rect 6188 30324 6244 30334
rect 6188 29876 6244 30268
rect 6300 30210 6356 30222
rect 6300 30158 6302 30210
rect 6354 30158 6356 30210
rect 6300 30100 6356 30158
rect 6300 30034 6356 30044
rect 6860 30210 6916 30222
rect 6860 30158 6862 30210
rect 6914 30158 6916 30210
rect 6860 29876 6916 30158
rect 6188 29820 6356 29876
rect 6300 28586 6356 29820
rect 6860 29810 6916 29820
rect 6972 30212 7028 30222
rect 7532 30210 7588 30222
rect 6300 28534 6302 28586
rect 6354 28534 6356 28586
rect 6076 27682 6132 27692
rect 6188 28308 6244 28318
rect 6188 27524 6244 28252
rect 5852 27132 6020 27188
rect 6076 27468 6244 27524
rect 4788 27010 4844 27020
rect 5628 27076 5684 27086
rect 5628 26982 5684 27020
rect 2604 26786 2660 26796
rect 5404 26852 5460 26862
rect 3052 26305 3108 26317
rect 2716 26290 2772 26302
rect 2716 26238 2718 26290
rect 2770 26238 2772 26290
rect 2716 26180 2772 26238
rect 1932 26124 2772 26180
rect 3052 26253 3054 26305
rect 3106 26253 3108 26305
rect 1820 25394 1876 25406
rect 1820 25342 1822 25394
rect 1874 25342 1876 25394
rect 1820 24724 1876 25342
rect 1820 24658 1876 24668
rect 2268 24724 2324 24734
rect 1596 23938 1652 23950
rect 1596 23886 1598 23938
rect 1650 23886 1652 23938
rect 1596 21586 1652 23886
rect 2268 22596 2324 24668
rect 2380 23938 2436 23950
rect 2380 23886 2382 23938
rect 2434 23886 2436 23938
rect 2380 23378 2436 23886
rect 2380 23326 2382 23378
rect 2434 23326 2436 23378
rect 2380 23314 2436 23326
rect 2492 23380 2548 26124
rect 3052 25844 3108 26253
rect 5012 26292 5068 26302
rect 5180 26292 5236 26302
rect 5012 26290 5180 26292
rect 5012 26238 5014 26290
rect 5066 26238 5180 26290
rect 5012 26236 5180 26238
rect 5012 26226 5068 26236
rect 5180 26198 5236 26236
rect 5404 26290 5460 26796
rect 5684 26404 5740 26414
rect 5852 26404 5908 27132
rect 6076 27035 6132 27468
rect 6076 26983 6078 27035
rect 6130 26983 6132 27035
rect 6300 27074 6356 28534
rect 6300 27022 6302 27074
rect 6354 27022 6356 27074
rect 6300 27010 6356 27022
rect 6636 29652 6692 29662
rect 6076 26971 6132 26983
rect 6412 26906 6468 26918
rect 6412 26854 6414 26906
rect 6466 26854 6468 26906
rect 6412 26628 6468 26854
rect 6468 26572 6580 26628
rect 6412 26562 6468 26572
rect 5684 26402 5908 26404
rect 5684 26350 5686 26402
rect 5738 26350 5908 26402
rect 5684 26348 5908 26350
rect 5684 26338 5740 26348
rect 5404 26238 5406 26290
rect 5458 26238 5460 26290
rect 5404 26226 5460 26238
rect 5964 26290 6020 26302
rect 5964 26238 5966 26290
rect 6018 26238 6020 26290
rect 3164 26180 3220 26190
rect 3164 26086 3220 26124
rect 3724 26180 3780 26190
rect 3052 25788 3556 25844
rect 3500 24836 3556 25788
rect 3724 25618 3780 26124
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 3724 25566 3726 25618
rect 3778 25566 3780 25618
rect 3724 25554 3780 25566
rect 4508 25508 4564 25518
rect 4508 25414 4564 25452
rect 5852 25506 5908 25518
rect 5852 25454 5854 25506
rect 5906 25454 5908 25506
rect 5740 25396 5796 25406
rect 5404 25284 5460 25294
rect 4844 25060 4900 25070
rect 3500 24770 3556 24780
rect 3948 24836 4004 24846
rect 2828 24724 2884 24762
rect 3948 24742 4004 24780
rect 4564 24836 4620 24846
rect 4564 24742 4620 24780
rect 2828 24658 2884 24668
rect 3704 24724 3760 24734
rect 3704 24722 3780 24724
rect 3704 24670 3706 24722
rect 3758 24670 3780 24722
rect 3704 24658 3780 24670
rect 4844 24722 4900 25004
rect 4844 24670 4846 24722
rect 4898 24670 4900 24722
rect 4844 24658 4900 24670
rect 4956 24836 5012 24846
rect 5404 24836 5460 25228
rect 3724 23716 3780 24658
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4284 23826 4340 23838
rect 4284 23774 4286 23826
rect 4338 23774 4340 23826
rect 3724 23660 3892 23716
rect 2492 23314 2548 23324
rect 3612 23322 3668 23334
rect 3612 23270 3614 23322
rect 3666 23270 3668 23322
rect 2716 23156 2772 23166
rect 2716 23062 2772 23100
rect 3500 23154 3556 23166
rect 3500 23102 3502 23154
rect 3554 23102 3556 23154
rect 3500 22820 3556 23102
rect 3612 23156 3668 23270
rect 3612 23090 3668 23100
rect 3836 23181 3892 23660
rect 3836 23129 3838 23181
rect 3890 23129 3892 23181
rect 3500 22764 3668 22820
rect 3444 22596 3500 22606
rect 2268 22540 3220 22596
rect 2268 22370 2324 22540
rect 2268 22318 2270 22370
rect 2322 22318 2324 22370
rect 2268 22306 2324 22318
rect 2380 22370 2436 22382
rect 2380 22318 2382 22370
rect 2434 22318 2436 22370
rect 2380 22260 2436 22318
rect 3052 22370 3108 22382
rect 3052 22318 3054 22370
rect 3106 22318 3108 22370
rect 2660 22260 2716 22270
rect 2380 22194 2436 22204
rect 2604 22258 2716 22260
rect 2604 22206 2662 22258
rect 2714 22206 2716 22258
rect 2604 22194 2716 22206
rect 1596 21534 1598 21586
rect 1650 21534 1652 21586
rect 1596 20018 1652 21534
rect 2380 21476 2436 21486
rect 2044 21474 2436 21476
rect 2044 21422 2382 21474
rect 2434 21422 2436 21474
rect 2044 21420 2436 21422
rect 2044 21026 2100 21420
rect 2380 21410 2436 21420
rect 2604 21252 2660 22194
rect 3052 21812 3108 22318
rect 3164 22370 3220 22540
rect 3444 22502 3500 22540
rect 3164 22318 3166 22370
rect 3218 22318 3220 22370
rect 3164 22306 3220 22318
rect 3052 21746 3108 21756
rect 3276 21252 3332 21262
rect 2604 21196 2772 21252
rect 2044 20974 2046 21026
rect 2098 20974 2100 21026
rect 2044 20962 2100 20974
rect 2604 20916 2660 20926
rect 2604 20822 2660 20860
rect 2380 20804 2436 20814
rect 2380 20710 2436 20748
rect 2716 20787 2772 21196
rect 2716 20735 2718 20787
rect 2770 20735 2772 20787
rect 3052 21028 3108 21038
rect 3052 20802 3108 20972
rect 3052 20750 3054 20802
rect 3106 20750 3108 20802
rect 3052 20738 3108 20750
rect 2716 20692 2772 20735
rect 2716 20626 2772 20636
rect 3276 20188 3332 21196
rect 3612 21028 3668 22764
rect 3836 22260 3892 23129
rect 3948 23492 4004 23502
rect 3948 22370 4004 23436
rect 4284 23492 4340 23774
rect 4284 23426 4340 23436
rect 4172 23154 4228 23166
rect 4172 23102 4174 23154
rect 4226 23102 4228 23154
rect 4172 22484 4228 23102
rect 4844 23154 4900 23166
rect 4844 23102 4846 23154
rect 4898 23102 4900 23154
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4284 22484 4340 22494
rect 4172 22482 4340 22484
rect 4172 22430 4286 22482
rect 4338 22430 4340 22482
rect 4172 22428 4340 22430
rect 4284 22418 4340 22428
rect 3948 22318 3950 22370
rect 4002 22318 4004 22370
rect 3948 22306 4004 22318
rect 4172 22326 4228 22338
rect 3836 22194 3892 22204
rect 4172 22274 4174 22326
rect 4226 22274 4228 22326
rect 4172 22148 4228 22274
rect 4676 22260 4732 22270
rect 4676 22166 4732 22204
rect 4172 22082 4228 22092
rect 3388 20972 3668 21028
rect 3388 20802 3444 20972
rect 3388 20750 3390 20802
rect 3442 20750 3444 20802
rect 3388 20738 3444 20750
rect 3500 20804 3556 20814
rect 3500 20634 3556 20748
rect 3500 20582 3502 20634
rect 3554 20582 3556 20634
rect 3500 20570 3556 20582
rect 3276 20132 3556 20188
rect 1596 19966 1598 20018
rect 1650 19966 1652 20018
rect 1596 18452 1652 19966
rect 2380 19908 2436 19918
rect 2044 19906 2436 19908
rect 2044 19854 2382 19906
rect 2434 19854 2436 19906
rect 2044 19852 2436 19854
rect 2044 19458 2100 19852
rect 2380 19842 2436 19852
rect 2044 19406 2046 19458
rect 2098 19406 2100 19458
rect 2044 19394 2100 19406
rect 2380 19460 2436 19470
rect 2380 19234 2436 19404
rect 2380 19182 2382 19234
rect 2434 19182 2436 19234
rect 2380 19170 2436 19182
rect 3052 18564 3108 18574
rect 1596 17666 1652 18396
rect 2044 18452 2100 18462
rect 2044 18358 2100 18396
rect 3052 18450 3108 18508
rect 3052 18398 3054 18450
rect 3106 18398 3108 18450
rect 3052 18386 3108 18398
rect 3500 18450 3556 20132
rect 3612 20020 3668 20972
rect 4284 21476 4340 21486
rect 4284 21028 4340 21420
rect 4844 21476 4900 23102
rect 4956 22370 5012 24780
rect 5068 24834 5460 24836
rect 5068 24782 5406 24834
rect 5458 24782 5460 24834
rect 5068 24780 5460 24782
rect 5068 24722 5124 24780
rect 5404 24770 5460 24780
rect 5068 24670 5070 24722
rect 5122 24670 5124 24722
rect 5068 24658 5124 24670
rect 5628 23938 5684 23950
rect 5628 23886 5630 23938
rect 5682 23886 5684 23938
rect 5180 23492 5236 23502
rect 5068 23154 5124 23166
rect 5068 23102 5070 23154
rect 5122 23102 5124 23154
rect 5068 22596 5124 23102
rect 5068 22530 5124 22540
rect 4956 22318 4958 22370
rect 5010 22318 5012 22370
rect 4956 22148 5012 22318
rect 5180 22370 5236 23436
rect 5628 23492 5684 23886
rect 5628 23426 5684 23436
rect 5348 23268 5404 23278
rect 5348 23174 5404 23212
rect 5516 23268 5572 23278
rect 5180 22318 5182 22370
rect 5234 22318 5236 22370
rect 5180 22306 5236 22318
rect 4956 22082 5012 22092
rect 5292 22260 5348 22270
rect 5292 21586 5348 22204
rect 5292 21534 5294 21586
rect 5346 21534 5348 21586
rect 5292 21522 5348 21534
rect 5516 21586 5572 23212
rect 5740 23156 5796 25340
rect 5852 24836 5908 25454
rect 5964 25338 6020 26238
rect 6188 26180 6244 26190
rect 6188 25479 6244 26124
rect 6188 25427 6190 25479
rect 6242 25427 6244 25479
rect 6188 25415 6244 25427
rect 6300 26066 6356 26078
rect 6300 26014 6302 26066
rect 6354 26014 6356 26066
rect 5964 25286 5966 25338
rect 6018 25286 6020 25338
rect 5964 25274 6020 25286
rect 6076 25284 6132 25294
rect 5852 24770 5908 24780
rect 5516 21534 5518 21586
rect 5570 21534 5572 21586
rect 5516 21522 5572 21534
rect 5628 23154 5796 23156
rect 5628 23102 5742 23154
rect 5794 23102 5796 23154
rect 5628 23100 5796 23102
rect 4844 21410 4900 21420
rect 5180 21476 5236 21486
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4284 20962 4340 20972
rect 3724 20916 3780 20926
rect 3724 20775 3780 20860
rect 3724 20723 3726 20775
rect 3778 20723 3780 20775
rect 3724 20711 3780 20723
rect 4060 20802 4116 20814
rect 4060 20750 4062 20802
rect 4114 20750 4116 20802
rect 4060 20692 4116 20750
rect 4956 20802 5012 20814
rect 4956 20750 4958 20802
rect 5010 20750 5012 20802
rect 4676 20692 4732 20702
rect 4060 20690 4732 20692
rect 4060 20638 4678 20690
rect 4730 20638 4732 20690
rect 4060 20636 4732 20638
rect 4060 20020 4116 20636
rect 4676 20626 4732 20636
rect 4956 20692 5012 20750
rect 5180 20802 5236 21420
rect 5628 21140 5684 23100
rect 5740 23090 5796 23100
rect 5964 24050 6020 24062
rect 5964 23998 5966 24050
rect 6018 23998 6020 24050
rect 5852 22372 5908 22382
rect 5852 22278 5908 22316
rect 5964 21476 6020 23998
rect 6076 23899 6132 25228
rect 6076 23847 6078 23899
rect 6130 23847 6132 23899
rect 6188 25060 6244 25070
rect 6188 23940 6244 25004
rect 6300 24948 6356 26014
rect 6412 25506 6468 25518
rect 6412 25454 6414 25506
rect 6466 25454 6468 25506
rect 6412 25396 6468 25454
rect 6412 25330 6468 25340
rect 6524 25060 6580 26572
rect 6636 25396 6692 29596
rect 6972 28644 7028 30156
rect 7196 30166 7252 30178
rect 7196 30114 7198 30166
rect 7250 30114 7252 30166
rect 7084 30100 7140 30110
rect 7084 30042 7140 30044
rect 7084 29990 7086 30042
rect 7138 29990 7140 30042
rect 7084 29978 7140 29990
rect 7196 29764 7252 30114
rect 7532 30158 7534 30210
rect 7586 30158 7588 30210
rect 7532 29988 7588 30158
rect 8316 30212 8372 30222
rect 8316 30118 8372 30156
rect 9100 30210 9156 30222
rect 9100 30158 9102 30210
rect 9154 30158 9156 30210
rect 7532 29922 7588 29932
rect 7868 29986 7924 29998
rect 7868 29934 7870 29986
rect 7922 29934 7924 29986
rect 7196 29698 7252 29708
rect 7868 29764 7924 29934
rect 9100 29876 9156 30158
rect 9100 29810 9156 29820
rect 7868 29698 7924 29708
rect 9044 29652 9100 29662
rect 9212 29652 9268 34636
rect 9380 34692 9436 34702
rect 9380 34598 9436 34636
rect 9604 34468 9660 34478
rect 9772 34468 9828 37214
rect 9996 36596 10052 38444
rect 10108 38164 10164 38174
rect 10108 38050 10164 38108
rect 10108 37998 10110 38050
rect 10162 37998 10164 38050
rect 10108 37986 10164 37998
rect 10220 37266 10276 38556
rect 10612 38276 10668 38286
rect 10612 38182 10668 38220
rect 11676 38274 11732 39788
rect 11788 40402 11844 40414
rect 11788 40350 11790 40402
rect 11842 40350 11844 40402
rect 11788 39396 11844 40350
rect 11788 39330 11844 39340
rect 11788 39172 11844 39182
rect 11788 39058 11844 39116
rect 11788 39006 11790 39058
rect 11842 39006 11844 39058
rect 11788 38994 11844 39006
rect 11676 38222 11678 38274
rect 11730 38222 11732 38274
rect 10332 38052 10388 38062
rect 10332 37958 10388 37996
rect 11676 38052 11732 38222
rect 11676 37986 11732 37996
rect 11900 37604 11956 40796
rect 12460 40628 12516 40796
rect 12236 40572 12516 40628
rect 12572 40628 12628 40638
rect 12012 39732 12068 39742
rect 12012 39583 12068 39676
rect 12012 39531 12014 39583
rect 12066 39531 12068 39583
rect 12012 39519 12068 39531
rect 12124 39562 12180 39574
rect 12124 39510 12126 39562
rect 12178 39510 12180 39562
rect 12124 39060 12180 39510
rect 12124 38994 12180 39004
rect 12124 38834 12180 38846
rect 12124 38782 12126 38834
rect 12178 38782 12180 38834
rect 12012 38052 12068 38062
rect 12124 38052 12180 38782
rect 12012 38050 12180 38052
rect 12012 37998 12014 38050
rect 12066 37998 12180 38050
rect 12012 37996 12180 37998
rect 12012 37986 12068 37996
rect 11900 37538 11956 37548
rect 10220 37214 10222 37266
rect 10274 37214 10276 37266
rect 10220 37202 10276 37214
rect 11004 37156 11060 37166
rect 11004 37154 11284 37156
rect 11004 37102 11006 37154
rect 11058 37102 11284 37154
rect 11004 37100 11284 37102
rect 11004 37090 11060 37100
rect 11228 36708 11284 37100
rect 12124 37044 12180 37996
rect 12124 36978 12180 36988
rect 12236 37492 12292 40572
rect 12572 39590 12628 40572
rect 12684 40404 12740 41244
rect 12796 41074 12852 41086
rect 12796 41022 12798 41074
rect 12850 41022 12852 41074
rect 12796 40740 12852 41022
rect 12796 40674 12852 40684
rect 13244 40740 13300 40750
rect 13244 40458 13300 40684
rect 13356 40628 13412 42700
rect 13468 42754 13524 42766
rect 13468 42702 13470 42754
rect 13522 42702 13524 42754
rect 13468 42644 13524 42702
rect 13468 42578 13524 42588
rect 13580 42756 13636 42766
rect 13580 42026 13636 42700
rect 13580 41974 13582 42026
rect 13634 41974 13636 42026
rect 14140 42026 14196 43148
rect 14364 42766 14420 43708
rect 14588 43988 14644 43998
rect 14344 42754 14420 42766
rect 14344 42702 14346 42754
rect 14398 42702 14420 42754
rect 14344 42700 14420 42702
rect 14476 43652 14532 43662
rect 14476 43428 14532 43596
rect 14344 42690 14400 42700
rect 14476 42644 14532 43372
rect 14588 42978 14644 43932
rect 14812 43538 14868 44380
rect 14812 43486 14814 43538
rect 14866 43486 14868 43538
rect 14812 43474 14868 43486
rect 14924 44322 14980 45838
rect 15148 45108 15204 46284
rect 15708 45890 15764 45902
rect 15708 45838 15710 45890
rect 15762 45838 15764 45890
rect 15596 45220 15652 45230
rect 15596 45150 15652 45164
rect 15372 45108 15428 45118
rect 15148 45106 15428 45108
rect 15148 45054 15374 45106
rect 15426 45054 15428 45106
rect 15596 45098 15598 45150
rect 15650 45098 15652 45150
rect 15596 45086 15652 45098
rect 15148 45052 15428 45054
rect 14924 44270 14926 44322
rect 14978 44270 14980 44322
rect 14924 43540 14980 44270
rect 15372 44100 15428 45052
rect 15708 44994 15764 45838
rect 17612 45780 17668 46622
rect 17612 45686 17668 45724
rect 17836 46564 17892 46574
rect 15708 44942 15710 44994
rect 15762 44942 15764 44994
rect 15708 44930 15764 44942
rect 16940 45106 16996 45118
rect 16940 45054 16942 45106
rect 16994 45054 16996 45106
rect 16940 44996 16996 45054
rect 17724 45108 17780 45118
rect 17724 45014 17780 45052
rect 17836 45106 17892 46508
rect 18172 46452 18228 46462
rect 17948 45890 18004 45902
rect 17948 45838 17950 45890
rect 18002 45838 18004 45890
rect 17948 45332 18004 45838
rect 17948 45266 18004 45276
rect 18172 45444 18228 46396
rect 18396 45780 18452 45790
rect 17836 45054 17838 45106
rect 17890 45054 17892 45106
rect 16940 44940 17332 44996
rect 16772 44884 16828 44894
rect 16772 44882 16996 44884
rect 16772 44830 16774 44882
rect 16826 44830 16996 44882
rect 16772 44828 16996 44830
rect 16772 44818 16828 44828
rect 16828 44660 16884 44670
rect 15820 44436 15876 44446
rect 15820 44342 15876 44380
rect 16156 44322 16212 44334
rect 15372 44034 15428 44044
rect 15932 44278 15988 44290
rect 15932 44226 15934 44278
rect 15986 44226 15988 44278
rect 15932 43988 15988 44226
rect 16156 44270 16158 44322
rect 16210 44270 16212 44322
rect 16156 44100 16212 44270
rect 16156 44034 16212 44044
rect 16268 44212 16324 44222
rect 15932 43922 15988 43932
rect 14924 43474 14980 43484
rect 16044 43540 16100 43550
rect 14588 42926 14590 42978
rect 14642 42926 14644 42978
rect 14588 42914 14644 42926
rect 16044 42978 16100 43484
rect 16044 42926 16046 42978
rect 16098 42926 16100 42978
rect 16044 42756 16100 42926
rect 14476 42578 14532 42588
rect 15372 42726 15428 42738
rect 15372 42674 15374 42726
rect 15426 42674 15428 42726
rect 16044 42690 16100 42700
rect 16156 43316 16212 43326
rect 15372 42644 15428 42674
rect 15372 42578 15428 42588
rect 13580 41962 13636 41974
rect 13692 41998 13748 42010
rect 13692 41972 13694 41998
rect 13746 41972 13748 41998
rect 13692 41906 13748 41916
rect 13916 41998 13972 42010
rect 13916 41972 13918 41998
rect 13970 41972 13972 41998
rect 14140 41974 14142 42026
rect 14194 41974 14196 42026
rect 16156 42026 16212 43260
rect 16268 42644 16324 44156
rect 16716 44100 16772 44110
rect 16268 42578 16324 42588
rect 16604 44098 16772 44100
rect 16604 44046 16718 44098
rect 16770 44046 16772 44098
rect 16604 44044 16772 44046
rect 16604 43652 16660 44044
rect 16716 44034 16772 44044
rect 15596 42005 15652 42017
rect 14140 41972 14196 41974
rect 15372 41972 15428 41982
rect 14140 41916 15092 41972
rect 13916 41906 13972 41916
rect 13468 41860 13524 41870
rect 13468 41153 13524 41804
rect 14420 41746 14476 41758
rect 14420 41694 14422 41746
rect 14474 41694 14476 41746
rect 13468 41101 13470 41153
rect 13522 41101 13524 41153
rect 13468 41089 13524 41101
rect 13804 41188 13860 41198
rect 14420 41188 14476 41694
rect 14420 41146 14618 41188
rect 13804 41101 13806 41132
rect 13858 41101 13860 41132
rect 13804 41089 13860 41101
rect 14308 41130 14364 41142
rect 14420 41132 14564 41146
rect 14308 41078 14310 41130
rect 14362 41078 14364 41130
rect 14308 41076 14364 41078
rect 14562 41094 14564 41132
rect 14616 41094 14618 41146
rect 15036 41186 15092 41916
rect 15036 41134 15038 41186
rect 15090 41134 15092 41186
rect 15036 41122 15092 41134
rect 15372 41142 15428 41916
rect 15596 41953 15598 42005
rect 15650 41953 15652 42005
rect 15596 41636 15652 41953
rect 15708 41998 15764 42010
rect 15708 41946 15710 41998
rect 15762 41946 15764 41998
rect 15708 41860 15764 41946
rect 15708 41794 15764 41804
rect 15932 41998 15988 42010
rect 15932 41946 15934 41998
rect 15986 41946 15988 41998
rect 16156 41974 16158 42026
rect 16210 41974 16212 42026
rect 16156 41962 16212 41974
rect 16436 41972 16492 41982
rect 15596 41570 15652 41580
rect 15932 41412 15988 41946
rect 16436 41878 16492 41916
rect 15932 41346 15988 41356
rect 16156 41748 16212 41758
rect 14308 41020 14420 41076
rect 13356 40572 13524 40628
rect 12908 40404 12964 40414
rect 12684 40348 12908 40404
rect 13244 40406 13246 40458
rect 13298 40406 13300 40458
rect 13244 40394 13300 40406
rect 12908 40310 12964 40348
rect 13132 40290 13188 40302
rect 13468 40292 13524 40572
rect 13132 40238 13134 40290
rect 13186 40238 13188 40290
rect 12404 39562 12460 39574
rect 12404 39510 12406 39562
rect 12458 39510 12460 39562
rect 12572 39538 12574 39590
rect 12626 39538 12628 39590
rect 12572 39526 12628 39538
rect 13020 40068 13076 40078
rect 12404 39508 12460 39510
rect 12852 39508 12908 39518
rect 12404 39452 12516 39508
rect 12460 39284 12516 39452
rect 12684 39506 12908 39508
rect 12684 39454 12854 39506
rect 12906 39454 12908 39506
rect 12684 39452 12908 39454
rect 12460 39228 12628 39284
rect 12572 39002 12628 39228
rect 12460 38948 12516 38958
rect 12572 38950 12574 39002
rect 12626 38950 12628 39002
rect 12572 38938 12628 38950
rect 12460 38834 12516 38892
rect 12460 38782 12462 38834
rect 12514 38782 12516 38834
rect 12460 38770 12516 38782
rect 12348 38052 12404 38062
rect 12348 37958 12404 37996
rect 12572 38050 12628 38062
rect 12572 37998 12574 38050
rect 12626 37998 12628 38050
rect 11452 36708 11508 36718
rect 11228 36706 11508 36708
rect 11228 36654 11454 36706
rect 11506 36654 11508 36706
rect 11228 36652 11508 36654
rect 11452 36642 11508 36652
rect 9884 36594 10052 36596
rect 9884 36542 9998 36594
rect 10050 36542 10052 36594
rect 9884 36540 10052 36542
rect 9884 35754 9940 36540
rect 9996 36530 10052 36540
rect 9884 35702 9886 35754
rect 9938 35702 9940 35754
rect 10780 36484 10836 36494
rect 9884 35690 9940 35702
rect 10108 35726 10164 35738
rect 10108 35674 10110 35726
rect 10162 35674 10164 35726
rect 10108 35140 10164 35674
rect 10332 35726 10388 35738
rect 10332 35674 10334 35726
rect 10386 35674 10388 35726
rect 10108 35084 10276 35140
rect 10108 34916 10164 34926
rect 10108 34822 10164 34860
rect 9940 34692 9996 34702
rect 10220 34692 10276 35084
rect 9940 34690 10052 34692
rect 9940 34638 9942 34690
rect 9994 34638 10052 34690
rect 9940 34626 10052 34638
rect 9996 34468 10052 34626
rect 9772 34412 9940 34468
rect 9604 34242 9660 34412
rect 9604 34190 9606 34242
rect 9658 34190 9660 34242
rect 9604 34178 9660 34190
rect 9884 34186 9940 34412
rect 9996 34402 10052 34412
rect 10108 34636 10276 34692
rect 9884 34134 9886 34186
rect 9938 34134 9940 34186
rect 9884 34132 9940 34134
rect 9884 34056 9940 34076
rect 10108 34158 10164 34636
rect 10108 34106 10110 34158
rect 10162 34106 10164 34158
rect 10108 33796 10164 34106
rect 9996 33740 10164 33796
rect 10332 34158 10388 35674
rect 10500 35714 10556 35726
rect 10500 35662 10502 35714
rect 10554 35700 10556 35714
rect 10554 35662 10612 35700
rect 10500 35644 10612 35662
rect 10556 35588 10612 35644
rect 10332 34106 10334 34158
rect 10386 34106 10388 34158
rect 10444 34468 10500 34478
rect 10444 34186 10500 34412
rect 10444 34134 10446 34186
rect 10498 34134 10500 34186
rect 10444 34122 10500 34134
rect 9996 33460 10052 33740
rect 10164 33572 10220 33582
rect 10164 33478 10220 33516
rect 10332 33572 10388 34106
rect 9996 33394 10052 33404
rect 9660 33348 9716 33358
rect 9660 33254 9716 33292
rect 10332 32788 10388 33516
rect 10444 33348 10500 33358
rect 10444 33266 10446 33292
rect 10498 33266 10500 33292
rect 10444 33254 10500 33266
rect 10332 32722 10388 32732
rect 9044 29650 9268 29652
rect 9044 29598 9046 29650
rect 9098 29598 9268 29650
rect 9044 29596 9268 29598
rect 9044 29586 9100 29596
rect 7532 29453 7588 29465
rect 7532 29401 7534 29453
rect 7586 29401 7588 29453
rect 7532 29316 7588 29401
rect 8204 29441 8260 29453
rect 8204 29389 8206 29441
rect 8258 29389 8260 29441
rect 8092 29316 8148 29326
rect 7532 29250 7588 29260
rect 7756 29314 8148 29316
rect 7756 29262 8094 29314
rect 8146 29262 8148 29314
rect 7756 29260 8148 29262
rect 7756 28754 7812 29260
rect 8092 29250 8148 29260
rect 8204 28980 8260 29389
rect 8540 29426 8596 29438
rect 8540 29374 8542 29426
rect 8594 29374 8596 29426
rect 8540 29316 8596 29374
rect 9212 29428 9268 29596
rect 9212 29362 9268 29372
rect 9324 32564 9380 32574
rect 9324 31778 9380 32508
rect 9996 32564 10052 32574
rect 10556 32564 10612 35532
rect 10780 34142 10836 36428
rect 11788 36484 11844 36494
rect 12068 36484 12124 36494
rect 11788 36482 12124 36484
rect 11788 36430 11790 36482
rect 11842 36430 12070 36482
rect 12122 36430 12124 36482
rect 11788 36428 12124 36430
rect 12236 36484 12292 37436
rect 12460 37604 12516 37614
rect 12236 36447 12348 36484
rect 12236 36428 12294 36447
rect 11788 36418 11844 36428
rect 12068 36418 12124 36428
rect 12292 36395 12294 36428
rect 12346 36395 12348 36447
rect 12292 36383 12348 36395
rect 12460 36260 12516 37548
rect 12572 37380 12628 37998
rect 12572 37314 12628 37324
rect 12236 36204 12516 36260
rect 12572 36484 12628 36494
rect 12572 36402 12574 36428
rect 12626 36402 12628 36428
rect 11116 35812 11172 35822
rect 10948 35588 11004 35598
rect 10948 35494 11004 35532
rect 10892 34914 10948 34926
rect 10892 34862 10894 34914
rect 10946 34862 10948 34914
rect 10892 34356 10948 34862
rect 10892 34290 10948 34300
rect 11116 34186 11172 35756
rect 12236 35754 12292 36204
rect 12572 36148 12628 36402
rect 12236 35702 12238 35754
rect 12290 35702 12292 35754
rect 11956 35476 12012 35486
rect 11956 35474 12068 35476
rect 11956 35422 11958 35474
rect 12010 35422 12068 35474
rect 11956 35410 12068 35422
rect 10780 34130 10892 34142
rect 10780 34078 10838 34130
rect 10890 34078 10892 34130
rect 11116 34134 11118 34186
rect 11170 34134 11172 34186
rect 11676 34692 11732 34702
rect 11116 34122 11172 34134
rect 11284 34165 11340 34177
rect 11284 34132 11286 34165
rect 10780 34076 10892 34078
rect 10836 34066 10892 34076
rect 11228 34113 11286 34132
rect 11338 34113 11340 34165
rect 11228 34076 11340 34113
rect 11564 34158 11620 34170
rect 11564 34106 11566 34158
rect 11618 34106 11620 34158
rect 11228 33796 11284 34076
rect 9996 32470 10052 32508
rect 10220 32508 10612 32564
rect 10668 33740 11284 33796
rect 10668 33460 10724 33740
rect 11564 33572 11620 34106
rect 11564 33506 11620 33516
rect 11676 34165 11732 34636
rect 11676 34113 11678 34165
rect 11730 34113 11732 34165
rect 11452 33460 11508 33470
rect 10668 33290 10724 33404
rect 10668 33238 10670 33290
rect 10722 33238 10724 33290
rect 9716 32452 9772 32462
rect 9716 32450 9828 32452
rect 9716 32398 9718 32450
rect 9770 32398 9828 32450
rect 9716 32386 9828 32398
rect 9660 32228 9716 32238
rect 9660 31890 9716 32172
rect 9660 31838 9662 31890
rect 9714 31838 9716 31890
rect 9660 31826 9716 31838
rect 9772 32116 9828 32386
rect 9324 31726 9326 31778
rect 9378 31726 9380 31778
rect 8540 29250 8596 29260
rect 7756 28702 7758 28754
rect 7810 28702 7812 28754
rect 7756 28690 7812 28702
rect 7868 28924 8260 28980
rect 6748 27860 6804 27870
rect 6748 27766 6804 27804
rect 6972 27076 7028 28588
rect 7252 28308 7308 28318
rect 7252 28082 7308 28252
rect 7252 28030 7254 28082
rect 7306 28030 7308 28082
rect 7252 28018 7308 28030
rect 7868 27970 7924 28924
rect 9212 28756 9268 28766
rect 7980 28644 8036 28654
rect 7980 28196 8036 28588
rect 7980 28140 8167 28196
rect 7868 27918 7870 27970
rect 7922 27918 7924 27970
rect 7868 27906 7924 27918
rect 8111 27914 8167 28140
rect 7084 27860 7140 27870
rect 8111 27862 8113 27914
rect 8165 27862 8167 27914
rect 8111 27850 8167 27862
rect 8988 27972 9044 27982
rect 8988 27858 9044 27916
rect 7084 27766 7140 27804
rect 8988 27806 8990 27858
rect 9042 27806 9044 27858
rect 8988 27794 9044 27806
rect 7084 27076 7140 27086
rect 6972 27074 7140 27076
rect 6972 27022 7086 27074
rect 7138 27022 7140 27074
rect 6972 27020 7140 27022
rect 7084 27010 7140 27020
rect 7868 27074 7924 27086
rect 7868 27022 7870 27074
rect 7922 27022 7924 27074
rect 7868 26908 7924 27022
rect 9212 26908 9268 28700
rect 9324 27860 9380 31726
rect 9772 31763 9828 32060
rect 9772 31711 9774 31763
rect 9826 31711 9828 31763
rect 9772 31699 9828 31711
rect 10108 31780 10164 31790
rect 10108 31686 10164 31724
rect 9548 29876 9604 29886
rect 9548 29314 9604 29820
rect 9660 29540 9716 29550
rect 9660 29470 9716 29484
rect 9660 29418 9662 29470
rect 9714 29418 9716 29470
rect 9660 29406 9716 29418
rect 9996 29426 10052 29438
rect 9548 29262 9550 29314
rect 9602 29262 9604 29314
rect 9548 29250 9604 29262
rect 9996 29374 9998 29426
rect 10050 29374 10052 29426
rect 9996 29316 10052 29374
rect 9996 28756 10052 29260
rect 10220 29092 10276 32508
rect 10668 32228 10724 33238
rect 10780 33458 11508 33460
rect 10780 33406 11454 33458
rect 11506 33406 11508 33458
rect 10780 33404 11508 33406
rect 10780 32562 10836 33404
rect 11452 33394 11508 33404
rect 11508 33320 11564 33328
rect 11116 33316 11564 33320
rect 10892 33290 10948 33302
rect 10892 33238 10894 33290
rect 10946 33238 10948 33290
rect 10892 32788 10948 33238
rect 11004 33290 11060 33302
rect 11004 33238 11006 33290
rect 11058 33238 11060 33290
rect 11004 33236 11060 33238
rect 11004 33170 11060 33180
rect 11116 33264 11510 33316
rect 11562 33264 11564 33316
rect 11116 32788 11172 33264
rect 11508 33252 11564 33264
rect 10892 32722 10948 32732
rect 11004 32732 11172 32788
rect 11676 32788 11732 34113
rect 11900 34132 11956 34142
rect 12012 34132 12068 35410
rect 12236 34804 12292 35702
rect 12460 36092 12628 36148
rect 12460 35754 12516 36092
rect 12684 35924 12740 39452
rect 12852 39442 12908 39452
rect 13020 39284 13076 40012
rect 12908 39228 13076 39284
rect 12908 38890 12964 39228
rect 12908 38838 12910 38890
rect 12962 38838 12964 38890
rect 12908 38826 12964 38838
rect 13132 38834 13188 40238
rect 13132 38782 13134 38834
rect 13186 38782 13188 38834
rect 13132 38770 13188 38782
rect 13356 40236 13524 40292
rect 13580 40402 13636 40414
rect 13580 40350 13582 40402
rect 13634 40350 13636 40402
rect 13356 38050 13412 40236
rect 13580 38836 13636 40350
rect 13916 40404 13972 40414
rect 14364 40404 14420 41020
rect 14562 40740 14618 41094
rect 15372 41090 15374 41142
rect 15426 41090 15428 41142
rect 14700 41076 14756 41086
rect 14700 41074 14980 41076
rect 14700 41022 14702 41074
rect 14754 41022 14980 41074
rect 14700 41020 14980 41022
rect 14700 41010 14756 41020
rect 14812 40740 14868 40750
rect 14562 40684 14756 40740
rect 14476 40404 14532 40414
rect 13916 40402 14196 40404
rect 13916 40350 13918 40402
rect 13970 40350 14196 40402
rect 13916 40348 14196 40350
rect 14364 40348 14476 40404
rect 13916 40338 13972 40348
rect 14140 39450 14196 40348
rect 14476 40310 14532 40348
rect 14252 40292 14308 40302
rect 14252 39618 14308 40236
rect 14700 39620 14756 40684
rect 14812 40402 14868 40684
rect 14812 40350 14814 40402
rect 14866 40350 14868 40402
rect 14812 40338 14868 40350
rect 14252 39566 14254 39618
rect 14306 39566 14308 39618
rect 14252 39554 14308 39566
rect 14644 39564 14756 39620
rect 14812 40234 14868 40246
rect 14812 40182 14814 40234
rect 14866 40182 14868 40234
rect 14812 39620 14868 40182
rect 14924 39844 14980 41020
rect 15372 40404 15428 41090
rect 15372 40338 15428 40348
rect 15484 41298 15540 41310
rect 15484 41246 15486 41298
rect 15538 41246 15540 41298
rect 15484 39844 15540 41246
rect 16044 41298 16100 41310
rect 16044 41246 16046 41298
rect 16098 41246 16100 41298
rect 15820 41076 15876 41086
rect 15820 40402 15876 41020
rect 16044 40628 16100 41246
rect 16156 41171 16212 41692
rect 16604 41636 16660 43596
rect 16716 43540 16772 43550
rect 16716 43446 16772 43484
rect 16604 41570 16660 41580
rect 16156 41119 16158 41171
rect 16210 41119 16212 41171
rect 16156 41107 16212 41119
rect 16492 41188 16548 41198
rect 16492 41094 16548 41132
rect 16828 41186 16884 44604
rect 16940 44324 16996 44828
rect 17276 44436 17332 44940
rect 17444 44882 17500 44894
rect 17836 44884 17892 45054
rect 17444 44830 17446 44882
rect 17498 44830 17500 44882
rect 17444 44660 17500 44830
rect 17444 44594 17500 44604
rect 17612 44828 17892 44884
rect 17948 45108 18004 45118
rect 17276 44380 17556 44436
rect 16940 44258 16996 44268
rect 17052 44322 17108 44334
rect 17052 44270 17054 44322
rect 17106 44270 17108 44322
rect 17052 43540 17108 44270
rect 17332 44210 17388 44222
rect 17332 44158 17334 44210
rect 17386 44158 17388 44210
rect 17332 43708 17388 44158
rect 17052 43474 17108 43484
rect 17164 43652 17388 43708
rect 17500 43708 17556 44380
rect 17612 44294 17668 44828
rect 17948 44772 18004 45052
rect 17612 44242 17614 44294
rect 17666 44242 17668 44294
rect 17612 44230 17668 44242
rect 17836 44716 18004 44772
rect 17836 44294 17892 44716
rect 18172 44660 18228 45388
rect 17836 44242 17838 44294
rect 17890 44242 17892 44294
rect 17836 44230 17892 44242
rect 17948 44604 18228 44660
rect 18284 45724 18396 45780
rect 17612 43764 17668 43774
rect 17500 43652 17668 43708
rect 17164 41198 17220 43652
rect 17276 43540 17332 43550
rect 17276 43446 17332 43484
rect 17500 43538 17556 43550
rect 17500 43486 17502 43538
rect 17554 43486 17556 43538
rect 16828 41134 16830 41186
rect 16882 41134 16884 41186
rect 16044 40562 16100 40572
rect 16156 40852 16212 40862
rect 15820 40350 15822 40402
rect 15874 40350 15876 40402
rect 15820 40338 15876 40350
rect 16156 40402 16212 40796
rect 16156 40350 16158 40402
rect 16210 40350 16212 40402
rect 16156 40338 16212 40350
rect 16380 40441 16436 40453
rect 16380 40389 16382 40441
rect 16434 40389 16436 40441
rect 16380 39956 16436 40389
rect 16828 40402 16884 41134
rect 16828 40350 16830 40402
rect 16882 40350 16884 40402
rect 16828 40338 16884 40350
rect 16940 41186 16996 41198
rect 16940 41134 16942 41186
rect 16994 41134 16996 41186
rect 14924 39788 15092 39844
rect 15036 39732 15092 39788
rect 15036 39666 15092 39676
rect 15372 39788 15540 39844
rect 15596 39900 16436 39956
rect 16492 40290 16548 40302
rect 16492 40238 16494 40290
rect 16546 40238 16548 40290
rect 16492 39956 16548 40238
rect 14644 39562 14700 39564
rect 14644 39510 14646 39562
rect 14698 39510 14700 39562
rect 14812 39554 14868 39564
rect 14924 39618 14980 39630
rect 14924 39566 14926 39618
rect 14978 39566 14980 39618
rect 14644 39498 14700 39510
rect 14924 39508 14980 39566
rect 14140 39398 14142 39450
rect 14194 39398 14196 39450
rect 14924 39442 14980 39452
rect 14140 39386 14196 39398
rect 13580 38770 13636 38780
rect 14644 39002 14700 39014
rect 14644 38950 14646 39002
rect 14698 38950 14700 39002
rect 14644 38836 14700 38950
rect 15372 38948 15428 39788
rect 15484 39618 15540 39630
rect 15484 39566 15486 39618
rect 15538 39566 15540 39618
rect 15484 39508 15540 39566
rect 15596 39618 15652 39900
rect 15596 39566 15598 39618
rect 15650 39566 15652 39618
rect 15596 39554 15652 39566
rect 15762 39620 15818 39630
rect 15762 39526 15818 39564
rect 16044 39508 16100 39900
rect 16492 39890 16548 39900
rect 16940 39844 16996 41134
rect 17108 41188 17220 41198
rect 17164 41132 17220 41188
rect 17276 43316 17332 43326
rect 17108 41094 17164 41132
rect 17276 40852 17332 43260
rect 17500 42532 17556 43486
rect 17500 42026 17556 42476
rect 17388 42005 17444 42017
rect 17388 41953 17390 42005
rect 17442 41953 17444 42005
rect 17388 41636 17444 41953
rect 17500 41974 17502 42026
rect 17554 41974 17556 42026
rect 17500 41860 17556 41974
rect 17612 42028 17668 43652
rect 17948 43540 18004 44604
rect 18060 44324 18116 44334
rect 18284 44324 18340 45724
rect 18396 45714 18452 45724
rect 18396 45332 18452 45342
rect 18396 45106 18452 45276
rect 18396 45054 18398 45106
rect 18450 45054 18452 45106
rect 18396 45042 18452 45054
rect 18060 44242 18062 44268
rect 18114 44242 18116 44268
rect 18228 44306 18340 44324
rect 18228 44254 18230 44306
rect 18282 44268 18340 44306
rect 18396 44324 18452 44334
rect 18282 44254 18284 44268
rect 18228 44242 18284 44254
rect 18060 44230 18116 44242
rect 18284 44100 18340 44110
rect 18172 43540 18228 43550
rect 17948 43538 18228 43540
rect 17948 43486 18174 43538
rect 18226 43486 18228 43538
rect 17948 43484 18228 43486
rect 17780 43316 17836 43326
rect 17780 43222 17836 43260
rect 17948 43092 18004 43484
rect 18172 43474 18228 43484
rect 17836 43036 18004 43092
rect 17724 42028 17780 42038
rect 17612 42026 17780 42028
rect 17612 41974 17726 42026
rect 17778 41974 17780 42026
rect 17612 41972 17780 41974
rect 17836 42028 17892 43036
rect 17948 42756 18004 42766
rect 17948 42662 18004 42700
rect 18060 42644 18116 42654
rect 17948 42028 18004 42038
rect 17836 42026 18004 42028
rect 17836 41974 17950 42026
rect 18002 41974 18004 42026
rect 17836 41972 18004 41974
rect 17724 41962 17780 41972
rect 17948 41962 18004 41972
rect 17500 41794 17556 41804
rect 17388 41570 17444 41580
rect 17500 41412 17556 41422
rect 17500 41318 17556 41356
rect 18060 40974 18116 42588
rect 18284 41972 18340 44044
rect 18396 43764 18452 44268
rect 18396 43540 18452 43708
rect 18508 43708 18564 47180
rect 19516 47170 19572 47180
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 19964 46676 20020 46686
rect 19852 46674 20020 46676
rect 19852 46622 19966 46674
rect 20018 46622 20020 46674
rect 19852 46620 20020 46622
rect 19628 46452 19684 46462
rect 18732 46450 19684 46452
rect 18732 46398 19630 46450
rect 19682 46398 19684 46450
rect 18732 46396 19684 46398
rect 18732 46002 18788 46396
rect 19628 46386 19684 46396
rect 18732 45950 18734 46002
rect 18786 45950 18788 46002
rect 18732 45938 18788 45950
rect 19852 45668 19908 46620
rect 19964 46610 20020 46620
rect 20188 46674 20244 46686
rect 20188 46622 20190 46674
rect 20242 46622 20244 46674
rect 19292 45612 19908 45668
rect 19180 44994 19236 45006
rect 19180 44942 19182 44994
rect 19234 44942 19236 44994
rect 19068 44548 19124 44558
rect 19180 44548 19236 44942
rect 19068 44546 19236 44548
rect 19068 44494 19070 44546
rect 19122 44494 19236 44546
rect 19068 44492 19236 44494
rect 19068 44482 19124 44492
rect 18676 44098 18732 44110
rect 18676 44046 18678 44098
rect 18730 44046 18732 44098
rect 18676 43876 18732 44046
rect 18676 43810 18732 43820
rect 19292 43708 19348 45612
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 20188 45332 20244 46622
rect 20188 45266 20244 45276
rect 20636 45778 20692 47628
rect 21084 47572 21140 47582
rect 20916 47236 20972 47246
rect 20636 45726 20638 45778
rect 20690 45726 20692 45778
rect 20524 44436 20580 44446
rect 19404 44324 19460 44334
rect 19684 44324 19740 44334
rect 19404 44322 19740 44324
rect 19404 44270 19406 44322
rect 19458 44270 19686 44322
rect 19738 44270 19740 44322
rect 19404 44268 19740 44270
rect 19404 44258 19460 44268
rect 19684 44258 19740 44268
rect 19964 44324 20020 44334
rect 20524 44287 20580 44380
rect 19964 44242 19966 44268
rect 20018 44242 20020 44268
rect 19964 44230 20020 44242
rect 20188 44266 20244 44278
rect 20188 44214 20190 44266
rect 20242 44214 20244 44266
rect 19628 44100 19684 44110
rect 18508 43652 18676 43708
rect 19292 43652 19572 43708
rect 18508 43540 18564 43550
rect 18396 43538 18564 43540
rect 18396 43486 18510 43538
rect 18562 43486 18564 43538
rect 18396 43484 18564 43486
rect 18508 43474 18564 43484
rect 18396 43370 18452 43382
rect 18396 43318 18398 43370
rect 18450 43318 18452 43370
rect 18396 43092 18452 43318
rect 18620 43316 18676 43652
rect 19404 43538 19460 43550
rect 19404 43486 19406 43538
rect 19458 43486 19460 43538
rect 19068 43316 19124 43326
rect 18396 43026 18452 43036
rect 18508 43260 18676 43316
rect 18732 43314 19124 43316
rect 18732 43262 19070 43314
rect 19122 43262 19124 43314
rect 18732 43260 19124 43262
rect 18284 41916 18452 41972
rect 18228 41748 18284 41758
rect 18228 41654 18284 41692
rect 18060 40964 18172 40974
rect 18060 40908 18116 40964
rect 18116 40870 18172 40908
rect 17276 40786 17332 40796
rect 17724 40404 17780 40414
rect 17724 40310 17780 40348
rect 17276 39844 17332 39854
rect 16940 39842 17332 39844
rect 16940 39790 17278 39842
rect 17330 39790 17332 39842
rect 16940 39788 17332 39790
rect 17276 39778 17332 39788
rect 16156 39732 16212 39742
rect 16716 39732 16772 39742
rect 16156 39730 16660 39732
rect 16156 39678 16158 39730
rect 16210 39678 16660 39730
rect 16156 39676 16660 39678
rect 16156 39666 16212 39676
rect 16604 39618 16660 39676
rect 16604 39566 16606 39618
rect 16658 39566 16660 39618
rect 16604 39554 16660 39566
rect 16716 39618 16772 39676
rect 16716 39566 16718 39618
rect 16770 39566 16772 39618
rect 18172 39618 18228 39630
rect 16716 39554 16772 39566
rect 16882 39564 16938 39574
rect 16828 39562 16938 39564
rect 16828 39510 16884 39562
rect 16936 39510 16938 39562
rect 16044 39452 16492 39508
rect 15484 39060 15540 39452
rect 15708 39396 15764 39406
rect 15484 39004 15652 39060
rect 15372 38882 15428 38892
rect 15260 38862 15316 38874
rect 14644 38770 14700 38780
rect 14812 38834 14868 38846
rect 14812 38782 14814 38834
rect 14866 38782 14868 38834
rect 14812 38388 14868 38782
rect 14812 38322 14868 38332
rect 15260 38810 15262 38862
rect 15314 38810 15316 38862
rect 15260 38164 15316 38810
rect 15484 38836 15540 38846
rect 15484 38742 15540 38780
rect 15596 38724 15652 39004
rect 15708 38946 15764 39340
rect 15708 38894 15710 38946
rect 15762 38894 15764 38946
rect 15708 38882 15764 38894
rect 15876 38948 15932 38958
rect 15876 38890 15932 38892
rect 15876 38838 15878 38890
rect 15930 38838 15932 38890
rect 16436 38946 16492 39452
rect 16436 38894 16438 38946
rect 16490 38894 16492 38946
rect 16436 38882 16492 38894
rect 16828 39498 16938 39510
rect 18172 39566 18174 39618
rect 18226 39566 18228 39618
rect 16828 38948 16884 39498
rect 18172 39060 18228 39566
rect 18172 38994 18228 39004
rect 16828 38882 16884 38892
rect 15876 38826 15932 38838
rect 16716 38834 16772 38846
rect 16716 38782 16718 38834
rect 16770 38782 16772 38834
rect 15596 38658 15652 38668
rect 16548 38724 16604 38734
rect 15260 38098 15316 38108
rect 15820 38388 15876 38398
rect 14140 38052 14196 38062
rect 13356 37998 13358 38050
rect 13410 37998 13412 38050
rect 13356 37986 13412 37998
rect 13580 38050 14196 38052
rect 13580 37998 14142 38050
rect 14194 37998 14196 38050
rect 13580 37996 14196 37998
rect 12852 37940 12908 37950
rect 12852 37938 13300 37940
rect 12852 37886 12854 37938
rect 12906 37886 13300 37938
rect 12852 37884 13300 37886
rect 12852 37874 12908 37884
rect 12908 37492 12964 37502
rect 12908 37378 12964 37436
rect 12908 37326 12910 37378
rect 12962 37326 12964 37378
rect 12908 37314 12964 37326
rect 13244 37266 13300 37884
rect 13580 37490 13636 37996
rect 14140 37986 14196 37996
rect 13580 37438 13582 37490
rect 13634 37438 13636 37490
rect 13580 37426 13636 37438
rect 15820 37490 15876 38332
rect 16548 38274 16604 38668
rect 16548 38222 16550 38274
rect 16602 38222 16604 38274
rect 16548 38210 16604 38222
rect 15820 37438 15822 37490
rect 15874 37438 15876 37490
rect 13244 37214 13246 37266
rect 13298 37214 13300 37266
rect 13244 37202 13300 37214
rect 15820 37268 15876 37438
rect 15820 37202 15876 37212
rect 15932 38164 15988 38174
rect 14924 36708 14980 36718
rect 14252 36706 14980 36708
rect 14252 36654 14926 36706
rect 14978 36654 14980 36706
rect 14252 36652 14980 36654
rect 12964 36466 13412 36484
rect 12460 35702 12462 35754
rect 12514 35702 12516 35754
rect 12460 35690 12516 35702
rect 12572 35868 12740 35924
rect 12796 36426 12852 36438
rect 12796 36374 12798 36426
rect 12850 36374 12852 36426
rect 12964 36414 12966 36466
rect 13018 36428 13412 36466
rect 13018 36414 13020 36428
rect 12964 36402 13020 36414
rect 12796 35924 12852 36374
rect 13356 35924 13412 36428
rect 13636 36258 13692 36270
rect 13636 36206 13638 36258
rect 13690 36206 13692 36258
rect 13636 35924 13692 36206
rect 12796 35868 12964 35924
rect 12236 34738 12292 34748
rect 12236 34356 12292 34366
rect 12236 34262 12292 34300
rect 11900 34130 12068 34132
rect 11900 34078 11902 34130
rect 11954 34078 12068 34130
rect 11900 34076 12068 34078
rect 11900 34066 11956 34076
rect 11900 33346 11956 33358
rect 11900 33294 11902 33346
rect 11954 33294 11956 33346
rect 11900 33236 11956 33294
rect 11900 33170 11956 33180
rect 12460 33346 12516 33358
rect 12460 33294 12462 33346
rect 12514 33294 12516 33346
rect 12460 33236 12516 33294
rect 12460 33170 12516 33180
rect 12572 33124 12628 35868
rect 12684 35754 12740 35766
rect 12684 35702 12686 35754
rect 12738 35702 12740 35754
rect 12684 35364 12740 35702
rect 12684 35298 12740 35308
rect 12796 35733 12852 35745
rect 12796 35681 12798 35733
rect 12850 35681 12852 35733
rect 12796 35028 12852 35681
rect 12908 35364 12964 35868
rect 12908 35298 12964 35308
rect 13356 35868 13692 35924
rect 12684 34972 12852 35028
rect 12684 34692 12740 34972
rect 12796 34804 12852 34814
rect 12796 34710 12852 34748
rect 12684 34626 12740 34636
rect 12908 34692 12964 34702
rect 12908 34366 12964 34636
rect 12852 34356 12964 34366
rect 12684 34354 12964 34356
rect 12684 34302 12854 34354
rect 12906 34302 12964 34354
rect 12684 34300 12964 34302
rect 13356 34468 13412 35868
rect 12684 33460 12740 34300
rect 12852 34290 12908 34300
rect 13020 34132 13076 34142
rect 12684 33394 12740 33404
rect 12908 33796 12964 33806
rect 12908 33458 12964 33740
rect 12908 33406 12910 33458
rect 12962 33406 12964 33458
rect 12908 33394 12964 33406
rect 12796 33348 12852 33358
rect 12796 33279 12798 33292
rect 12850 33279 12852 33292
rect 12796 33254 12852 33279
rect 12572 33068 12964 33124
rect 10780 32510 10782 32562
rect 10834 32510 10836 32562
rect 10780 32498 10836 32510
rect 10668 32162 10724 32172
rect 10332 32116 10388 32126
rect 10332 31230 10388 32060
rect 11004 32002 11060 32732
rect 11676 32722 11732 32732
rect 11004 31950 11006 32002
rect 11058 31950 11060 32002
rect 11004 31938 11060 31950
rect 12684 32450 12740 32462
rect 12684 32398 12686 32450
rect 12738 32398 12740 32450
rect 12684 31948 12740 32398
rect 12348 31892 12740 31948
rect 10612 31780 10668 31790
rect 10612 31556 10668 31724
rect 11247 31780 11303 31790
rect 11247 31686 11303 31724
rect 12124 31778 12180 31790
rect 12124 31726 12126 31778
rect 12178 31726 12180 31778
rect 12124 31556 12180 31726
rect 10612 31554 10948 31556
rect 10612 31502 10614 31554
rect 10666 31502 10948 31554
rect 10612 31500 10948 31502
rect 10612 31490 10668 31500
rect 10332 31218 10444 31230
rect 10332 31166 10390 31218
rect 10442 31166 10444 31218
rect 10332 31164 10444 31166
rect 10388 31154 10444 31164
rect 10668 30324 10724 30334
rect 10668 30100 10724 30268
rect 10668 30044 10743 30100
rect 10444 29540 10500 29550
rect 10444 29446 10500 29484
rect 10687 29482 10743 30044
rect 10687 29430 10689 29482
rect 10741 29430 10743 29482
rect 10687 29418 10743 29430
rect 10220 29036 10836 29092
rect 9996 28690 10052 28700
rect 10220 28868 10276 28878
rect 10220 28644 10276 28812
rect 9660 28532 9716 28542
rect 9660 28530 9940 28532
rect 9660 28478 9662 28530
rect 9714 28478 9940 28530
rect 9660 28476 9940 28478
rect 9660 28466 9716 28476
rect 9884 27972 9940 28476
rect 9492 27916 9828 27972
rect 9492 27914 9548 27916
rect 9492 27862 9494 27914
rect 9546 27862 9548 27914
rect 9492 27850 9548 27862
rect 9324 27794 9380 27804
rect 7868 26852 8260 26908
rect 6972 26628 7028 26638
rect 6972 26334 7028 26572
rect 6972 26282 6974 26334
rect 7026 26282 7028 26334
rect 6972 26270 7028 26282
rect 7196 26290 7252 26302
rect 7196 26238 7198 26290
rect 7250 26238 7252 26290
rect 6860 26180 6916 26190
rect 6860 26086 6916 26124
rect 6636 25330 6692 25340
rect 7196 25284 7252 26238
rect 8204 26178 8260 26852
rect 8316 26852 8372 26862
rect 8316 26334 8372 26796
rect 8316 26282 8318 26334
rect 8370 26282 8372 26334
rect 8316 26270 8372 26282
rect 8652 26852 9268 26908
rect 9660 27746 9716 27758
rect 9660 27694 9662 27746
rect 9714 27694 9716 27746
rect 9660 26964 9716 27694
rect 9772 27188 9828 27916
rect 9884 27858 9940 27916
rect 9884 27806 9886 27858
rect 9938 27806 9940 27858
rect 10220 27914 10276 28588
rect 10220 27862 10222 27914
rect 10274 27862 10276 27914
rect 10220 27850 10276 27862
rect 9884 27636 9940 27806
rect 9884 27580 10164 27636
rect 10108 27188 10164 27580
rect 9772 27186 10052 27188
rect 9772 27134 9774 27186
rect 9826 27134 10052 27186
rect 9772 27132 10052 27134
rect 9772 27122 9828 27132
rect 9660 26898 9716 26908
rect 9996 26908 10052 27132
rect 10276 27242 10332 27254
rect 10276 27190 10278 27242
rect 10330 27190 10332 27242
rect 10276 27188 10332 27190
rect 10276 27132 10724 27188
rect 10108 27074 10164 27132
rect 10108 27022 10110 27074
rect 10162 27022 10164 27074
rect 10108 27010 10164 27022
rect 10668 27074 10724 27132
rect 10668 27022 10670 27074
rect 10722 27022 10724 27074
rect 10668 27010 10724 27022
rect 9996 26852 10164 26908
rect 8652 26290 8708 26852
rect 8652 26238 8654 26290
rect 8706 26238 8708 26290
rect 8652 26226 8708 26238
rect 9996 26292 10052 26302
rect 9996 26198 10052 26236
rect 10108 26290 10164 26852
rect 10276 26852 10332 26862
rect 10276 26514 10332 26796
rect 10276 26462 10278 26514
rect 10330 26462 10332 26514
rect 10276 26450 10332 26462
rect 10444 26516 10500 26526
rect 10108 26238 10110 26290
rect 10162 26238 10164 26290
rect 10108 26226 10164 26238
rect 8204 26126 8206 26178
rect 8258 26126 8260 26178
rect 8204 26114 8260 26126
rect 9660 26068 9716 26078
rect 9100 26066 9716 26068
rect 9100 26014 9662 26066
rect 9714 26014 9716 26066
rect 9100 26012 9716 26014
rect 9100 25618 9156 26012
rect 9660 26002 9716 26012
rect 9100 25566 9102 25618
rect 9154 25566 9156 25618
rect 9100 25554 9156 25566
rect 7196 25218 7252 25228
rect 7980 25508 8036 25518
rect 6524 24994 6580 25004
rect 6300 24882 6356 24892
rect 7308 24948 7364 24958
rect 7308 24722 7364 24892
rect 7308 24670 7310 24722
rect 7362 24670 7364 24722
rect 7308 24658 7364 24670
rect 7980 24724 8036 25452
rect 8316 25508 8372 25518
rect 8316 25414 8372 25452
rect 10444 24778 10500 26460
rect 10780 25508 10836 29036
rect 10892 28980 10948 31500
rect 11676 31444 11732 31454
rect 11004 30994 11060 31006
rect 11004 30942 11006 30994
rect 11058 30942 11060 30994
rect 11004 30212 11060 30942
rect 11340 30770 11396 30782
rect 11340 30718 11342 30770
rect 11394 30718 11396 30770
rect 11340 30212 11396 30718
rect 11676 30324 11732 31388
rect 11900 31220 11956 31230
rect 12124 31220 12180 31500
rect 11900 31218 12180 31220
rect 11900 31166 11902 31218
rect 11954 31166 12180 31218
rect 11900 31164 12180 31166
rect 12348 31444 12404 31892
rect 12796 31780 12852 31790
rect 12796 31686 12852 31724
rect 12516 31668 12572 31678
rect 12516 31574 12572 31612
rect 11900 31154 11956 31164
rect 12236 30996 12292 31006
rect 12348 30996 12404 31388
rect 12516 31108 12572 31118
rect 12740 31052 12796 31062
rect 12516 31014 12572 31052
rect 12684 31050 12796 31052
rect 12236 30994 12404 30996
rect 12236 30942 12238 30994
rect 12290 30942 12404 30994
rect 12236 30940 12404 30942
rect 12684 30998 12742 31050
rect 12794 30998 12796 31050
rect 12684 30986 12796 30998
rect 12236 30930 12292 30940
rect 12684 30884 12740 30986
rect 12404 30436 12460 30446
rect 12684 30436 12740 30828
rect 12404 30434 12740 30436
rect 12404 30382 12406 30434
rect 12458 30382 12740 30434
rect 12404 30380 12740 30382
rect 12404 30370 12460 30380
rect 11452 30212 11508 30222
rect 11340 30210 11508 30212
rect 11340 30158 11454 30210
rect 11506 30158 11508 30210
rect 11340 30156 11508 30158
rect 11004 30118 11060 30156
rect 11452 29988 11508 30156
rect 11676 30210 11732 30268
rect 11676 30158 11678 30210
rect 11730 30158 11732 30210
rect 11676 30146 11732 30158
rect 12236 30212 12292 30222
rect 12236 30118 12292 30156
rect 11956 30100 12012 30110
rect 11452 29428 11508 29932
rect 11788 30098 12012 30100
rect 11788 30046 11958 30098
rect 12010 30046 12012 30098
rect 11788 30044 12012 30046
rect 11564 29428 11620 29438
rect 11452 29426 11620 29428
rect 11452 29374 11566 29426
rect 11618 29374 11620 29426
rect 11452 29372 11620 29374
rect 11564 29362 11620 29372
rect 11564 29092 11620 29102
rect 11788 29092 11844 30044
rect 11956 30034 12012 30044
rect 12796 29876 12852 29886
rect 12684 29594 12740 29606
rect 12684 29542 12686 29594
rect 12738 29542 12740 29594
rect 12348 29465 12404 29477
rect 10892 28924 11284 28980
rect 11228 27188 11284 28924
rect 11396 28868 11452 28878
rect 11396 28774 11452 28812
rect 11340 27746 11396 27758
rect 11340 27694 11342 27746
rect 11394 27694 11396 27746
rect 11340 27412 11396 27694
rect 11340 27346 11396 27356
rect 11228 27132 11396 27188
rect 10892 27076 10948 27086
rect 10892 26290 10948 27020
rect 11116 27074 11172 27086
rect 11116 27022 11118 27074
rect 11170 27022 11172 27074
rect 11116 26628 11172 27022
rect 10892 26238 10894 26290
rect 10946 26238 10948 26290
rect 10892 26226 10948 26238
rect 11004 26572 11116 26628
rect 11004 25618 11060 26572
rect 11116 26562 11172 26572
rect 11228 26516 11284 26526
rect 11228 26404 11284 26460
rect 11116 26348 11284 26404
rect 11116 26334 11172 26348
rect 11116 26282 11118 26334
rect 11170 26282 11172 26334
rect 11116 26270 11172 26282
rect 11228 26180 11284 26190
rect 11228 26086 11284 26124
rect 11004 25566 11006 25618
rect 11058 25566 11060 25618
rect 11004 25554 11060 25566
rect 10780 25452 10948 25508
rect 10892 25284 10948 25452
rect 10892 25228 11172 25284
rect 8092 24724 8148 24734
rect 7980 24722 8148 24724
rect 7980 24670 8094 24722
rect 8146 24670 8148 24722
rect 7980 24668 8148 24670
rect 6300 23940 6356 23950
rect 6188 23938 6356 23940
rect 6188 23886 6302 23938
rect 6354 23886 6356 23938
rect 6188 23884 6356 23886
rect 6300 23874 6356 23884
rect 6636 23938 6692 23950
rect 6636 23886 6638 23938
rect 6690 23886 6692 23938
rect 6076 23835 6132 23847
rect 6636 23268 6692 23886
rect 6636 23202 6692 23212
rect 7868 23940 7924 23950
rect 7980 23940 8036 24668
rect 8092 24658 8148 24668
rect 9100 24724 9156 24734
rect 9100 24630 9156 24668
rect 10164 24724 10220 24734
rect 10164 24630 10220 24668
rect 10444 24726 10446 24778
rect 10498 24726 10500 24778
rect 8764 24498 8820 24510
rect 8764 24446 8766 24498
rect 8818 24446 8820 24498
rect 8652 24052 8708 24062
rect 8764 24052 8820 24446
rect 8652 24050 8820 24052
rect 8652 23998 8654 24050
rect 8706 23998 8820 24050
rect 8652 23996 8820 23998
rect 10444 24052 10500 24726
rect 10668 25172 10724 25182
rect 10668 24778 10724 25116
rect 10668 24726 10670 24778
rect 10722 24726 10724 24778
rect 10668 24714 10724 24726
rect 10892 25060 10948 25070
rect 10892 24778 10948 25004
rect 10892 24726 10894 24778
rect 10946 24726 10948 24778
rect 10892 24714 10948 24726
rect 11004 24836 11060 24846
rect 11004 24778 11060 24780
rect 11004 24726 11006 24778
rect 11058 24726 11060 24778
rect 11004 24714 11060 24726
rect 10556 24052 10612 24062
rect 10444 24050 10612 24052
rect 10444 23998 10558 24050
rect 10610 23998 10612 24050
rect 10444 23996 10612 23998
rect 8652 23986 8708 23996
rect 10556 23986 10612 23996
rect 7868 23938 8036 23940
rect 7868 23886 7870 23938
rect 7922 23886 8036 23938
rect 7868 23884 8036 23886
rect 7868 23378 7924 23884
rect 11116 23828 11172 25228
rect 11116 23762 11172 23772
rect 11228 24722 11284 24734
rect 11228 24670 11230 24722
rect 11282 24670 11284 24722
rect 7868 23326 7870 23378
rect 7922 23326 7924 23378
rect 6860 23181 6916 23193
rect 6076 23169 6132 23181
rect 6076 23117 6078 23169
rect 6130 23117 6132 23169
rect 6076 21700 6132 23117
rect 6860 23156 6862 23181
rect 6914 23156 6916 23181
rect 6188 23044 6244 23054
rect 6188 23042 6692 23044
rect 6188 22990 6190 23042
rect 6242 22990 6692 23042
rect 6188 22988 6692 22990
rect 6188 22978 6244 22988
rect 6636 22482 6692 22988
rect 6636 22430 6638 22482
rect 6690 22430 6692 22482
rect 6636 22418 6692 22430
rect 6412 21700 6468 21710
rect 6076 21698 6468 21700
rect 6076 21646 6414 21698
rect 6466 21646 6468 21698
rect 6076 21644 6468 21646
rect 6412 21634 6468 21644
rect 6655 21586 6711 21598
rect 6655 21534 6657 21586
rect 6709 21534 6711 21586
rect 6655 21476 6711 21534
rect 5964 21420 6711 21476
rect 5796 21364 5852 21374
rect 5628 21074 5684 21084
rect 5740 21362 5852 21364
rect 5740 21310 5798 21362
rect 5850 21310 5852 21362
rect 5740 21298 5852 21310
rect 5180 20750 5182 20802
rect 5234 20750 5236 20802
rect 5180 20692 5236 20750
rect 5180 20636 5572 20692
rect 4956 20626 5012 20636
rect 5292 20186 5348 20198
rect 4956 20132 5012 20142
rect 3612 19954 3668 19964
rect 3724 19964 4116 20020
rect 4732 20020 4788 20030
rect 4788 19964 4900 20020
rect 3500 18398 3502 18450
rect 3554 18398 3556 18450
rect 3724 18494 3780 19964
rect 4732 19926 4788 19964
rect 4284 19906 4340 19918
rect 4284 19854 4286 19906
rect 4338 19854 4340 19906
rect 4060 19346 4116 19358
rect 4060 19294 4062 19346
rect 4114 19294 4116 19346
rect 3724 18442 3726 18494
rect 3778 18442 3780 18494
rect 3724 18430 3780 18442
rect 3836 18900 3892 18910
rect 3500 18340 3556 18398
rect 3500 18274 3556 18284
rect 3836 18338 3892 18844
rect 4060 18452 4116 19294
rect 4284 19236 4340 19854
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4732 19348 4788 19358
rect 4284 19180 4564 19236
rect 4284 18618 4340 18630
rect 4284 18566 4286 18618
rect 4338 18566 4340 18618
rect 4284 18564 4340 18566
rect 4284 18498 4340 18508
rect 4060 18386 4116 18396
rect 4396 18450 4452 18462
rect 4396 18398 4398 18450
rect 4450 18398 4452 18450
rect 3836 18286 3838 18338
rect 3890 18286 3892 18338
rect 3836 18274 3892 18286
rect 2716 18228 2772 18238
rect 4396 18228 4452 18398
rect 4508 18340 4564 19180
rect 4732 18506 4788 19292
rect 4732 18454 4734 18506
rect 4786 18454 4788 18506
rect 4732 18442 4788 18454
rect 4508 18274 4564 18284
rect 2380 18226 2772 18228
rect 2380 18174 2718 18226
rect 2770 18174 2772 18226
rect 2380 18172 2772 18174
rect 2380 17778 2436 18172
rect 2716 18162 2772 18172
rect 4060 18172 4396 18228
rect 2380 17726 2382 17778
rect 2434 17726 2436 17778
rect 2380 17714 2436 17726
rect 1596 17614 1598 17666
rect 1650 17614 1652 17666
rect 1596 16882 1652 17614
rect 1596 16830 1598 16882
rect 1650 16830 1652 16882
rect 1596 16818 1652 16830
rect 3948 17108 4004 17118
rect 2380 16770 2436 16782
rect 2380 16718 2382 16770
rect 2434 16718 2436 16770
rect 2380 16324 2436 16718
rect 2492 16324 2548 16334
rect 2380 16322 2548 16324
rect 2380 16270 2494 16322
rect 2546 16270 2548 16322
rect 2380 16268 2548 16270
rect 2492 16258 2548 16268
rect 3388 16324 3444 16334
rect 2828 16100 2884 16110
rect 2828 16006 2884 16044
rect 3164 16098 3220 16110
rect 3164 16046 3166 16098
rect 3218 16046 3220 16098
rect 3164 15988 3220 16046
rect 3388 16083 3444 16268
rect 3388 16031 3390 16083
rect 3442 16031 3444 16083
rect 3388 16019 3444 16031
rect 3500 16210 3556 16222
rect 3500 16158 3502 16210
rect 3554 16158 3556 16210
rect 3164 15922 3220 15932
rect 3500 15764 3556 16158
rect 3948 16098 4004 17052
rect 3948 16046 3950 16098
rect 4002 16046 4004 16098
rect 3948 16034 4004 16046
rect 4060 16100 4116 18172
rect 4396 18162 4452 18172
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4844 18004 4900 19964
rect 4956 19206 5012 20076
rect 5292 20134 5294 20186
rect 5346 20134 5348 20186
rect 4956 19154 4958 19206
rect 5010 19154 5012 19206
rect 4956 19142 5012 19154
rect 5068 20045 5124 20057
rect 5068 19993 5070 20045
rect 5122 19993 5124 20045
rect 5068 18900 5124 19993
rect 5292 19460 5348 20134
rect 5404 20020 5460 20030
rect 5404 19926 5460 19964
rect 5516 19796 5572 20636
rect 5740 20020 5796 21298
rect 6468 21028 6524 21038
rect 6655 21028 6711 21420
rect 6655 20972 6804 21028
rect 6468 20858 6524 20972
rect 6188 20804 6244 20814
rect 6020 20802 6244 20804
rect 6020 20750 6190 20802
rect 6242 20750 6244 20802
rect 6468 20806 6470 20858
rect 6522 20806 6524 20858
rect 6468 20794 6524 20806
rect 6636 20802 6692 20814
rect 6020 20748 6244 20750
rect 5908 20690 5964 20702
rect 5908 20638 5910 20690
rect 5962 20638 5964 20690
rect 5908 20244 5964 20638
rect 5908 20178 5964 20188
rect 5740 19954 5796 19964
rect 5852 20018 5908 20030
rect 5852 19966 5854 20018
rect 5906 19966 5908 20018
rect 5852 19796 5908 19966
rect 5516 19740 5908 19796
rect 6020 19850 6076 20748
rect 6188 20738 6244 20748
rect 6636 20750 6638 20802
rect 6690 20750 6692 20802
rect 6300 20690 6356 20702
rect 6300 20638 6302 20690
rect 6354 20638 6356 20690
rect 6020 19798 6022 19850
rect 6074 19798 6076 19850
rect 6020 19786 6076 19798
rect 6188 20244 6244 20254
rect 6188 19460 6244 20188
rect 5292 19394 5348 19404
rect 6076 19404 6244 19460
rect 5628 19348 5684 19358
rect 5628 19254 5684 19292
rect 5964 19236 6020 19246
rect 5852 19234 6020 19236
rect 5068 18834 5124 18844
rect 5740 19190 5796 19202
rect 5740 19138 5742 19190
rect 5794 19138 5796 19190
rect 4844 17890 4900 17948
rect 4844 17838 4846 17890
rect 4898 17838 4900 17890
rect 4844 17826 4900 17838
rect 4956 18450 5012 18462
rect 4956 18398 4958 18450
rect 5010 18398 5012 18450
rect 4284 17668 4340 17678
rect 4284 17574 4340 17612
rect 4284 17108 4340 17118
rect 4284 16994 4340 17052
rect 4284 16942 4286 16994
rect 4338 16942 4340 16994
rect 4284 16930 4340 16942
rect 4172 16884 4228 16894
rect 4172 16212 4228 16828
rect 4844 16884 4900 16894
rect 4956 16884 5012 18398
rect 5740 18450 5796 19138
rect 5740 18398 5742 18450
rect 5794 18398 5796 18450
rect 5460 18228 5516 18238
rect 5460 18134 5516 18172
rect 5740 18228 5796 18398
rect 5740 18162 5796 18172
rect 5852 19182 5966 19234
rect 6018 19182 6020 19234
rect 5852 19180 6020 19182
rect 5852 18450 5908 19180
rect 5964 19170 6020 19180
rect 6076 18676 6132 19404
rect 6300 19348 6356 20638
rect 6636 20356 6692 20750
rect 6636 20290 6692 20300
rect 6748 20188 6804 20972
rect 5852 18398 5854 18450
rect 5906 18398 5908 18450
rect 5180 17892 5236 17902
rect 5180 17666 5236 17836
rect 5180 17614 5182 17666
rect 5234 17614 5236 17666
rect 5180 17602 5236 17614
rect 5516 17892 5572 17902
rect 5404 17556 5460 17566
rect 5180 17444 5236 17454
rect 4844 16882 5012 16884
rect 4844 16830 4846 16882
rect 4898 16830 5012 16882
rect 4844 16828 5012 16830
rect 5068 16909 5124 16922
rect 5068 16884 5070 16909
rect 5122 16884 5124 16909
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4732 16324 4788 16334
rect 4284 16212 4340 16222
rect 4172 16210 4340 16212
rect 4172 16158 4286 16210
rect 4338 16158 4340 16210
rect 4172 16156 4340 16158
rect 4284 16146 4340 16156
rect 4060 16068 4172 16100
rect 4060 16044 4118 16068
rect 4116 16016 4118 16044
rect 4170 16016 4172 16068
rect 4116 16004 4172 16016
rect 4620 16098 4676 16110
rect 4620 16046 4622 16098
rect 4674 16046 4676 16098
rect 3500 15698 3556 15708
rect 4284 15988 4340 15998
rect 2828 15316 2884 15326
rect 2828 15222 2884 15260
rect 2492 15092 2548 15102
rect 2380 15090 2548 15092
rect 2380 15038 2494 15090
rect 2546 15038 2548 15090
rect 2380 15036 2548 15038
rect 2380 14642 2436 15036
rect 2492 15026 2548 15036
rect 2380 14590 2382 14642
rect 2434 14590 2436 14642
rect 2380 14578 2436 14590
rect 4284 14642 4340 15932
rect 4620 15988 4676 16046
rect 4732 16098 4788 16268
rect 4732 16046 4734 16098
rect 4786 16046 4788 16098
rect 4732 16034 4788 16046
rect 4620 15922 4676 15932
rect 4620 15764 4676 15774
rect 4844 15764 4900 16828
rect 5068 16818 5124 16828
rect 5180 16436 5236 17388
rect 5012 16380 5236 16436
rect 5012 16322 5068 16380
rect 5012 16270 5014 16322
rect 5066 16270 5068 16322
rect 5012 16258 5068 16270
rect 4676 15708 4788 15764
rect 4844 15708 5012 15764
rect 4620 15698 4676 15708
rect 4620 15482 4676 15494
rect 4620 15430 4622 15482
rect 4674 15430 4676 15482
rect 4508 15314 4564 15326
rect 4508 15262 4510 15314
rect 4562 15262 4564 15314
rect 4508 15092 4564 15262
rect 4620 15316 4676 15430
rect 4732 15428 4788 15708
rect 4732 15372 4844 15428
rect 4788 15370 4844 15372
rect 4788 15318 4790 15370
rect 4842 15318 4844 15370
rect 4788 15306 4844 15318
rect 4620 15250 4676 15260
rect 4956 15148 5012 15708
rect 5180 15314 5236 16380
rect 5292 17050 5348 17062
rect 5292 16998 5294 17050
rect 5346 16998 5348 17050
rect 5292 16100 5348 16998
rect 5404 16882 5460 17500
rect 5404 16830 5406 16882
rect 5458 16830 5460 16882
rect 5404 16324 5460 16830
rect 5404 16258 5460 16268
rect 5292 16034 5348 16044
rect 5180 15262 5182 15314
rect 5234 15262 5236 15314
rect 5180 15250 5236 15262
rect 4956 15092 5124 15148
rect 4508 15036 5124 15092
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4284 14590 4286 14642
rect 4338 14590 4340 14642
rect 4284 14578 4340 14590
rect 1596 14530 1652 14542
rect 1596 14478 1598 14530
rect 1650 14478 1652 14530
rect 1596 12292 1652 14478
rect 4844 14306 4900 15036
rect 5180 14530 5236 14542
rect 5180 14478 5182 14530
rect 5234 14478 5236 14530
rect 5180 14420 5236 14478
rect 5180 14354 5236 14364
rect 5516 14420 5572 17836
rect 5852 17780 5908 18398
rect 5740 17724 5908 17780
rect 5964 18620 6132 18676
rect 6244 19292 6356 19348
rect 6412 20132 6468 20142
rect 5964 17780 6020 18620
rect 6076 18450 6132 18462
rect 6076 18398 6078 18450
rect 6130 18398 6132 18450
rect 6076 18340 6132 18398
rect 6076 18274 6132 18284
rect 6244 18282 6300 19292
rect 6244 18230 6246 18282
rect 6298 18230 6300 18282
rect 6244 18218 6300 18230
rect 5740 17668 5796 17724
rect 5964 17714 6020 17724
rect 6300 18116 6356 18126
rect 5740 16098 5796 17612
rect 6188 17666 6244 17678
rect 6188 17614 6190 17666
rect 6242 17614 6244 17666
rect 5908 17556 5964 17566
rect 6188 17556 6244 17614
rect 6300 17666 6356 18060
rect 6300 17614 6302 17666
rect 6354 17614 6356 17666
rect 6300 17602 6356 17614
rect 5908 17462 5964 17500
rect 6020 17500 6244 17556
rect 6020 17332 6076 17500
rect 6412 17444 6468 20076
rect 6636 20132 6804 20188
rect 6860 20244 6916 23100
rect 7868 22372 7924 23326
rect 9660 23380 9716 23390
rect 9660 23286 9716 23324
rect 9996 23154 10052 23166
rect 9996 23102 9998 23154
rect 10050 23102 10052 23154
rect 9996 23044 10052 23102
rect 10836 23156 10892 23166
rect 10836 23062 10892 23100
rect 10388 23044 10444 23054
rect 9996 23042 10444 23044
rect 9996 22990 10390 23042
rect 10442 22990 10444 23042
rect 9996 22988 10444 22990
rect 9996 22708 10052 22988
rect 10388 22978 10444 22988
rect 9548 22652 10052 22708
rect 10892 22932 10948 22942
rect 7868 22306 7924 22316
rect 8876 22372 8932 22382
rect 8876 22278 8932 22316
rect 8540 22258 8596 22270
rect 8540 22206 8542 22258
rect 8594 22206 8596 22258
rect 7532 21588 7588 21598
rect 7532 21586 7812 21588
rect 7532 21534 7534 21586
rect 7586 21534 7812 21586
rect 7532 21532 7812 21534
rect 7532 21522 7588 21532
rect 7084 21140 7140 21150
rect 6860 20178 6916 20188
rect 6972 21028 7028 21038
rect 6636 20018 6692 20132
rect 6636 19966 6638 20018
rect 6690 19966 6692 20018
rect 6972 20074 7028 20972
rect 7084 21026 7140 21084
rect 7756 21038 7812 21532
rect 7084 20974 7086 21026
rect 7138 20974 7140 21026
rect 7084 20962 7140 20974
rect 7700 21028 7812 21038
rect 7756 20972 7812 21028
rect 7700 20934 7756 20972
rect 7420 20804 7476 20814
rect 6972 20022 6974 20074
rect 7026 20022 7028 20074
rect 6972 20010 7028 20022
rect 7084 20802 7476 20804
rect 7084 20750 7422 20802
rect 7474 20750 7476 20802
rect 7084 20748 7476 20750
rect 6636 19954 6692 19966
rect 6636 19234 6692 19246
rect 6636 19182 6638 19234
rect 6690 19182 6692 19234
rect 6636 18788 6692 19182
rect 6524 18732 6692 18788
rect 6524 18452 6580 18732
rect 7084 18676 7140 20748
rect 7420 20738 7476 20748
rect 7868 20804 7924 20814
rect 7868 20710 7924 20748
rect 8092 20804 8148 20814
rect 7308 20244 7364 20254
rect 6972 18620 7140 18676
rect 7196 20186 7252 20198
rect 7196 20134 7198 20186
rect 7250 20134 7252 20186
rect 6524 18386 6580 18396
rect 6636 18450 6692 18462
rect 6636 18398 6638 18450
rect 6690 18398 6692 18450
rect 6636 18004 6692 18398
rect 6636 17938 6692 17948
rect 6972 17892 7028 18620
rect 7084 18489 7140 18501
rect 7084 18437 7086 18489
rect 7138 18437 7140 18489
rect 7084 18228 7140 18437
rect 7084 18162 7140 18172
rect 6972 17826 7028 17836
rect 5964 17276 6076 17332
rect 6132 17388 6468 17444
rect 6524 17780 6580 17790
rect 5740 16046 5742 16098
rect 5794 16046 5796 16098
rect 5740 15316 5796 16046
rect 5852 17108 5908 17118
rect 5852 16098 5908 17052
rect 5964 16996 6020 17276
rect 5964 16324 6020 16940
rect 6132 17106 6188 17388
rect 6132 17054 6134 17106
rect 6186 17054 6188 17106
rect 6132 16884 6188 17054
rect 6412 16884 6468 16894
rect 6132 16818 6188 16828
rect 6300 16882 6468 16884
rect 6300 16830 6414 16882
rect 6466 16830 6468 16882
rect 6300 16828 6468 16830
rect 6132 16324 6188 16334
rect 5964 16322 6188 16324
rect 5964 16270 6134 16322
rect 6186 16270 6188 16322
rect 5964 16268 6188 16270
rect 6132 16258 6188 16268
rect 5852 16046 5854 16098
rect 5906 16046 5908 16098
rect 5852 16034 5908 16046
rect 6300 15988 6356 16828
rect 6412 16818 6468 16828
rect 6524 16548 6580 17724
rect 7084 17778 7140 17790
rect 7084 17726 7086 17778
rect 7138 17726 7140 17778
rect 6636 17666 6692 17678
rect 6636 17614 6638 17666
rect 6690 17614 6692 17666
rect 6636 17108 6692 17614
rect 6972 17622 7028 17634
rect 6972 17570 6974 17622
rect 7026 17570 7028 17622
rect 6972 17332 7028 17570
rect 6636 17042 6692 17052
rect 6860 17276 6972 17332
rect 6860 16938 6916 17276
rect 6972 17266 7028 17276
rect 7084 17108 7140 17726
rect 6860 16886 6862 16938
rect 6914 16886 6916 16938
rect 6860 16874 6916 16886
rect 6972 17052 7140 17108
rect 7196 17668 7252 20134
rect 7308 20018 7364 20188
rect 7308 19966 7310 20018
rect 7362 19966 7364 20018
rect 7308 19954 7364 19966
rect 7756 20056 7812 20068
rect 7756 20020 7758 20056
rect 7810 20020 7812 20056
rect 7756 19954 7812 19964
rect 8092 20018 8148 20748
rect 8540 20804 8596 22206
rect 8540 20738 8596 20748
rect 9324 20804 9380 20814
rect 9324 20710 9380 20748
rect 8820 20244 8876 20254
rect 8820 20150 8876 20188
rect 8092 19966 8094 20018
rect 8146 19966 8148 20018
rect 8092 19954 8148 19966
rect 8484 20020 8540 20030
rect 8988 20020 9044 20030
rect 8484 20018 9044 20020
rect 8484 19966 8486 20018
rect 8538 19966 8990 20018
rect 9042 19966 9044 20018
rect 8484 19964 9044 19966
rect 8484 19954 8540 19964
rect 8316 19908 8372 19918
rect 8204 19906 8372 19908
rect 8204 19854 8318 19906
rect 8370 19854 8372 19906
rect 8204 19852 8372 19854
rect 8204 19572 8260 19852
rect 8316 19842 8372 19852
rect 7308 19516 8260 19572
rect 7308 18450 7364 19516
rect 8988 19348 9044 19964
rect 9324 19348 9380 19358
rect 8988 19346 9380 19348
rect 8988 19294 9326 19346
rect 9378 19294 9380 19346
rect 8988 19292 9380 19294
rect 9324 19282 9380 19292
rect 7420 19236 7476 19246
rect 7420 19234 7700 19236
rect 7420 19182 7422 19234
rect 7474 19182 7700 19234
rect 7420 19180 7700 19182
rect 7420 19170 7476 19180
rect 7644 18788 7700 19180
rect 7644 18732 8148 18788
rect 8092 18674 8148 18732
rect 7308 18398 7310 18450
rect 7362 18398 7364 18450
rect 7308 18386 7364 18398
rect 7420 18618 7476 18630
rect 7420 18566 7422 18618
rect 7474 18566 7476 18618
rect 8092 18622 8094 18674
rect 8146 18622 8148 18674
rect 8092 18610 8148 18622
rect 7420 18452 7476 18566
rect 7756 18452 7812 18462
rect 7420 18450 7812 18452
rect 7420 18398 7758 18450
rect 7810 18398 7812 18450
rect 7420 18396 7812 18398
rect 7756 18386 7812 18396
rect 7644 18228 7700 18238
rect 7644 17890 7700 18172
rect 7644 17838 7646 17890
rect 7698 17838 7700 17890
rect 7644 17826 7700 17838
rect 8316 17780 8372 17790
rect 7308 17668 7364 17678
rect 7196 17666 7364 17668
rect 7196 17614 7310 17666
rect 7362 17614 7364 17666
rect 7196 17612 7364 17614
rect 6748 16772 6804 16782
rect 6748 16678 6804 16716
rect 6524 16492 6748 16548
rect 6692 16154 6748 16492
rect 6300 15358 6356 15932
rect 5964 15316 6020 15326
rect 5740 15314 6020 15316
rect 5740 15262 5966 15314
rect 6018 15262 6020 15314
rect 6300 15306 6302 15358
rect 6354 15306 6356 15358
rect 6300 15294 6356 15306
rect 6524 16098 6580 16110
rect 6524 16046 6526 16098
rect 6578 16046 6580 16098
rect 6692 16102 6694 16154
rect 6746 16102 6748 16154
rect 6692 16090 6748 16102
rect 6972 16098 7028 17052
rect 7084 16884 7140 16894
rect 7196 16884 7252 17612
rect 7308 17602 7364 17612
rect 8316 17651 8372 17724
rect 8988 17780 9044 17790
rect 8988 17686 9044 17724
rect 8316 17599 8318 17651
rect 8370 17599 8372 17651
rect 8652 17668 8708 17678
rect 8876 17668 8932 17678
rect 8652 17666 8876 17668
rect 8652 17614 8654 17666
rect 8706 17614 8876 17666
rect 8652 17612 8876 17614
rect 9324 17666 9380 17678
rect 8652 17602 8708 17612
rect 8316 17587 8372 17599
rect 8428 17498 8484 17510
rect 8428 17446 8430 17498
rect 8482 17446 8484 17498
rect 7084 16882 7252 16884
rect 7084 16830 7086 16882
rect 7138 16830 7252 16882
rect 7084 16828 7252 16830
rect 7420 16996 7476 17006
rect 7420 16882 7476 16940
rect 7420 16830 7422 16882
rect 7474 16830 7476 16882
rect 7084 16818 7140 16828
rect 7420 16818 7476 16830
rect 8204 16882 8260 16894
rect 8204 16830 8206 16882
rect 8258 16830 8260 16882
rect 8204 16772 8260 16830
rect 8428 16882 8484 17446
rect 8428 16830 8430 16882
rect 8482 16830 8484 16882
rect 8428 16818 8484 16830
rect 8540 17108 8596 17118
rect 8204 16706 8260 16716
rect 5740 15260 6020 15262
rect 5964 15250 6020 15260
rect 6412 15204 6468 15242
rect 6412 15138 6468 15148
rect 5964 14868 6020 14878
rect 5964 14530 6020 14812
rect 6524 14868 6580 16046
rect 6972 16046 6974 16098
rect 7026 16046 7028 16098
rect 6972 16034 7028 16046
rect 7084 16660 7140 16670
rect 6860 15986 6916 15998
rect 6860 15934 6862 15986
rect 6914 15934 6916 15986
rect 6860 15204 6916 15934
rect 6972 15316 7028 15326
rect 6972 15222 7028 15260
rect 6860 15138 6916 15148
rect 7084 15092 7140 16604
rect 8540 16210 8596 17052
rect 8708 16996 8764 17006
rect 8876 16996 8932 17612
rect 9100 17622 9156 17634
rect 9100 17570 9102 17622
rect 9154 17570 9156 17622
rect 9100 17444 9156 17570
rect 9100 17378 9156 17388
rect 9324 17614 9326 17666
rect 9378 17614 9380 17666
rect 9324 17108 9380 17614
rect 9548 17668 9604 22652
rect 9660 22372 9716 22382
rect 9660 22370 9940 22372
rect 9660 22318 9662 22370
rect 9714 22318 9940 22370
rect 9660 22316 9940 22318
rect 9660 22306 9716 22316
rect 9884 21810 9940 22316
rect 9884 21758 9886 21810
rect 9938 21758 9940 21810
rect 9884 21746 9940 21758
rect 10220 22148 10276 22158
rect 10220 21586 10276 22092
rect 10220 21534 10222 21586
rect 10274 21534 10276 21586
rect 10220 21522 10276 21534
rect 10892 21586 10948 22876
rect 11228 22372 11284 24670
rect 11340 24724 11396 27132
rect 11452 27074 11508 27086
rect 11452 27022 11454 27074
rect 11506 27022 11508 27074
rect 11452 26516 11508 27022
rect 11564 26908 11620 29036
rect 11676 29036 11844 29092
rect 12124 29426 12180 29438
rect 12124 29374 12126 29426
rect 12178 29374 12180 29426
rect 11676 28644 11732 29036
rect 12124 28754 12180 29374
rect 12348 29413 12350 29465
rect 12402 29413 12404 29465
rect 12348 28868 12404 29413
rect 12684 29204 12740 29542
rect 12796 29426 12852 29820
rect 12796 29374 12798 29426
rect 12850 29374 12852 29426
rect 12796 29362 12852 29374
rect 12684 29138 12740 29148
rect 12348 28802 12404 28812
rect 12124 28702 12126 28754
rect 12178 28702 12180 28754
rect 12124 28690 12180 28702
rect 11676 28550 11732 28588
rect 11900 28642 11956 28654
rect 11900 28590 11902 28642
rect 11954 28590 11956 28642
rect 11900 28532 11956 28590
rect 12236 28644 12292 28654
rect 12236 28575 12238 28588
rect 12290 28575 12292 28588
rect 12236 28550 12292 28575
rect 12460 28642 12516 28654
rect 12460 28590 12462 28642
rect 12514 28590 12516 28642
rect 11676 27524 11732 27534
rect 11676 27186 11732 27468
rect 11900 27412 11956 28476
rect 12460 28532 12516 28590
rect 12460 28466 12516 28476
rect 12908 28084 12964 33068
rect 13020 32564 13076 34076
rect 13020 32498 13076 32508
rect 13244 32577 13300 32589
rect 13244 32525 13246 32577
rect 13298 32525 13300 32577
rect 13132 32450 13188 32462
rect 13132 32398 13134 32450
rect 13186 32398 13188 32450
rect 13020 31778 13076 31790
rect 13020 31726 13022 31778
rect 13074 31726 13076 31778
rect 13020 31668 13076 31726
rect 13132 31780 13188 32398
rect 13244 32340 13300 32525
rect 13244 32274 13300 32284
rect 13356 31948 13412 34412
rect 13468 35698 13524 35710
rect 13468 35646 13470 35698
rect 13522 35646 13524 35698
rect 13468 34132 13524 35646
rect 14252 35698 14308 36652
rect 14924 36642 14980 36652
rect 14588 36484 14644 36494
rect 14252 35646 14254 35698
rect 14306 35646 14308 35698
rect 14252 35634 14308 35646
rect 14476 36482 14644 36484
rect 14476 36430 14590 36482
rect 14642 36430 14644 36482
rect 14476 36428 14644 36430
rect 14252 35476 14308 35486
rect 14252 34916 14308 35420
rect 14476 35150 14532 36428
rect 14588 36418 14644 36428
rect 15372 36484 15428 36494
rect 15148 35364 15204 35374
rect 14420 35138 14532 35150
rect 14420 35086 14422 35138
rect 14474 35086 14532 35138
rect 14420 35084 14532 35086
rect 14924 35252 14980 35262
rect 14420 35074 14476 35084
rect 14252 34879 14700 34916
rect 14252 34860 14646 34879
rect 14644 34827 14646 34860
rect 14698 34827 14700 34879
rect 14644 34815 14700 34827
rect 14924 34886 14980 35196
rect 14924 34834 14926 34886
rect 14978 34834 14980 34886
rect 14924 34822 14980 34834
rect 15148 34886 15204 35308
rect 15372 35252 15428 36428
rect 15932 35812 15988 38108
rect 16044 38052 16100 38062
rect 16044 37268 16100 37996
rect 16716 37828 16772 38782
rect 16940 38834 16996 38846
rect 16940 38782 16942 38834
rect 16994 38782 16996 38834
rect 16940 38612 16996 38782
rect 17556 38722 17612 38734
rect 17556 38670 17558 38722
rect 17610 38670 17612 38722
rect 17556 38668 17612 38670
rect 17948 38722 18004 38734
rect 17948 38670 17950 38722
rect 18002 38670 18004 38722
rect 17556 38612 17892 38668
rect 16940 38276 16996 38556
rect 16828 38220 16996 38276
rect 16828 38022 16884 38220
rect 17500 38164 17556 38174
rect 17388 38052 17444 38062
rect 16828 37970 16830 38022
rect 16882 37970 16884 38022
rect 16828 37958 16884 37970
rect 16940 38015 17052 38052
rect 16940 37963 16998 38015
rect 17050 37963 17052 38015
rect 16940 37951 17052 37963
rect 17276 37994 17332 38006
rect 16940 37828 16996 37951
rect 16716 37772 16996 37828
rect 17276 37942 17278 37994
rect 17330 37942 17332 37994
rect 17500 38052 17556 38108
rect 17612 38052 17668 38062
rect 17500 38050 17668 38052
rect 17500 37998 17614 38050
rect 17666 37998 17668 38050
rect 17500 37996 17668 37998
rect 17836 38052 17892 38612
rect 17948 38612 18004 38670
rect 17948 38276 18004 38556
rect 17948 38210 18004 38220
rect 18396 38052 18452 41916
rect 18508 39564 18564 43260
rect 18732 42866 18788 43260
rect 19068 43250 19124 43260
rect 18732 42814 18734 42866
rect 18786 42814 18788 42866
rect 18732 42802 18788 42814
rect 18956 43092 19012 43102
rect 19404 43092 19460 43486
rect 19516 43540 19572 43652
rect 19628 43652 19684 44044
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19628 43596 19964 43652
rect 19908 43594 19964 43596
rect 19908 43542 19910 43594
rect 19962 43542 19964 43594
rect 19516 43484 19740 43540
rect 19908 43530 19964 43542
rect 20188 43566 20244 44214
rect 19684 43426 19740 43484
rect 19684 43374 19686 43426
rect 19738 43374 19740 43426
rect 19684 43362 19740 43374
rect 20188 43514 20190 43566
rect 20242 43514 20244 43566
rect 19404 43036 19908 43092
rect 18956 42082 19012 43036
rect 19852 42532 19908 43036
rect 19628 42476 19908 42532
rect 19628 42196 19684 42476
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 20076 42196 20132 42206
rect 19628 42140 19852 42196
rect 18956 42030 18958 42082
rect 19010 42030 19012 42082
rect 18956 42018 19012 42030
rect 19796 42082 19852 42140
rect 19796 42030 19798 42082
rect 19850 42030 19852 42082
rect 19796 42018 19852 42030
rect 20076 42026 20132 42140
rect 18620 41972 18676 41982
rect 19068 41970 19124 41982
rect 18620 41878 18676 41916
rect 18788 41914 18844 41926
rect 18788 41862 18790 41914
rect 18842 41862 18844 41914
rect 18788 41412 18844 41862
rect 18788 41346 18844 41356
rect 19068 41918 19070 41970
rect 19122 41918 19124 41970
rect 20076 41974 20078 42026
rect 20130 41974 20132 42026
rect 20076 41962 20132 41974
rect 20188 42038 20244 43514
rect 20412 44266 20468 44278
rect 20412 44214 20414 44266
rect 20466 44214 20468 44266
rect 20524 44235 20526 44287
rect 20578 44235 20580 44287
rect 20524 44223 20580 44235
rect 20412 43566 20468 44214
rect 20636 44100 20692 45726
rect 20748 47234 20972 47236
rect 20748 47182 20918 47234
rect 20970 47182 20972 47234
rect 20748 47180 20972 47182
rect 20748 44660 20804 47180
rect 20916 47170 20972 47180
rect 20972 46676 21028 46686
rect 21084 46676 21140 47516
rect 21196 47458 21252 47740
rect 22652 47628 23492 47684
rect 22428 47572 22484 47582
rect 22428 47478 22484 47516
rect 22652 47460 22708 47628
rect 21196 47406 21198 47458
rect 21250 47406 21252 47458
rect 21196 47394 21252 47406
rect 22596 47404 22708 47460
rect 22764 47460 22820 47470
rect 23100 47460 23156 47470
rect 22596 47402 22652 47404
rect 22596 47350 22598 47402
rect 22650 47350 22652 47402
rect 22596 47338 22652 47350
rect 21364 47236 21420 47246
rect 20972 46674 21140 46676
rect 20972 46622 20974 46674
rect 21026 46622 21140 46674
rect 20972 46620 21140 46622
rect 21196 47234 21420 47236
rect 21196 47182 21366 47234
rect 21418 47182 21420 47234
rect 21196 47180 21420 47182
rect 20972 46610 21028 46620
rect 21196 45108 21252 47180
rect 21364 47170 21420 47180
rect 21924 47236 21980 47246
rect 21924 47234 22148 47236
rect 21924 47182 21926 47234
rect 21978 47182 22148 47234
rect 21924 47180 22148 47182
rect 21924 47170 21980 47180
rect 21308 45890 21364 45902
rect 21308 45838 21310 45890
rect 21362 45838 21364 45890
rect 21308 45332 21364 45838
rect 21308 45108 21364 45276
rect 21532 45108 21588 45118
rect 22092 45108 22148 47180
rect 22764 46452 22820 47404
rect 22876 47458 23156 47460
rect 22876 47406 23102 47458
rect 23154 47406 23156 47458
rect 22876 47404 23156 47406
rect 22876 46786 22932 47404
rect 23100 47394 23156 47404
rect 23268 47236 23324 47246
rect 23268 47142 23324 47180
rect 22876 46734 22878 46786
rect 22930 46734 22932 46786
rect 22876 46722 22932 46734
rect 23436 46786 23492 47628
rect 26236 47628 26516 47684
rect 24892 47460 24948 47470
rect 24668 47414 24724 47426
rect 24668 47362 24670 47414
rect 24722 47362 24724 47414
rect 24892 47366 24948 47404
rect 26236 47458 26292 47628
rect 26236 47406 26238 47458
rect 26290 47406 26292 47458
rect 26236 47394 26292 47406
rect 26348 47458 26404 47470
rect 26348 47406 26350 47458
rect 26402 47406 26404 47458
rect 23436 46734 23438 46786
rect 23490 46734 23492 46786
rect 23436 46722 23492 46734
rect 23884 47236 23940 47246
rect 23679 46674 23735 46686
rect 23679 46622 23681 46674
rect 23733 46622 23735 46674
rect 23679 46564 23735 46622
rect 23679 46508 23828 46564
rect 22764 46396 23156 46452
rect 22652 46004 22708 46014
rect 22540 46002 22708 46004
rect 22540 45950 22654 46002
rect 22706 45950 22708 46002
rect 22540 45948 22708 45950
rect 21308 45106 21588 45108
rect 21308 45054 21534 45106
rect 21586 45054 21588 45106
rect 21308 45052 21588 45054
rect 21196 45042 21252 45052
rect 20748 44436 20804 44604
rect 20748 44370 20804 44380
rect 21084 44994 21140 45006
rect 21084 44942 21086 44994
rect 21138 44942 21140 44994
rect 21084 44324 21140 44942
rect 21532 44436 21588 45052
rect 21532 44370 21588 44380
rect 21756 45052 22148 45108
rect 22316 45108 22372 45118
rect 22540 45108 22596 45948
rect 22652 45938 22708 45948
rect 23100 45892 23156 46396
rect 23100 45890 23492 45892
rect 22764 45846 22820 45858
rect 22764 45794 22766 45846
rect 22818 45794 22820 45846
rect 23100 45838 23102 45890
rect 23154 45838 23492 45890
rect 23100 45836 23492 45838
rect 23100 45826 23156 45836
rect 22764 45332 22820 45794
rect 22764 45266 22820 45276
rect 22316 45106 22596 45108
rect 22316 45054 22318 45106
rect 22370 45054 22596 45106
rect 22316 45052 22596 45054
rect 21756 44296 21812 45052
rect 22316 45042 22372 45052
rect 21084 44258 21140 44268
rect 21308 44294 21812 44296
rect 20636 44034 20692 44044
rect 21308 44242 21758 44294
rect 21810 44242 21812 44294
rect 21308 44240 21812 44242
rect 20636 43764 20692 43774
rect 20636 43606 20692 43708
rect 20412 43514 20414 43566
rect 20466 43514 20468 43566
rect 20599 43594 20692 43606
rect 20599 43542 20601 43594
rect 20653 43542 20692 43594
rect 20599 43540 20692 43542
rect 20599 43530 20655 43540
rect 20188 42026 20300 42038
rect 20188 41974 20246 42026
rect 20298 41974 20300 42026
rect 20188 41962 20300 41974
rect 20412 42028 20468 43514
rect 20748 43428 20804 43438
rect 20636 42756 20692 42766
rect 20636 42642 20692 42700
rect 20636 42590 20638 42642
rect 20690 42590 20692 42642
rect 20636 42196 20692 42590
rect 20636 42130 20692 42140
rect 20748 42038 20804 43372
rect 21028 43428 21084 43438
rect 21028 43334 21084 43372
rect 21196 42756 21252 42766
rect 21308 42756 21364 44240
rect 21756 44230 21812 44240
rect 22764 44772 22820 44782
rect 23436 44772 23492 45836
rect 21644 44100 21700 44110
rect 21532 43540 21588 43550
rect 21532 43446 21588 43484
rect 21308 42700 21588 42756
rect 21196 42662 21252 42700
rect 21364 42532 21420 42542
rect 21364 42438 21420 42476
rect 20412 41998 20580 42028
rect 20412 41972 20526 41998
rect 19068 40852 19124 41918
rect 19348 41748 19404 41758
rect 19348 41746 19460 41748
rect 19348 41694 19350 41746
rect 19402 41694 19460 41746
rect 19348 41682 19460 41694
rect 19068 40786 19124 40796
rect 19292 39844 19348 39854
rect 19404 39844 19460 41682
rect 19964 41188 20020 41198
rect 19348 39788 19460 39844
rect 19516 41186 20020 41188
rect 19516 41134 19966 41186
rect 20018 41134 20020 41186
rect 19516 41132 20020 41134
rect 19516 39844 19572 41132
rect 19964 41122 20020 41132
rect 19628 40962 19684 40974
rect 19628 40910 19630 40962
rect 19682 40910 19684 40962
rect 19628 40402 19684 40910
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19628 40350 19630 40402
rect 19682 40350 19684 40402
rect 19628 40338 19684 40350
rect 19964 40404 20020 40414
rect 19684 39844 19740 39854
rect 19516 39842 19740 39844
rect 19516 39790 19686 39842
rect 19738 39790 19740 39842
rect 19516 39788 19740 39790
rect 19292 39778 19348 39788
rect 19684 39778 19740 39788
rect 19404 39620 19460 39630
rect 18508 39508 18676 39564
rect 19404 39526 19460 39564
rect 19964 39590 20020 40348
rect 19964 39538 19966 39590
rect 20018 39538 20020 39590
rect 19964 39526 20020 39538
rect 20188 39562 20244 41962
rect 20524 41946 20526 41972
rect 20578 41946 20580 41998
rect 20711 42026 20804 42038
rect 20711 41974 20713 42026
rect 20765 41974 20804 42026
rect 20711 41972 20804 41974
rect 20711 41962 20767 41972
rect 20524 41636 20580 41946
rect 21140 41860 21196 41870
rect 21084 41858 21196 41860
rect 21084 41806 21142 41858
rect 21194 41806 21196 41858
rect 21084 41794 21196 41806
rect 20524 41580 20692 41636
rect 20524 41188 20580 41198
rect 20356 40964 20412 40974
rect 20356 40870 20412 40908
rect 20412 40404 20468 40414
rect 20524 40404 20580 41132
rect 20636 40740 20692 41580
rect 20804 40964 20860 40974
rect 20804 40962 21028 40964
rect 20804 40910 20806 40962
rect 20858 40910 21028 40962
rect 20804 40908 21028 40910
rect 20804 40898 20860 40908
rect 20636 40684 20916 40740
rect 20748 40516 20804 40526
rect 20748 40422 20804 40460
rect 20412 40402 20692 40404
rect 20412 40350 20414 40402
rect 20466 40350 20692 40402
rect 20412 40348 20692 40350
rect 20412 40338 20468 40348
rect 18508 39396 18564 39406
rect 18508 39302 18564 39340
rect 18620 38164 18676 39508
rect 19068 39508 19124 39518
rect 19068 39414 19124 39452
rect 20188 39510 20190 39562
rect 20242 39510 20244 39562
rect 20188 39508 20244 39510
rect 20188 39442 20244 39452
rect 20300 39620 20356 39630
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19852 38722 19908 38734
rect 19852 38670 19854 38722
rect 19906 38670 19908 38722
rect 19852 38500 19908 38670
rect 18620 38098 18676 38108
rect 18732 38444 19908 38500
rect 19964 38724 20020 38734
rect 18732 38162 18788 38444
rect 18732 38110 18734 38162
rect 18786 38110 18788 38162
rect 18732 38098 18788 38110
rect 18844 38164 18900 38174
rect 19964 38164 20020 38668
rect 20300 38724 20356 39564
rect 20412 39562 20468 39574
rect 20412 39510 20414 39562
rect 20466 39510 20468 39562
rect 20412 39396 20468 39510
rect 20524 39562 20580 39574
rect 20524 39510 20526 39562
rect 20578 39510 20580 39562
rect 20524 39508 20580 39510
rect 20524 39442 20580 39452
rect 20412 39330 20468 39340
rect 20636 38834 20692 40348
rect 20860 39396 20916 40684
rect 20860 39330 20916 39340
rect 20972 39284 21028 40908
rect 21084 39508 21140 41794
rect 21084 39442 21140 39452
rect 21196 41300 21252 41310
rect 21196 39284 21252 41244
rect 21420 41188 21476 41198
rect 20972 39218 21028 39228
rect 21084 39228 21252 39284
rect 21308 39284 21364 39294
rect 20636 38782 20638 38834
rect 20690 38782 20692 38834
rect 20972 39060 21028 39070
rect 20972 38878 21028 39004
rect 20972 38826 20974 38878
rect 21026 38826 21028 38878
rect 20972 38814 21028 38826
rect 20636 38770 20692 38782
rect 20300 38658 20356 38668
rect 20860 38724 20916 38734
rect 20860 38630 20916 38668
rect 17836 37996 18004 38052
rect 17388 37963 17390 37996
rect 17442 37963 17444 37996
rect 17612 37986 17668 37996
rect 17388 37951 17444 37963
rect 17276 37828 17332 37942
rect 17780 37828 17836 37838
rect 17276 37826 17836 37828
rect 17276 37774 17782 37826
rect 17834 37774 17836 37826
rect 17276 37772 17836 37774
rect 16716 37502 16772 37772
rect 17780 37762 17836 37772
rect 16716 37490 16828 37502
rect 16716 37438 16774 37490
rect 16826 37438 16828 37490
rect 16716 37436 16828 37438
rect 16772 37426 16828 37436
rect 17500 37380 17556 37390
rect 17500 37286 17556 37324
rect 17743 37380 17799 37390
rect 17743 37322 17799 37324
rect 16156 37268 16212 37278
rect 16044 37266 16212 37268
rect 16044 37214 16158 37266
rect 16210 37214 16212 37266
rect 16044 37212 16212 37214
rect 16156 37202 16212 37212
rect 16940 37266 16996 37278
rect 16940 37214 16942 37266
rect 16994 37214 16996 37266
rect 17743 37270 17745 37322
rect 17797 37270 17799 37322
rect 17743 37258 17799 37270
rect 17948 37380 18004 37996
rect 18396 37958 18452 37996
rect 18620 38006 18676 38018
rect 18620 37954 18622 38006
rect 18674 37954 18676 38006
rect 18620 37492 18676 37954
rect 18620 37426 18676 37436
rect 16940 36596 16996 37214
rect 17836 37044 17892 37054
rect 17724 36596 17780 36606
rect 16940 36594 17780 36596
rect 16940 36542 17726 36594
rect 17778 36542 17780 36594
rect 16940 36540 17780 36542
rect 16716 36484 16772 36494
rect 16380 36426 16436 36438
rect 16380 36374 16382 36426
rect 16434 36374 16436 36426
rect 16100 36260 16156 36270
rect 16380 36260 16436 36374
rect 16100 36258 16436 36260
rect 16100 36206 16102 36258
rect 16154 36206 16436 36258
rect 16100 36204 16436 36206
rect 16100 36194 16156 36204
rect 16156 35812 16212 35822
rect 15932 35810 16212 35812
rect 15932 35758 16158 35810
rect 16210 35758 16212 35810
rect 15932 35756 16212 35758
rect 15932 35476 15988 35756
rect 16156 35746 16212 35756
rect 16380 35588 16436 36204
rect 16380 35522 16436 35532
rect 16492 36426 16548 36438
rect 16492 36374 16494 36426
rect 16546 36374 16548 36426
rect 16716 36402 16718 36428
rect 16770 36402 16772 36428
rect 16716 36390 16772 36402
rect 16940 36454 16996 36540
rect 17724 36530 17780 36540
rect 16940 36402 16942 36454
rect 16994 36402 16996 36454
rect 16940 36390 16996 36402
rect 16492 35924 16548 36374
rect 15932 35410 15988 35420
rect 16492 35364 16548 35868
rect 17220 36370 17276 36382
rect 17220 36318 17222 36370
rect 17274 36318 17276 36370
rect 17220 35812 17276 36318
rect 17220 35746 17276 35756
rect 17500 35698 17556 35710
rect 17500 35646 17502 35698
rect 17554 35646 17556 35698
rect 16492 35298 16548 35308
rect 16884 35586 16940 35598
rect 16884 35534 16886 35586
rect 16938 35534 16940 35586
rect 16884 35364 16940 35534
rect 16884 35298 16940 35308
rect 17500 35364 17556 35646
rect 17500 35298 17556 35308
rect 17724 35698 17780 35710
rect 17724 35646 17726 35698
rect 17778 35646 17780 35698
rect 15372 35186 15428 35196
rect 15148 34834 15150 34886
rect 15202 34834 15204 34886
rect 15820 34914 15876 34926
rect 15148 34822 15204 34834
rect 15260 34858 15316 34870
rect 15260 34806 15262 34858
rect 15314 34806 15316 34858
rect 15260 34692 15316 34806
rect 15820 34862 15822 34914
rect 15874 34862 15876 34914
rect 15652 34692 15708 34702
rect 15260 34626 15316 34636
rect 15596 34690 15708 34692
rect 15596 34638 15654 34690
rect 15706 34638 15708 34690
rect 15596 34626 15708 34638
rect 13468 34066 13524 34076
rect 13804 34018 13860 34030
rect 13804 33966 13806 34018
rect 13858 33966 13860 34018
rect 13804 33796 13860 33966
rect 13804 33730 13860 33740
rect 15036 33514 15092 33526
rect 15036 33462 15038 33514
rect 15090 33462 15092 33514
rect 13580 33348 13636 33358
rect 14700 33346 14756 33358
rect 13580 33254 13636 33292
rect 13823 33290 13879 33302
rect 13823 33238 13825 33290
rect 13877 33238 13879 33290
rect 13580 33124 13636 33134
rect 13580 32562 13636 33068
rect 13823 32788 13879 33238
rect 14700 33294 14702 33346
rect 14754 33294 14756 33346
rect 14700 33124 14756 33294
rect 14700 33058 14756 33068
rect 13580 32510 13582 32562
rect 13634 32510 13636 32562
rect 13580 32498 13636 32510
rect 13804 32732 13879 32788
rect 13804 32340 13860 32732
rect 13804 32274 13860 32284
rect 14252 32676 14308 32686
rect 13132 31714 13188 31724
rect 13244 31892 13412 31948
rect 13020 31602 13076 31612
rect 13244 31220 13300 31892
rect 13356 31778 13412 31790
rect 13356 31726 13358 31778
rect 13410 31726 13412 31778
rect 14252 31750 14308 32620
rect 15036 32676 15092 33462
rect 15148 33348 15204 33358
rect 15148 33254 15204 33292
rect 15484 33348 15540 33358
rect 15596 33348 15652 34626
rect 15820 34356 15876 34862
rect 17500 34914 17556 34926
rect 17500 34862 17502 34914
rect 17554 34862 17556 34914
rect 15484 33346 15652 33348
rect 15484 33294 15486 33346
rect 15538 33294 15652 33346
rect 15484 33292 15652 33294
rect 15708 34300 15876 34356
rect 16156 34692 16268 34702
rect 16212 34690 16268 34692
rect 16212 34638 16214 34690
rect 16266 34638 16268 34690
rect 16212 34636 16268 34638
rect 16156 34626 16268 34636
rect 16492 34692 16548 34702
rect 15708 34018 15764 34300
rect 15708 33966 15710 34018
rect 15762 33966 15764 34018
rect 15484 33124 15540 33292
rect 15484 33058 15540 33068
rect 15708 33012 15764 33966
rect 15708 32946 15764 32956
rect 15820 34132 15876 34142
rect 15820 33346 15876 34076
rect 15820 33294 15822 33346
rect 15874 33294 15876 33346
rect 15036 32610 15092 32620
rect 14364 32589 14420 32602
rect 14364 32564 14366 32589
rect 14418 32564 14420 32589
rect 14364 32498 14420 32508
rect 15820 32564 15876 33294
rect 15820 32498 15876 32508
rect 16156 32340 16212 34626
rect 16380 34130 16436 34142
rect 16380 34078 16382 34130
rect 16434 34078 16436 34130
rect 16380 33908 16436 34078
rect 16380 33236 16436 33852
rect 16268 32564 16324 32574
rect 16268 32470 16324 32508
rect 16156 32284 16324 32340
rect 13356 31444 13412 31726
rect 13916 31722 13972 31734
rect 13916 31670 13918 31722
rect 13970 31670 13972 31722
rect 13916 31668 13972 31670
rect 13916 31602 13972 31612
rect 14028 31722 14084 31734
rect 14028 31670 14030 31722
rect 14082 31670 14084 31722
rect 14252 31698 14254 31750
rect 14306 31698 14308 31750
rect 14252 31686 14308 31698
rect 14476 31892 14532 31902
rect 14476 31750 14532 31836
rect 14476 31698 14478 31750
rect 14530 31698 14532 31750
rect 14476 31686 14532 31698
rect 13356 31378 13412 31388
rect 13524 31554 13580 31566
rect 13524 31502 13526 31554
rect 13578 31502 13580 31554
rect 13132 31164 13300 31220
rect 13020 31022 13076 31034
rect 13020 30970 13022 31022
rect 13074 30970 13076 31022
rect 13020 30772 13076 30970
rect 13020 30706 13076 30716
rect 12908 28028 13076 28084
rect 11900 27346 11956 27356
rect 12460 27412 12516 27422
rect 11676 27134 11678 27186
rect 11730 27134 11732 27186
rect 11676 27122 11732 27134
rect 11788 27076 11844 27086
rect 11788 26982 11844 27020
rect 12460 27074 12516 27356
rect 12852 27300 12908 27310
rect 12852 27206 12908 27244
rect 12460 27022 12462 27074
rect 12514 27022 12516 27074
rect 12460 27010 12516 27022
rect 12572 27076 12628 27086
rect 12572 26982 12628 27020
rect 11956 26964 12012 26974
rect 11564 26852 11732 26908
rect 11452 26450 11508 26460
rect 11508 26292 11564 26302
rect 11508 25730 11564 26236
rect 11508 25678 11510 25730
rect 11562 25678 11564 25730
rect 11508 25666 11564 25678
rect 11340 24658 11396 24668
rect 11676 24836 11732 26852
rect 11788 26628 11844 26638
rect 11788 26290 11844 26572
rect 11956 26514 12012 26908
rect 11956 26462 11958 26514
rect 12010 26462 12012 26514
rect 11956 26450 12012 26462
rect 12236 26292 12292 26302
rect 11788 26238 11790 26290
rect 11842 26238 11844 26290
rect 11788 25478 11844 26238
rect 11788 25426 11790 25478
rect 11842 25426 11844 25478
rect 12124 26290 12292 26292
rect 12124 26238 12238 26290
rect 12290 26238 12292 26290
rect 12124 26236 12292 26238
rect 11788 25414 11844 25426
rect 12012 25450 12068 25462
rect 12012 25398 12014 25450
rect 12066 25398 12068 25450
rect 12012 25172 12068 25398
rect 12012 25106 12068 25116
rect 11676 24052 11732 24780
rect 12012 24948 12068 24958
rect 12012 24722 12068 24892
rect 12012 24670 12014 24722
rect 12066 24670 12068 24722
rect 12012 24658 12068 24670
rect 12124 24174 12180 26236
rect 12236 26226 12292 26236
rect 12572 26066 12628 26078
rect 12572 26014 12574 26066
rect 12626 26014 12628 26066
rect 12236 25564 12516 25620
rect 12236 25478 12292 25564
rect 12236 25426 12238 25478
rect 12290 25426 12292 25478
rect 12236 25414 12292 25426
rect 12348 25450 12404 25462
rect 12348 25398 12350 25450
rect 12402 25398 12404 25450
rect 12348 25284 12404 25398
rect 12348 25218 12404 25228
rect 12068 24162 12180 24174
rect 12068 24110 12070 24162
rect 12122 24110 12180 24162
rect 12068 24108 12180 24110
rect 12236 25172 12292 25182
rect 12068 24098 12124 24108
rect 11676 23986 11732 23996
rect 12236 23940 12292 25116
rect 12460 25060 12516 25564
rect 12460 24994 12516 25004
rect 12572 24948 12628 26014
rect 13020 25396 13076 28028
rect 13132 25508 13188 31164
rect 13244 31022 13300 31034
rect 13244 30970 13246 31022
rect 13298 30970 13300 31022
rect 13244 30436 13300 30970
rect 13356 31029 13412 31041
rect 13356 30996 13358 31029
rect 13410 30996 13412 31029
rect 13356 30930 13412 30940
rect 13524 30996 13580 31502
rect 14028 31220 14084 31670
rect 14756 31668 14812 31678
rect 14028 31154 14084 31164
rect 14700 31666 14812 31668
rect 14700 31614 14758 31666
rect 14810 31614 14812 31666
rect 14700 31602 14812 31614
rect 15596 31668 15652 31678
rect 13524 30930 13580 30940
rect 13692 30994 13748 31006
rect 14028 30996 14084 31006
rect 13692 30942 13694 30994
rect 13746 30942 13748 30994
rect 13692 30884 13748 30942
rect 13692 30818 13748 30828
rect 13916 30994 14084 30996
rect 13916 30942 14030 30994
rect 14082 30942 14084 30994
rect 13916 30940 14084 30942
rect 13244 30370 13300 30380
rect 13916 30772 13972 30940
rect 14028 30930 14084 30940
rect 14588 30994 14644 31006
rect 14588 30942 14590 30994
rect 14642 30942 14644 30994
rect 13916 30210 13972 30716
rect 14588 30436 14644 30942
rect 14588 30370 14644 30380
rect 13916 30158 13918 30210
rect 13970 30158 13972 30210
rect 13356 29204 13412 29214
rect 13244 28644 13300 28654
rect 13244 27858 13300 28588
rect 13356 28642 13412 29148
rect 13356 28590 13358 28642
rect 13410 28590 13412 28642
rect 13356 28578 13412 28590
rect 13692 28644 13748 28654
rect 13692 28550 13748 28588
rect 13244 27806 13246 27858
rect 13298 27806 13300 27858
rect 13244 27794 13300 27806
rect 13468 27188 13524 27198
rect 13300 27076 13356 27086
rect 13300 26514 13356 27020
rect 13468 27039 13524 27132
rect 13468 26987 13470 27039
rect 13522 26987 13524 27039
rect 13804 27076 13860 27086
rect 13468 26975 13524 26987
rect 13580 27018 13636 27030
rect 13580 26966 13582 27018
rect 13634 26966 13636 27018
rect 13804 26994 13806 27020
rect 13858 26994 13860 27020
rect 13804 26982 13860 26994
rect 13580 26964 13636 26966
rect 13580 26898 13636 26908
rect 13300 26462 13302 26514
rect 13354 26462 13356 26514
rect 13300 26450 13356 26462
rect 13692 26516 13748 26526
rect 13692 26346 13748 26460
rect 13468 26290 13524 26302
rect 13468 26238 13470 26290
rect 13522 26238 13524 26290
rect 13692 26294 13694 26346
rect 13746 26294 13748 26346
rect 13916 26516 13972 30158
rect 14700 30212 14756 31602
rect 14924 31220 14980 31230
rect 14812 30996 14868 31006
rect 14812 30902 14868 30940
rect 14700 30175 14812 30212
rect 14700 30156 14758 30175
rect 14756 30123 14758 30156
rect 14810 30123 14812 30175
rect 14756 30111 14812 30123
rect 14084 30100 14140 30110
rect 14084 30042 14140 30044
rect 14084 29990 14086 30042
rect 14138 29990 14140 30042
rect 14532 30100 14588 30110
rect 14532 30098 14644 30100
rect 14532 30046 14534 30098
rect 14586 30046 14644 30098
rect 14532 30034 14644 30046
rect 14084 29978 14140 29990
rect 14476 28644 14532 28654
rect 14364 27972 14420 27982
rect 14028 27860 14084 27870
rect 14028 27766 14084 27804
rect 14028 27412 14084 27422
rect 14028 27046 14084 27356
rect 14364 27310 14420 27916
rect 14308 27298 14420 27310
rect 14308 27246 14310 27298
rect 14362 27246 14420 27298
rect 14308 27244 14420 27246
rect 14308 27234 14364 27244
rect 14028 26994 14030 27046
rect 14082 26994 14084 27046
rect 14028 26982 14084 26994
rect 14476 26908 14532 28588
rect 14588 28420 14644 30034
rect 14924 29662 14980 31164
rect 15596 31050 15652 31612
rect 15596 30998 15598 31050
rect 15650 30998 15652 31050
rect 15596 30986 15652 30998
rect 15820 31220 15876 31230
rect 15820 31050 15876 31164
rect 15820 30998 15822 31050
rect 15874 30998 15876 31050
rect 15820 30986 15876 30998
rect 16044 31108 16100 31118
rect 16044 31050 16100 31052
rect 16044 30998 16046 31050
rect 16098 30998 16100 31050
rect 16044 30986 16100 30998
rect 16156 31029 16212 31041
rect 16156 30977 16158 31029
rect 16210 30977 16212 31029
rect 15036 30882 15092 30894
rect 15036 30830 15038 30882
rect 15090 30830 15092 30882
rect 15036 30182 15092 30830
rect 15316 30772 15372 30782
rect 15316 30770 16042 30772
rect 15316 30718 15318 30770
rect 15370 30718 16042 30770
rect 15316 30716 16042 30718
rect 15316 30706 15372 30716
rect 15484 30548 15540 30558
rect 15036 30130 15038 30182
rect 15090 30130 15092 30182
rect 15036 30118 15092 30130
rect 15148 30436 15204 30446
rect 14924 29650 15036 29662
rect 14924 29598 14982 29650
rect 15034 29598 15036 29650
rect 14924 29596 15036 29598
rect 14980 29586 15036 29596
rect 15148 29426 15204 30380
rect 15260 30154 15316 30166
rect 15260 30102 15262 30154
rect 15314 30102 15316 30154
rect 15260 30100 15316 30102
rect 15260 30034 15316 30044
rect 15372 30154 15428 30166
rect 15372 30102 15374 30154
rect 15426 30102 15428 30154
rect 15372 29988 15428 30102
rect 15372 29922 15428 29932
rect 15148 29374 15150 29426
rect 15202 29374 15204 29426
rect 15148 29362 15204 29374
rect 15484 29428 15540 30492
rect 15708 30210 15764 30222
rect 15708 30158 15710 30210
rect 15762 30158 15764 30210
rect 15708 29988 15764 30158
rect 15820 30210 15876 30222
rect 15820 30158 15822 30210
rect 15874 30158 15876 30210
rect 15820 30100 15876 30158
rect 15986 30210 16042 30716
rect 15986 30158 15988 30210
rect 16040 30158 16042 30210
rect 15986 30146 16042 30158
rect 15820 30034 15876 30044
rect 15708 29922 15764 29932
rect 16156 29764 16212 30977
rect 15652 29708 16212 29764
rect 15652 29650 15708 29708
rect 15652 29598 15654 29650
rect 15706 29598 15708 29650
rect 15652 29586 15708 29598
rect 15764 29428 15820 29438
rect 15484 29426 15820 29428
rect 15484 29374 15766 29426
rect 15818 29374 15820 29426
rect 15484 29372 15820 29374
rect 15764 29362 15820 29372
rect 15932 29428 15988 29438
rect 15932 29334 15988 29372
rect 15260 29204 15316 29214
rect 16268 29204 16324 32284
rect 16380 32004 16436 33180
rect 16380 31938 16436 31948
rect 16492 32452 16548 34636
rect 16772 34692 16828 34702
rect 16772 34598 16828 34636
rect 17332 34692 17388 34702
rect 17332 34690 17444 34692
rect 17332 34638 17334 34690
rect 17386 34638 17444 34690
rect 17332 34626 17444 34638
rect 16716 34244 16772 34254
rect 16716 34174 16772 34188
rect 16716 34122 16718 34174
rect 16770 34122 16772 34174
rect 16716 34110 16772 34122
rect 16940 34132 16996 34142
rect 16828 34020 16884 34030
rect 16604 34018 16884 34020
rect 16604 33966 16830 34018
rect 16882 33966 16884 34018
rect 16604 33964 16884 33966
rect 16604 33458 16660 33964
rect 16828 33954 16884 33964
rect 16940 33796 16996 34076
rect 16604 33406 16606 33458
rect 16658 33406 16660 33458
rect 16604 33394 16660 33406
rect 16828 33740 16996 33796
rect 17388 33796 17444 34626
rect 17500 34468 17556 34862
rect 17724 34916 17780 35646
rect 17836 35530 17892 36988
rect 17836 35478 17838 35530
rect 17890 35478 17892 35530
rect 17836 35466 17892 35478
rect 17724 34850 17780 34860
rect 17948 34804 18004 37324
rect 18620 37268 18676 37278
rect 18620 37174 18676 37212
rect 18844 36820 18900 38108
rect 19628 38108 20020 38164
rect 18956 38050 19012 38062
rect 18956 37998 18958 38050
rect 19010 37998 19012 38050
rect 18956 37044 19012 37998
rect 19292 38052 19348 38062
rect 19292 37958 19348 37996
rect 19124 37940 19180 37950
rect 19124 37490 19180 37884
rect 19124 37438 19126 37490
rect 19178 37438 19180 37490
rect 19124 37426 19180 37438
rect 19628 37268 19684 38108
rect 20300 38050 20356 38062
rect 20300 37998 20302 38050
rect 20354 37998 20356 38050
rect 20020 37940 20076 37950
rect 20300 37940 20356 37998
rect 20580 38052 20636 38062
rect 20748 38052 20804 38062
rect 20580 38050 20692 38052
rect 20580 37998 20582 38050
rect 20634 37998 20692 38050
rect 20580 37986 20692 37998
rect 20020 37938 20244 37940
rect 20020 37886 20022 37938
rect 20074 37886 20244 37938
rect 20020 37884 20244 37886
rect 20020 37874 20076 37884
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20076 37492 20132 37502
rect 19852 37268 19908 37278
rect 19628 37266 19908 37268
rect 19628 37214 19854 37266
rect 19906 37214 19908 37266
rect 19628 37212 19908 37214
rect 19852 37202 19908 37212
rect 20076 37098 20132 37436
rect 20188 37266 20244 37884
rect 20300 37874 20356 37884
rect 20412 37938 20468 37950
rect 20412 37886 20414 37938
rect 20466 37886 20468 37938
rect 20188 37214 20190 37266
rect 20242 37214 20244 37266
rect 20188 37202 20244 37214
rect 18956 36978 19012 36988
rect 19516 37042 19572 37054
rect 19516 36990 19518 37042
rect 19570 36990 19572 37042
rect 20076 37046 20078 37098
rect 20130 37046 20132 37098
rect 20076 37034 20132 37046
rect 18508 36764 18900 36820
rect 18396 35924 18452 35934
rect 18396 35830 18452 35868
rect 18172 34804 18228 34814
rect 17948 34748 18116 34804
rect 17668 34692 17724 34702
rect 17668 34690 18004 34692
rect 17668 34638 17670 34690
rect 17722 34638 18004 34690
rect 17668 34636 18004 34638
rect 17668 34626 17724 34636
rect 17500 34412 17668 34468
rect 17500 34244 17556 34254
rect 17500 34150 17556 34188
rect 17612 33908 17668 34412
rect 17743 34132 17799 34142
rect 17743 34038 17799 34076
rect 17612 33852 17780 33908
rect 16492 31892 16548 32396
rect 16604 31892 16660 31902
rect 16492 31890 16660 31892
rect 16492 31838 16606 31890
rect 16658 31838 16660 31890
rect 16492 31836 16660 31838
rect 16380 30322 16436 30334
rect 16380 30270 16382 30322
rect 16434 30270 16436 30322
rect 16380 29540 16436 30270
rect 16380 29474 16436 29484
rect 16492 29428 16548 31836
rect 16604 31826 16660 31836
rect 16716 31332 16772 31342
rect 16604 31220 16660 31230
rect 16604 31126 16660 31164
rect 16716 30548 16772 31276
rect 16828 30660 16884 33740
rect 17388 33730 17444 33740
rect 17724 33348 17780 33852
rect 17388 33124 17444 33134
rect 17052 32732 17332 32788
rect 16828 30594 16884 30604
rect 16940 30994 16996 31006
rect 16940 30942 16942 30994
rect 16994 30942 16996 30994
rect 16716 30482 16772 30492
rect 16940 30436 16996 30942
rect 16940 30370 16996 30380
rect 16940 30210 16996 30222
rect 16940 30158 16942 30210
rect 16994 30158 16996 30210
rect 16940 29876 16996 30158
rect 16940 29810 16996 29820
rect 16492 29362 16548 29372
rect 16828 29428 16884 29438
rect 16268 29148 16548 29204
rect 14812 28644 14868 28654
rect 15260 28642 15316 29148
rect 16268 28756 16324 28766
rect 14812 28550 14868 28588
rect 14980 28586 15036 28598
rect 14980 28534 14982 28586
rect 15034 28534 15036 28586
rect 15260 28590 15262 28642
rect 15314 28590 15316 28642
rect 15260 28578 15316 28590
rect 15932 28644 15988 28654
rect 15932 28550 15988 28588
rect 16268 28627 16324 28700
rect 16268 28575 16270 28627
rect 16322 28575 16324 28627
rect 16268 28563 16324 28575
rect 14980 28532 15036 28534
rect 14980 28476 15092 28532
rect 14588 28364 14980 28420
rect 14812 28196 14868 28206
rect 14812 27860 14868 28140
rect 14700 27858 14868 27860
rect 14700 27806 14814 27858
rect 14866 27806 14868 27858
rect 14700 27804 14868 27806
rect 14700 27300 14756 27804
rect 14812 27794 14868 27804
rect 14924 27858 14980 28364
rect 15036 28196 15092 28476
rect 15036 28130 15092 28140
rect 15148 28530 15204 28542
rect 15148 28478 15150 28530
rect 15202 28478 15204 28530
rect 15148 28084 15204 28478
rect 15540 28532 15596 28542
rect 15540 28530 15876 28532
rect 15540 28478 15542 28530
rect 15594 28478 15876 28530
rect 15540 28476 15876 28478
rect 15540 28466 15596 28476
rect 15820 28084 15876 28476
rect 16156 28474 16212 28486
rect 16156 28422 16158 28474
rect 16210 28422 16212 28474
rect 15148 28028 15316 28084
rect 15820 28028 15988 28084
rect 15036 27972 15092 27982
rect 15092 27916 15126 27972
rect 15036 27906 15126 27916
rect 14924 27806 14926 27858
rect 14978 27806 14980 27858
rect 15070 27896 15126 27906
rect 15070 27844 15072 27896
rect 15124 27844 15126 27896
rect 15070 27832 15126 27844
rect 14924 27794 14980 27806
rect 15260 27636 15316 28028
rect 15820 27858 15876 27870
rect 15820 27806 15822 27858
rect 15874 27806 15876 27858
rect 14700 27234 14756 27244
rect 14868 27580 15316 27636
rect 15484 27636 15540 27646
rect 15484 27634 15764 27636
rect 15484 27582 15486 27634
rect 15538 27582 15764 27634
rect 15484 27580 15764 27582
rect 14868 27298 14924 27580
rect 15484 27570 15540 27580
rect 14868 27246 14870 27298
rect 14922 27246 14924 27298
rect 14868 27234 14924 27246
rect 15148 27412 15204 27422
rect 15148 27074 15204 27356
rect 15596 27300 15652 27310
rect 15148 27022 15150 27074
rect 15202 27022 15204 27074
rect 15148 27010 15204 27022
rect 15372 27074 15428 27086
rect 15372 27022 15374 27074
rect 15426 27022 15428 27074
rect 14364 26852 14532 26908
rect 15372 26908 15428 27022
rect 15596 27074 15652 27244
rect 15596 27022 15598 27074
rect 15650 27022 15652 27074
rect 15596 27010 15652 27022
rect 15708 27074 15764 27580
rect 15820 27300 15876 27806
rect 15820 27234 15876 27244
rect 15932 27086 15988 28028
rect 16044 27860 16100 27870
rect 16044 27766 16100 27804
rect 15708 27022 15710 27074
rect 15762 27022 15764 27074
rect 15708 27010 15764 27022
rect 15876 27074 15988 27086
rect 15876 27022 15878 27074
rect 15930 27022 15988 27074
rect 15876 27020 15988 27022
rect 15876 27010 15932 27020
rect 16156 26908 16212 28422
rect 16324 27634 16380 27646
rect 16324 27582 16326 27634
rect 16378 27582 16380 27634
rect 16324 27412 16380 27582
rect 16324 27346 16380 27356
rect 15372 26852 16212 26908
rect 16268 27186 16324 27198
rect 16268 27134 16270 27186
rect 16322 27134 16324 27186
rect 16268 26964 16324 27134
rect 16268 26898 16324 26908
rect 16492 26908 16548 29148
rect 16828 28094 16884 29372
rect 16940 28868 16996 28878
rect 16940 28774 16996 28812
rect 16828 28082 16940 28094
rect 16828 28030 16886 28082
rect 16938 28030 16940 28082
rect 16828 28028 16940 28030
rect 16884 28018 16940 28028
rect 17052 27860 17108 32732
rect 17164 32564 17220 32574
rect 17164 31556 17220 32508
rect 17276 32450 17332 32732
rect 17388 32562 17444 33068
rect 17388 32510 17390 32562
rect 17442 32510 17444 32562
rect 17388 32498 17444 32510
rect 17724 33124 17780 33292
rect 17724 32562 17780 33068
rect 17724 32510 17726 32562
rect 17778 32510 17780 32562
rect 17724 32498 17780 32510
rect 17836 33796 17892 33806
rect 17276 32398 17278 32450
rect 17330 32398 17332 32450
rect 17276 32386 17332 32398
rect 17836 31948 17892 33740
rect 17948 33348 18004 34636
rect 18060 34468 18116 34748
rect 18172 34710 18228 34748
rect 18060 34402 18116 34412
rect 18508 34244 18564 36764
rect 19516 36484 19572 36990
rect 20412 36708 20468 37886
rect 20524 37716 20580 37726
rect 20524 37266 20580 37660
rect 20524 37214 20526 37266
rect 20578 37214 20580 37266
rect 20524 37202 20580 37214
rect 20636 37268 20692 37986
rect 20748 37958 20804 37996
rect 20636 37202 20692 37212
rect 20972 37940 21028 37950
rect 20804 36708 20860 36718
rect 20412 36652 20580 36708
rect 19516 36418 19572 36428
rect 19628 36482 19684 36494
rect 19628 36430 19630 36482
rect 19682 36430 19684 36482
rect 19180 35924 19236 35934
rect 19628 35924 19684 36430
rect 20412 36482 20468 36494
rect 20412 36430 20414 36482
rect 20466 36430 20468 36482
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19180 35922 19684 35924
rect 19180 35870 19182 35922
rect 19234 35870 19684 35922
rect 19180 35868 19684 35870
rect 19180 35858 19236 35868
rect 18844 35812 18900 35822
rect 18732 35698 18788 35710
rect 18732 35646 18734 35698
rect 18786 35646 18788 35698
rect 18732 35588 18788 35646
rect 18844 35698 18900 35756
rect 18844 35646 18846 35698
rect 18898 35646 18900 35698
rect 18844 35634 18900 35646
rect 20076 35698 20132 35710
rect 20076 35646 20078 35698
rect 20130 35646 20132 35698
rect 18732 35522 18788 35532
rect 20076 35140 20132 35646
rect 20300 35700 20356 35710
rect 20300 35606 20356 35644
rect 20076 35074 20132 35084
rect 20188 35530 20244 35542
rect 20188 35478 20190 35530
rect 20242 35478 20244 35530
rect 20076 34916 20132 34926
rect 19852 34914 20132 34916
rect 19852 34862 20078 34914
rect 20130 34862 20132 34914
rect 19852 34860 20132 34862
rect 19852 34692 19908 34860
rect 20076 34850 20132 34860
rect 19628 34636 19908 34692
rect 18508 34178 18564 34188
rect 18620 34580 18676 34590
rect 18620 34130 18676 34524
rect 19628 34356 19684 34636
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 20188 34356 20244 35478
rect 20412 34916 20468 36430
rect 20524 36148 20580 36652
rect 20804 36594 20860 36652
rect 20804 36542 20806 36594
rect 20858 36542 20860 36594
rect 20804 36530 20860 36542
rect 20524 36082 20580 36092
rect 20972 36484 21028 37884
rect 21084 37490 21140 39228
rect 21308 38834 21364 39228
rect 21308 38782 21310 38834
rect 21362 38782 21364 38834
rect 21308 38770 21364 38782
rect 21420 38668 21476 41132
rect 21532 40964 21588 42700
rect 21644 42754 21700 44044
rect 21980 43706 22036 43718
rect 21868 43652 21924 43662
rect 21868 43594 21924 43596
rect 21644 42702 21646 42754
rect 21698 42702 21700 42754
rect 21644 42690 21700 42702
rect 21756 43540 21812 43550
rect 21868 43542 21870 43594
rect 21922 43542 21924 43594
rect 21868 43530 21924 43542
rect 21980 43654 21982 43706
rect 22034 43654 22036 43706
rect 21644 42196 21700 42206
rect 21644 41970 21700 42140
rect 21644 41918 21646 41970
rect 21698 41918 21700 41970
rect 21644 41906 21700 41918
rect 21756 41300 21812 43484
rect 21980 41970 22036 43654
rect 22204 43652 22260 43662
rect 22092 43540 22148 43550
rect 22092 43446 22148 43484
rect 22204 42094 22260 43596
rect 22764 43650 22820 44716
rect 23212 44716 23492 44772
rect 23660 45890 23716 45902
rect 23660 45838 23662 45890
rect 23714 45838 23716 45890
rect 22764 43598 22766 43650
rect 22818 43598 22820 43650
rect 22764 43586 22820 43598
rect 23007 43652 23063 43662
rect 23007 43594 23063 43596
rect 23007 43542 23009 43594
rect 23061 43542 23063 43594
rect 23007 43530 23063 43542
rect 23212 43092 23268 44716
rect 23436 44324 23492 44334
rect 23436 44230 23492 44268
rect 23660 44324 23716 45838
rect 23772 44436 23828 46508
rect 23884 45108 23940 47180
rect 24556 47236 24612 47246
rect 24556 46674 24612 47180
rect 24668 47124 24724 47362
rect 24668 47058 24724 47068
rect 24780 47290 24836 47302
rect 24780 47238 24782 47290
rect 24834 47238 24836 47290
rect 24556 46622 24558 46674
rect 24610 46622 24612 46674
rect 24556 46610 24612 46622
rect 24780 46340 24836 47238
rect 25340 47124 25396 47134
rect 25340 46786 25396 47068
rect 26348 47012 26404 47406
rect 25340 46734 25342 46786
rect 25394 46734 25396 46786
rect 25340 46722 25396 46734
rect 25788 46956 26404 47012
rect 25583 46705 25639 46717
rect 25583 46653 25585 46705
rect 25637 46676 25639 46705
rect 25788 46676 25844 46956
rect 25637 46653 25844 46676
rect 25583 46620 25844 46653
rect 26460 46676 26516 47628
rect 30660 47570 30716 47966
rect 30660 47518 30662 47570
rect 30714 47518 30716 47570
rect 30660 47506 30716 47518
rect 31836 48018 31892 50200
rect 31836 47966 31838 48018
rect 31890 47966 31892 48018
rect 26628 47460 26684 47470
rect 26628 47366 26684 47404
rect 28364 47458 28420 47470
rect 28364 47406 28366 47458
rect 28418 47406 28420 47458
rect 27580 46676 27636 46686
rect 26460 46674 26740 46676
rect 26460 46622 26462 46674
rect 26514 46622 26740 46674
rect 26460 46620 26740 46622
rect 24556 46284 24836 46340
rect 24444 46004 24500 46014
rect 24556 46004 24612 46284
rect 24444 46002 24612 46004
rect 24444 45950 24446 46002
rect 24498 45950 24612 46002
rect 24444 45948 24612 45950
rect 24444 45938 24500 45948
rect 25564 45121 25620 45133
rect 23884 45042 23940 45052
rect 25228 45108 25284 45118
rect 25228 45014 25284 45052
rect 25564 45069 25566 45121
rect 25618 45069 25620 45121
rect 23772 44370 23828 44380
rect 24220 44996 24276 45006
rect 24220 44994 25060 44996
rect 24220 44942 24222 44994
rect 24274 44942 25060 44994
rect 24220 44940 25060 44942
rect 23660 44258 23716 44268
rect 24220 43708 24276 44940
rect 24780 44436 24836 44446
rect 24780 44342 24836 44380
rect 23884 43652 24276 43708
rect 24444 44322 24500 44334
rect 24444 44270 24446 44322
rect 24498 44270 24500 44322
rect 25004 44322 25060 44940
rect 25564 44436 25620 45069
rect 25676 44994 25732 46620
rect 26460 46610 26516 46620
rect 26348 45892 26404 45902
rect 26348 45798 26404 45836
rect 26684 45892 26740 46620
rect 27580 46582 27636 46620
rect 28364 46676 28420 47406
rect 29240 47460 29296 47470
rect 29240 47366 29296 47404
rect 30492 47460 30548 47470
rect 29484 47348 29540 47358
rect 29372 47346 29540 47348
rect 29372 47294 29486 47346
rect 29538 47294 29540 47346
rect 29372 47292 29540 47294
rect 28364 46610 28420 46620
rect 29260 47236 29316 47246
rect 26684 45826 26740 45836
rect 27692 46060 28420 46116
rect 27692 45890 27748 46060
rect 27692 45838 27694 45890
rect 27746 45838 27748 45890
rect 27692 45826 27748 45838
rect 27804 45892 27860 45902
rect 27804 45798 27860 45836
rect 26684 45668 26740 45678
rect 25676 44942 25678 44994
rect 25730 44942 25732 44994
rect 25676 44930 25732 44942
rect 25900 45106 25956 45118
rect 25900 45054 25902 45106
rect 25954 45054 25956 45106
rect 25564 44370 25620 44380
rect 23884 43538 23940 43652
rect 24444 43606 24500 44270
rect 24388 43596 24500 43606
rect 24332 43594 24500 43596
rect 23884 43486 23886 43538
rect 23938 43486 23940 43538
rect 23884 43474 23940 43486
rect 24220 43540 24276 43550
rect 24220 43426 24276 43484
rect 24220 43374 24222 43426
rect 24274 43374 24276 43426
rect 24220 43362 24276 43374
rect 24332 43542 24390 43594
rect 24442 43542 24500 43594
rect 24668 44266 24724 44278
rect 24668 44214 24670 44266
rect 24722 44214 24724 44266
rect 24332 43540 24500 43542
rect 24556 43540 24612 43550
rect 24668 43540 24724 44214
rect 25004 44270 25006 44322
rect 25058 44270 25060 44322
rect 25004 43708 25060 44270
rect 24332 43530 24444 43540
rect 24556 43538 24724 43540
rect 23212 43036 23604 43092
rect 22428 42754 22484 42766
rect 22428 42702 22430 42754
rect 22482 42702 22484 42754
rect 22428 42196 22484 42702
rect 23548 42532 23604 43036
rect 24332 42868 24388 43530
rect 22428 42130 22484 42140
rect 23100 42476 23604 42532
rect 24220 42812 24388 42868
rect 24556 43486 24558 43538
rect 24610 43486 24724 43538
rect 24556 43484 24724 43486
rect 24780 43652 25060 43708
rect 25228 44324 25284 44334
rect 25116 43652 25172 43662
rect 22204 42082 22316 42094
rect 22204 42030 22262 42082
rect 22314 42030 22316 42082
rect 22204 42028 22316 42030
rect 22260 42018 22316 42028
rect 21980 41918 21982 41970
rect 22034 41918 22036 41970
rect 21980 41906 22036 41918
rect 22540 41970 22596 41982
rect 22540 41918 22542 41970
rect 22594 41918 22596 41970
rect 22540 41860 22596 41918
rect 22764 41972 22820 41982
rect 22764 41878 22820 41916
rect 22540 41794 22596 41804
rect 21756 41234 21812 41244
rect 21868 41188 21924 41198
rect 22876 41188 22932 41198
rect 21868 41094 21924 41132
rect 22540 41186 22932 41188
rect 22540 41134 22878 41186
rect 22930 41134 22932 41186
rect 22540 41132 22932 41134
rect 22372 40964 22428 40974
rect 21532 39592 21588 40908
rect 22316 40962 22428 40964
rect 22316 40910 22374 40962
rect 22426 40910 22428 40962
rect 22316 40898 22428 40910
rect 22316 40740 22372 40898
rect 22316 40674 22372 40684
rect 22428 40628 22484 40638
rect 21980 40068 22036 40078
rect 22428 40068 22484 40572
rect 21644 39592 21700 39602
rect 21532 39590 21812 39592
rect 21532 39538 21646 39590
rect 21698 39538 21812 39590
rect 21532 39536 21812 39538
rect 21644 39526 21700 39536
rect 21420 38612 21588 38668
rect 21420 38162 21476 38174
rect 21420 38110 21422 38162
rect 21474 38110 21476 38162
rect 21308 38052 21364 38062
rect 21308 37958 21364 37996
rect 21420 37716 21476 38110
rect 21420 37650 21476 37660
rect 21084 37438 21086 37490
rect 21138 37438 21140 37490
rect 21084 37426 21140 37438
rect 21420 37268 21476 37278
rect 21420 37174 21476 37212
rect 21532 37266 21588 38612
rect 21644 37994 21700 38006
rect 21644 37942 21646 37994
rect 21698 37942 21700 37994
rect 21644 37380 21700 37942
rect 21644 37314 21700 37324
rect 21532 37214 21534 37266
rect 21586 37214 21588 37266
rect 21532 37202 21588 37214
rect 21756 36606 21812 39536
rect 21700 36594 21812 36606
rect 21700 36542 21702 36594
rect 21754 36542 21812 36594
rect 21700 36530 21812 36542
rect 20804 35700 20860 35710
rect 20972 35700 21028 36428
rect 21196 36148 21252 36158
rect 21196 35810 21252 36092
rect 21196 35758 21198 35810
rect 21250 35758 21252 35810
rect 21196 35746 21252 35758
rect 21084 35700 21140 35710
rect 20972 35698 21140 35700
rect 20972 35646 21086 35698
rect 21138 35646 21140 35698
rect 21532 35698 21588 35710
rect 20972 35644 21140 35646
rect 20804 35606 20860 35644
rect 21084 35634 21140 35644
rect 21364 35642 21420 35654
rect 21364 35590 21366 35642
rect 21418 35590 21420 35642
rect 21364 35364 21420 35590
rect 21084 35308 21420 35364
rect 21532 35646 21534 35698
rect 21586 35646 21588 35698
rect 20972 35140 21028 35150
rect 20860 34916 20916 34926
rect 20412 34914 20916 34916
rect 20412 34862 20862 34914
rect 20914 34862 20916 34914
rect 20412 34860 20916 34862
rect 19628 34300 19908 34356
rect 19852 34298 19908 34300
rect 19852 34246 19854 34298
rect 19906 34246 19908 34298
rect 19852 34234 19908 34246
rect 20076 34300 20244 34356
rect 20076 34174 20132 34300
rect 18620 34078 18622 34130
rect 18674 34078 18676 34130
rect 18620 34066 18676 34078
rect 19012 34132 19068 34142
rect 19012 34038 19068 34076
rect 19292 34130 19348 34142
rect 19292 34078 19294 34130
rect 19346 34078 19348 34130
rect 17948 33282 18004 33292
rect 18172 33684 18228 33694
rect 17612 31892 18116 31948
rect 17612 31750 17668 31892
rect 17612 31698 17614 31750
rect 17666 31698 17668 31750
rect 17612 31686 17668 31698
rect 17836 31778 17892 31790
rect 17836 31726 17838 31778
rect 17890 31726 17892 31778
rect 17836 31556 17892 31726
rect 17164 31500 17892 31556
rect 17164 29428 17220 31500
rect 17388 31332 17444 31342
rect 17388 30994 17444 31276
rect 17388 30942 17390 30994
rect 17442 30942 17444 30994
rect 17388 30930 17444 30942
rect 17276 30660 17332 30670
rect 17276 30183 17332 30604
rect 17276 30131 17278 30183
rect 17330 30131 17332 30183
rect 17276 30119 17332 30131
rect 17388 30548 17444 30558
rect 18060 30548 18116 31892
rect 18172 31220 18228 33628
rect 18508 33460 18564 33470
rect 19292 33460 19348 34078
rect 19516 34130 19572 34142
rect 19516 34078 19518 34130
rect 19570 34078 19572 34130
rect 18508 33366 18564 33404
rect 19068 33404 19348 33460
rect 19404 33572 19460 33582
rect 18284 32562 18340 32574
rect 18284 32510 18286 32562
rect 18338 32510 18340 32562
rect 18284 31780 18340 32510
rect 18284 31714 18340 31724
rect 18508 32564 18564 32574
rect 19068 32564 19124 33404
rect 19404 33346 19460 33516
rect 19404 33294 19406 33346
rect 19458 33294 19460 33346
rect 19404 33282 19460 33294
rect 19236 33236 19292 33246
rect 19236 33178 19292 33180
rect 19236 33126 19238 33178
rect 19290 33126 19292 33178
rect 19236 33114 19292 33126
rect 19516 32676 19572 34078
rect 19740 34130 19796 34142
rect 19740 34078 19742 34130
rect 19794 34078 19796 34130
rect 20076 34122 20078 34174
rect 20130 34122 20132 34174
rect 20076 34110 20132 34122
rect 20636 34132 20692 34142
rect 19740 33908 19796 34078
rect 19740 33842 19796 33852
rect 20188 33460 20244 33470
rect 19740 33348 19796 33358
rect 19628 33290 19684 33302
rect 19628 33238 19630 33290
rect 19682 33238 19684 33290
rect 20188 33318 20244 33404
rect 19740 33266 19742 33292
rect 19794 33266 19796 33292
rect 19740 33254 19796 33266
rect 19964 33290 20020 33302
rect 19628 33012 19684 33238
rect 19964 33238 19966 33290
rect 20018 33238 20020 33290
rect 19964 33236 20020 33238
rect 19964 33170 20020 33180
rect 20188 33266 20190 33318
rect 20242 33266 20244 33318
rect 20636 33348 20692 34076
rect 20860 33908 20916 34860
rect 20972 34020 21028 35084
rect 20972 33926 21028 33964
rect 21084 34169 21140 35308
rect 21084 34117 21086 34169
rect 21138 34117 21140 34169
rect 20860 33842 20916 33852
rect 20636 33292 21028 33348
rect 19628 32946 19684 32956
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19404 32620 19572 32676
rect 19404 32601 19460 32620
rect 19180 32564 19236 32574
rect 19068 32562 19236 32564
rect 19068 32510 19182 32562
rect 19234 32510 19236 32562
rect 19068 32508 19236 32510
rect 18172 31164 18340 31220
rect 18284 31108 18340 31164
rect 18264 31050 18340 31108
rect 18264 30998 18266 31050
rect 18318 30998 18340 31050
rect 18264 30986 18340 30998
rect 18508 30996 18564 32508
rect 19180 32116 19236 32508
rect 19404 32564 19406 32601
rect 19458 32564 19460 32601
rect 19404 32498 19460 32508
rect 19852 32564 19908 32574
rect 20188 32564 20244 33266
rect 19852 32562 20244 32564
rect 19852 32510 19854 32562
rect 19906 32510 20190 32562
rect 20242 32510 20244 32562
rect 19852 32508 20244 32510
rect 19852 32498 19908 32508
rect 20188 32498 20244 32508
rect 20300 33236 20356 33246
rect 20468 33236 20524 33246
rect 20300 32562 20356 33180
rect 20300 32510 20302 32562
rect 20354 32510 20356 32562
rect 20300 32498 20356 32510
rect 20412 33234 20524 33236
rect 20412 33182 20470 33234
rect 20522 33182 20524 33234
rect 20412 33170 20524 33182
rect 19516 32450 19572 32462
rect 19516 32398 19518 32450
rect 19570 32398 19572 32450
rect 19516 32340 19572 32398
rect 20412 32340 20468 33170
rect 20860 32562 20916 32574
rect 20860 32510 20862 32562
rect 20914 32510 20916 32562
rect 19516 32274 19572 32284
rect 20188 32284 20468 32340
rect 20580 32340 20636 32350
rect 20580 32338 20692 32340
rect 20580 32286 20582 32338
rect 20634 32286 20692 32338
rect 19180 32050 19236 32060
rect 18620 31778 18676 31790
rect 18620 31726 18622 31778
rect 18674 31726 18676 31778
rect 18620 31220 18676 31726
rect 20188 31556 20244 32284
rect 20580 32274 20692 32286
rect 20524 32004 20580 32014
rect 20524 31892 20580 31948
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 18620 31154 18676 31164
rect 19124 31162 19180 31174
rect 17276 29428 17332 29438
rect 17164 29426 17332 29428
rect 17164 29374 17278 29426
rect 17330 29374 17332 29426
rect 17164 29372 17332 29374
rect 17276 29362 17332 29372
rect 17388 28868 17444 30492
rect 17948 30492 18116 30548
rect 17836 30324 17892 30334
rect 17612 30212 17668 30222
rect 17612 30118 17668 30156
rect 17724 30042 17780 30054
rect 17724 29990 17726 30042
rect 17778 29990 17780 30042
rect 17052 27794 17108 27804
rect 17164 28812 17444 28868
rect 17500 29876 17556 29886
rect 17164 27636 17220 28812
rect 17052 27580 17220 27636
rect 17276 28644 17332 28654
rect 17388 28644 17444 28654
rect 17276 28642 17444 28644
rect 17276 28590 17278 28642
rect 17330 28590 17390 28642
rect 17442 28590 17444 28642
rect 17276 28588 17444 28590
rect 16492 26852 16660 26908
rect 13916 26460 14308 26516
rect 13692 26282 13748 26294
rect 13804 26318 13860 26330
rect 13132 25452 13300 25508
rect 13020 25340 13188 25396
rect 12852 25284 12908 25294
rect 12852 25190 12908 25228
rect 12572 24882 12628 24892
rect 12236 23874 12292 23884
rect 12348 24388 12404 24398
rect 12348 23910 12404 24332
rect 12348 23858 12350 23910
rect 12402 23858 12404 23910
rect 12348 23846 12404 23858
rect 12460 24052 12516 24062
rect 11732 23828 11788 23838
rect 11732 23734 11788 23772
rect 12460 23716 12516 23996
rect 12572 23940 12628 23950
rect 12572 23858 12574 23884
rect 12626 23858 12628 23884
rect 12572 23846 12628 23858
rect 12796 23940 12852 23950
rect 12796 23858 12798 23884
rect 12850 23858 12852 23884
rect 12796 23846 12852 23858
rect 12908 23882 12964 23894
rect 12908 23830 12910 23882
rect 12962 23830 12964 23882
rect 12908 23828 12964 23830
rect 12460 23660 12628 23716
rect 11396 23268 11452 23278
rect 11396 23174 11452 23212
rect 12572 23210 12628 23660
rect 11956 23189 12012 23201
rect 11956 23156 11958 23189
rect 11900 23137 11958 23156
rect 12010 23137 12012 23189
rect 11900 23100 12012 23137
rect 12236 23182 12292 23194
rect 12236 23130 12238 23182
rect 12290 23130 12292 23182
rect 11732 22932 11788 22942
rect 11732 22838 11788 22876
rect 11900 22708 11956 23100
rect 11788 22652 11956 22708
rect 11228 22306 11284 22316
rect 11564 22372 11620 22382
rect 11564 22278 11620 22316
rect 11396 21812 11452 21822
rect 11396 21718 11452 21756
rect 11788 21700 11844 22652
rect 11900 22372 11956 22382
rect 11900 22036 11956 22316
rect 12068 22260 12124 22270
rect 12068 22166 12124 22204
rect 12236 22148 12292 23130
rect 12460 23182 12516 23194
rect 12460 23130 12462 23182
rect 12514 23130 12516 23182
rect 12572 23158 12574 23210
rect 12626 23158 12628 23210
rect 12572 23146 12628 23158
rect 12460 22484 12516 23130
rect 12460 22418 12516 22428
rect 12348 22372 12404 22382
rect 12796 22372 12852 22382
rect 12348 22290 12350 22316
rect 12402 22290 12404 22316
rect 12348 22278 12404 22290
rect 12572 22314 12628 22326
rect 12236 22082 12292 22092
rect 12572 22262 12574 22314
rect 12626 22262 12628 22314
rect 12796 22290 12798 22316
rect 12850 22290 12852 22316
rect 12796 22278 12852 22290
rect 12908 22335 12964 23772
rect 13132 23828 13188 25340
rect 13244 25284 13300 25452
rect 13356 25284 13412 25294
rect 13244 25228 13356 25284
rect 13244 25060 13300 25070
rect 13244 23940 13300 25004
rect 13244 23874 13300 23884
rect 13132 23762 13188 23772
rect 13356 23492 13412 25228
rect 13468 24388 13524 26238
rect 13804 26266 13806 26318
rect 13858 26266 13860 26318
rect 13804 25060 13860 26266
rect 13916 25618 13972 26460
rect 14084 26325 14140 26337
rect 14084 26273 14086 26325
rect 14138 26292 14140 26325
rect 14252 26318 14308 26460
rect 14138 26273 14196 26292
rect 14084 26236 14196 26273
rect 14252 26266 14254 26318
rect 14306 26266 14308 26318
rect 14252 26254 14308 26266
rect 13916 25566 13918 25618
rect 13970 25566 13972 25618
rect 13916 25554 13972 25566
rect 13804 24994 13860 25004
rect 14140 25172 14196 26236
rect 14364 26180 14420 26852
rect 15764 26516 15820 26526
rect 14532 26292 14588 26302
rect 14812 26292 14868 26302
rect 14532 26290 14868 26292
rect 14532 26238 14534 26290
rect 14586 26238 14814 26290
rect 14866 26238 14868 26290
rect 14532 26236 14868 26238
rect 14532 26226 14588 26236
rect 14812 26226 14868 26236
rect 14364 26114 14420 26124
rect 15764 26180 15820 26460
rect 16604 26516 16660 26852
rect 16604 26450 16660 26460
rect 16660 26180 16716 26190
rect 15764 26178 15988 26180
rect 15764 26126 15766 26178
rect 15818 26126 15988 26178
rect 15764 26124 15988 26126
rect 15764 26114 15820 26124
rect 15148 26068 15204 26078
rect 15148 26066 15652 26068
rect 15148 26014 15150 26066
rect 15202 26014 15652 26066
rect 15148 26012 15652 26014
rect 15148 26002 15204 26012
rect 15596 25732 15652 26012
rect 15596 25676 15876 25732
rect 15820 25618 15876 25676
rect 15820 25566 15822 25618
rect 15874 25566 15876 25618
rect 15820 25554 15876 25566
rect 13468 24322 13524 24332
rect 13916 24610 13972 24622
rect 13916 24558 13918 24610
rect 13970 24558 13972 24610
rect 13916 24388 13972 24558
rect 14140 24612 14196 25116
rect 15260 25060 15316 25070
rect 15260 24946 15316 25004
rect 15260 24894 15262 24946
rect 15314 24894 15316 24946
rect 15260 24882 15316 24894
rect 14476 24836 14532 24846
rect 14476 24766 14532 24780
rect 14476 24714 14478 24766
rect 14530 24714 14532 24766
rect 15596 24836 15652 24846
rect 14476 24702 14532 24714
rect 14700 24724 14756 24734
rect 14364 24612 14420 24622
rect 14140 24610 14420 24612
rect 14140 24558 14366 24610
rect 14418 24558 14420 24610
rect 14140 24556 14420 24558
rect 14364 24546 14420 24556
rect 13916 24322 13972 24332
rect 13916 24164 13972 24174
rect 13580 24052 13636 24062
rect 13580 23958 13636 23996
rect 13356 23426 13412 23436
rect 13916 23938 13972 24108
rect 14700 24062 14756 24668
rect 15596 24722 15652 24780
rect 15596 24670 15598 24722
rect 15650 24670 15652 24722
rect 15596 24062 15652 24670
rect 15932 24500 15988 26124
rect 16492 26124 16660 26180
rect 16492 24722 16548 26124
rect 16660 26086 16716 26124
rect 16492 24670 16494 24722
rect 16546 24670 16548 24722
rect 16492 24658 16548 24670
rect 16604 25508 16660 25518
rect 16940 25508 16996 25518
rect 16604 25506 16996 25508
rect 16604 25454 16606 25506
rect 16658 25454 16942 25506
rect 16994 25454 16996 25506
rect 16604 25452 16996 25454
rect 16604 24722 16660 25452
rect 16940 25442 16996 25452
rect 17052 25172 17108 27580
rect 17164 27186 17220 27198
rect 17164 27134 17166 27186
rect 17218 27134 17220 27186
rect 17164 26908 17220 27134
rect 17276 26908 17332 28588
rect 17388 28578 17444 28588
rect 17500 27858 17556 29820
rect 17724 28644 17780 29990
rect 17724 28578 17780 28588
rect 17724 28420 17780 28430
rect 17836 28420 17892 30268
rect 17724 28418 17892 28420
rect 17724 28366 17726 28418
rect 17778 28366 17892 28418
rect 17724 28364 17892 28366
rect 17724 28354 17780 28364
rect 17836 28084 17892 28094
rect 17500 27806 17502 27858
rect 17554 27806 17556 27858
rect 17164 26852 17332 26908
rect 17052 25106 17108 25116
rect 17164 26516 17220 26526
rect 16604 24670 16606 24722
rect 16658 24670 16660 24722
rect 16156 24500 16212 24510
rect 15932 24498 16212 24500
rect 15932 24446 16158 24498
rect 16210 24446 16212 24498
rect 15932 24444 16212 24446
rect 14644 24050 14756 24062
rect 14644 23998 14646 24050
rect 14698 23998 14756 24050
rect 14644 23986 14756 23998
rect 15092 24052 15148 24062
rect 15540 24052 15652 24062
rect 15092 24050 15652 24052
rect 15092 23998 15094 24050
rect 15146 23998 15542 24050
rect 15594 23998 15652 24050
rect 15092 23996 15652 23998
rect 15988 24276 16044 24286
rect 15988 24050 16044 24220
rect 15988 23998 15990 24050
rect 16042 23998 16044 24050
rect 15092 23986 15148 23996
rect 15540 23986 15596 23996
rect 13916 23886 13918 23938
rect 13970 23886 13972 23938
rect 13188 23380 13244 23390
rect 13188 23286 13244 23324
rect 13916 23380 13972 23886
rect 13916 23314 13972 23324
rect 14252 23492 14308 23502
rect 12908 22283 12910 22335
rect 12962 22283 12964 22335
rect 12572 22148 12628 22262
rect 12572 22082 12628 22092
rect 12348 22036 12404 22046
rect 11900 21980 12068 22036
rect 10892 21534 10894 21586
rect 10946 21534 10948 21586
rect 10892 21522 10948 21534
rect 11676 21644 11844 21700
rect 10556 21364 10612 21374
rect 10108 21362 10612 21364
rect 10108 21310 10558 21362
rect 10610 21310 10612 21362
rect 10108 21308 10612 21310
rect 10108 20914 10164 21308
rect 10556 21298 10612 21308
rect 11676 21252 11732 21644
rect 12012 21586 12068 21980
rect 12012 21534 12014 21586
rect 12066 21534 12068 21586
rect 12012 21522 12068 21534
rect 11844 21476 11900 21486
rect 11844 21382 11900 21420
rect 12348 21476 12404 21980
rect 12908 21812 12964 22283
rect 12908 21746 12964 21756
rect 13020 23156 13076 23166
rect 12348 21410 12404 21420
rect 12460 21586 12516 21598
rect 12460 21534 12462 21586
rect 12514 21534 12516 21586
rect 12180 21364 12236 21374
rect 12180 21362 12292 21364
rect 12180 21310 12182 21362
rect 12234 21310 12292 21362
rect 12180 21298 12292 21310
rect 11676 21196 11956 21252
rect 10108 20862 10110 20914
rect 10162 20862 10164 20914
rect 10108 20850 10164 20862
rect 9660 20804 9716 20814
rect 9660 19234 9716 20748
rect 11900 20692 11956 21196
rect 12012 20692 12068 20702
rect 11900 20690 12068 20692
rect 11900 20638 12014 20690
rect 12066 20638 12068 20690
rect 11900 20636 12068 20638
rect 11508 20047 11564 20059
rect 11508 19995 11510 20047
rect 11562 20020 11564 20047
rect 11562 19995 11620 20020
rect 11508 19964 11620 19995
rect 11340 19908 11396 19918
rect 10444 19906 11396 19908
rect 10444 19854 11342 19906
rect 11394 19854 11396 19906
rect 10444 19852 11396 19854
rect 10444 19346 10500 19852
rect 11340 19842 11396 19852
rect 10444 19294 10446 19346
rect 10498 19294 10500 19346
rect 10444 19282 10500 19294
rect 9660 19182 9662 19234
rect 9714 19182 9716 19234
rect 9660 19170 9716 19182
rect 11564 18564 11620 19964
rect 11788 20018 11844 20030
rect 11788 19966 11790 20018
rect 11842 19966 11844 20018
rect 11676 18564 11732 18574
rect 11564 18562 11732 18564
rect 11564 18510 11678 18562
rect 11730 18510 11732 18562
rect 11564 18508 11732 18510
rect 11676 18498 11732 18508
rect 11564 17780 11620 17790
rect 9548 17602 9604 17612
rect 9940 17668 9996 17678
rect 9940 17574 9996 17612
rect 11228 17666 11284 17678
rect 11228 17614 11230 17666
rect 11282 17614 11284 17666
rect 9324 17042 9380 17052
rect 11228 17108 11284 17614
rect 11452 17668 11508 17691
rect 11564 17686 11620 17724
rect 11788 17668 11844 19966
rect 11900 19236 11956 20636
rect 12012 20626 12068 20636
rect 12236 20132 12292 21298
rect 12348 20802 12404 20814
rect 12348 20750 12350 20802
rect 12402 20750 12404 20802
rect 12348 20244 12404 20750
rect 12460 20804 12516 21534
rect 12460 20738 12516 20748
rect 12572 20916 12628 20926
rect 12572 20802 12628 20860
rect 12572 20750 12574 20802
rect 12626 20750 12628 20802
rect 12572 20738 12628 20750
rect 12852 20692 12908 20702
rect 12684 20690 12908 20692
rect 12684 20638 12854 20690
rect 12906 20638 12908 20690
rect 12684 20636 12908 20638
rect 12572 20244 12628 20254
rect 12348 20188 12516 20244
rect 12068 20074 12124 20086
rect 12236 20076 12348 20132
rect 12068 20022 12070 20074
rect 12122 20022 12124 20074
rect 12068 19572 12124 20022
rect 12292 20074 12348 20076
rect 12292 20022 12294 20074
rect 12346 20022 12348 20074
rect 12292 20010 12348 20022
rect 12460 19572 12516 20188
rect 12572 20074 12628 20188
rect 12572 20022 12574 20074
rect 12626 20022 12628 20074
rect 12684 20132 12740 20636
rect 12852 20626 12908 20636
rect 12684 20066 12740 20076
rect 12572 20010 12628 20022
rect 13020 20020 13076 23100
rect 13356 23156 13412 23166
rect 13356 23154 13580 23156
rect 13356 23102 13358 23154
rect 13410 23102 13580 23154
rect 13356 23100 13580 23102
rect 13356 23090 13412 23100
rect 13524 22594 13580 23100
rect 13524 22542 13526 22594
rect 13578 22542 13580 22594
rect 13524 22530 13580 22542
rect 13692 22930 13748 22942
rect 13692 22878 13694 22930
rect 13746 22878 13748 22930
rect 13692 22260 13748 22878
rect 14252 22932 14308 23436
rect 14588 23268 14644 23278
rect 14588 23154 14644 23212
rect 14588 23102 14590 23154
rect 14642 23102 14644 23154
rect 14252 22930 14420 22932
rect 14252 22878 14254 22930
rect 14306 22878 14420 22930
rect 14252 22876 14420 22878
rect 14252 22866 14308 22876
rect 14252 22372 14308 22382
rect 13244 22204 13748 22260
rect 13804 22314 13860 22326
rect 13804 22262 13806 22314
rect 13858 22262 13860 22314
rect 13244 21586 13300 22204
rect 13804 21924 13860 22262
rect 14028 22314 14084 22326
rect 14028 22262 14030 22314
rect 14082 22262 14084 22314
rect 14252 22290 14254 22316
rect 14306 22290 14308 22316
rect 14252 22278 14308 22290
rect 14364 22314 14420 22876
rect 14588 22820 14644 23102
rect 14700 22932 14756 23986
rect 15988 23828 16044 23998
rect 15988 23762 16044 23772
rect 15260 23154 15316 23166
rect 15260 23102 15262 23154
rect 15314 23102 15316 23154
rect 15092 23044 15148 23054
rect 15260 23044 15316 23102
rect 15092 23042 15316 23044
rect 15092 22990 15094 23042
rect 15146 22990 15316 23042
rect 15092 22988 15316 22990
rect 15092 22978 15148 22988
rect 14700 22866 14756 22876
rect 14588 22754 14644 22764
rect 15260 22708 15316 22988
rect 15260 22642 15316 22652
rect 15484 23156 15540 23166
rect 14028 22148 14084 22262
rect 14028 22082 14084 22092
rect 14364 22262 14366 22314
rect 14418 22262 14420 22314
rect 14364 22036 14420 22262
rect 14364 21970 14420 21980
rect 14924 22370 14980 22382
rect 14924 22318 14926 22370
rect 14978 22318 14980 22370
rect 13804 21858 13860 21868
rect 13244 21534 13246 21586
rect 13298 21534 13300 21586
rect 13244 21522 13300 21534
rect 14588 21700 14644 21710
rect 14028 20916 14084 20926
rect 13356 20804 13412 20814
rect 13356 20710 13412 20748
rect 13468 20132 13524 20142
rect 13468 20045 13524 20076
rect 13468 20020 13470 20045
rect 12068 19516 12404 19572
rect 12348 19348 12404 19516
rect 12460 19506 12516 19516
rect 12908 19993 13470 20020
rect 13522 19993 13524 20045
rect 12908 19964 13524 19993
rect 12908 19358 12964 19964
rect 13020 19796 13076 19806
rect 13020 19702 13076 19740
rect 13916 19572 13972 19582
rect 12348 19346 12852 19348
rect 12348 19294 12350 19346
rect 12402 19294 12852 19346
rect 12348 19292 12852 19294
rect 12908 19346 13020 19358
rect 12908 19294 12966 19346
rect 13018 19294 13020 19346
rect 12908 19292 13020 19294
rect 12348 19282 12404 19292
rect 11900 19170 11956 19180
rect 11919 18450 11975 18462
rect 11919 18398 11921 18450
rect 11973 18398 11975 18450
rect 11919 18004 11975 18398
rect 12796 18452 12852 19292
rect 12964 19282 13020 19292
rect 13356 19236 13412 19246
rect 13356 19142 13412 19180
rect 13916 19234 13972 19516
rect 13916 19182 13918 19234
rect 13970 19182 13972 19234
rect 13748 19124 13804 19134
rect 13524 19012 13580 19022
rect 13524 18462 13580 18956
rect 13356 18452 13412 18462
rect 12796 18450 13188 18452
rect 12796 18398 12798 18450
rect 12850 18398 13188 18450
rect 12796 18396 13188 18398
rect 12796 18386 12852 18396
rect 11919 17938 11975 17948
rect 12796 18116 12852 18126
rect 12236 17780 12292 17790
rect 11900 17668 11956 17678
rect 11788 17666 11956 17668
rect 11788 17614 11902 17666
rect 11954 17614 11956 17666
rect 11788 17612 11956 17614
rect 11452 17599 11454 17612
rect 11506 17599 11508 17612
rect 11452 17587 11508 17599
rect 11900 17444 11956 17612
rect 12236 17639 12292 17724
rect 12236 17587 12238 17639
rect 12290 17587 12292 17639
rect 12236 17575 12292 17587
rect 12572 17666 12628 17678
rect 12572 17614 12574 17666
rect 12626 17614 12628 17666
rect 12572 17556 12628 17614
rect 11900 17378 11956 17388
rect 12012 17498 12068 17510
rect 12012 17446 12014 17498
rect 12066 17446 12068 17498
rect 12572 17490 12628 17500
rect 11228 17042 11284 17052
rect 8708 16902 8764 16940
rect 8820 16940 8932 16996
rect 9436 16996 9492 17006
rect 8820 16772 8876 16940
rect 9436 16882 9492 16940
rect 9436 16830 9438 16882
rect 9490 16830 9492 16882
rect 9436 16818 9492 16830
rect 10108 16884 10164 16894
rect 10108 16882 10276 16884
rect 10108 16830 10110 16882
rect 10162 16830 10276 16882
rect 10108 16828 10276 16830
rect 10108 16818 10164 16828
rect 8540 16158 8542 16210
rect 8594 16158 8596 16210
rect 8540 16146 8596 16158
rect 8764 16716 8876 16772
rect 7252 15988 7308 15998
rect 7252 15986 7364 15988
rect 7252 15934 7254 15986
rect 7306 15934 7364 15986
rect 7252 15922 7364 15934
rect 6524 14802 6580 14812
rect 6972 15036 7140 15092
rect 7196 15314 7252 15326
rect 7196 15262 7198 15314
rect 7250 15262 7252 15314
rect 5964 14478 5966 14530
rect 6018 14478 6020 14530
rect 5964 14466 6020 14478
rect 6076 14756 6132 14766
rect 5516 14354 5572 14364
rect 4844 14254 4846 14306
rect 4898 14254 4900 14306
rect 4844 14196 4900 14254
rect 4844 14140 5236 14196
rect 2604 13748 2660 13758
rect 2604 13746 2772 13748
rect 2604 13694 2606 13746
rect 2658 13694 2772 13746
rect 2604 13692 2772 13694
rect 2604 13682 2660 13692
rect 2548 13188 2604 13198
rect 2548 13074 2604 13132
rect 2548 13022 2550 13074
rect 2602 13022 2604 13074
rect 2548 13010 2604 13022
rect 2716 12962 2772 13692
rect 3388 13634 3444 13646
rect 3388 13582 3390 13634
rect 3442 13582 3444 13634
rect 3388 13186 3444 13582
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 3388 13134 3390 13186
rect 3442 13134 3444 13186
rect 3388 13122 3444 13134
rect 4396 13188 4452 13198
rect 2716 12910 2718 12962
rect 2770 12910 2772 12962
rect 2716 12404 2772 12910
rect 3724 12964 3780 12974
rect 3724 12870 3780 12908
rect 4396 12962 4452 13132
rect 4396 12910 4398 12962
rect 4450 12910 4452 12962
rect 4396 12898 4452 12910
rect 4620 13074 4676 13086
rect 4620 13022 4622 13074
rect 4674 13022 4676 13074
rect 4060 12740 4116 12750
rect 4060 12738 4228 12740
rect 4060 12686 4062 12738
rect 4114 12686 4228 12738
rect 4060 12684 4228 12686
rect 4060 12674 4116 12684
rect 2716 12338 2772 12348
rect 1596 12178 1652 12236
rect 1596 12126 1598 12178
rect 1650 12126 1652 12178
rect 1596 10610 1652 12126
rect 2380 12066 2436 12078
rect 2380 12014 2382 12066
rect 2434 12014 2436 12066
rect 2380 11618 2436 12014
rect 2380 11566 2382 11618
rect 2434 11566 2436 11618
rect 2380 11554 2436 11566
rect 3500 11506 3556 11518
rect 3500 11454 3502 11506
rect 3554 11454 3556 11506
rect 2716 11396 2772 11406
rect 2716 11302 2772 11340
rect 3164 11394 3220 11406
rect 3164 11342 3166 11394
rect 3218 11342 3220 11394
rect 3164 10836 3220 11342
rect 3388 11350 3444 11362
rect 3388 11298 3390 11350
rect 3442 11298 3444 11350
rect 3388 11284 3444 11298
rect 3388 11218 3444 11228
rect 3164 10770 3220 10780
rect 1596 10558 1598 10610
rect 1650 10558 1652 10610
rect 1596 10546 1652 10558
rect 3500 10612 3556 11454
rect 3948 11396 4004 11406
rect 3948 11226 4004 11340
rect 3948 11174 3950 11226
rect 4002 11174 4004 11226
rect 3948 11162 4004 11174
rect 4060 11394 4116 11406
rect 4060 11342 4062 11394
rect 4114 11342 4116 11394
rect 4060 11284 4116 11342
rect 4060 10612 4116 11228
rect 3500 10556 4004 10612
rect 2380 10498 2436 10510
rect 2380 10446 2382 10498
rect 2434 10446 2436 10498
rect 2380 10050 2436 10446
rect 2380 9998 2382 10050
rect 2434 9998 2436 10050
rect 2380 9986 2436 9998
rect 3724 10052 3780 10062
rect 2716 9828 2772 9838
rect 2716 9734 2772 9772
rect 3612 9828 3668 9838
rect 3612 9658 3668 9772
rect 3612 9606 3614 9658
rect 3666 9606 3668 9658
rect 3612 9594 3668 9606
rect 3724 9826 3780 9996
rect 3724 9774 3726 9826
rect 3778 9774 3780 9826
rect 1596 9042 1652 9054
rect 1596 8990 1598 9042
rect 1650 8990 1652 9042
rect 1596 7700 1652 8990
rect 2380 8930 2436 8942
rect 2380 8878 2382 8930
rect 2434 8878 2436 8930
rect 2380 8372 2436 8878
rect 2380 8306 2436 8316
rect 3388 8708 3444 8718
rect 3388 8230 3444 8652
rect 3724 8708 3780 9774
rect 3948 9787 4004 10556
rect 4060 10546 4116 10556
rect 4172 10276 4228 12684
rect 4284 12180 4340 12190
rect 4284 12086 4340 12124
rect 4620 11956 4676 13022
rect 5068 12962 5124 12974
rect 4788 12906 4844 12918
rect 4788 12854 4790 12906
rect 4842 12854 4844 12906
rect 4788 12852 4844 12854
rect 5068 12910 5070 12962
rect 5122 12910 5124 12962
rect 4788 12796 4900 12852
rect 4340 11900 4676 11956
rect 4844 12068 4900 12796
rect 4340 11844 4396 11900
rect 4284 11788 4396 11844
rect 4476 11788 4740 11798
rect 4284 11355 4340 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4844 11788 4900 12012
rect 4956 12205 5012 12217
rect 4956 12153 4958 12205
rect 5010 12153 5012 12205
rect 4956 11956 5012 12153
rect 5068 12180 5124 12910
rect 5180 12964 5236 14140
rect 6076 13790 6132 14700
rect 6412 14756 6468 14766
rect 6412 14642 6468 14700
rect 6412 14590 6414 14642
rect 6466 14590 6468 14642
rect 6412 14578 6468 14590
rect 6300 14532 6356 14542
rect 6300 14463 6302 14476
rect 6354 14463 6356 14476
rect 6300 14438 6356 14463
rect 6972 14532 7028 15036
rect 7084 14868 7140 14878
rect 7084 14532 7140 14812
rect 7196 14756 7252 15262
rect 7196 14690 7252 14700
rect 7196 14532 7252 14542
rect 7084 14530 7252 14532
rect 7084 14478 7198 14530
rect 7250 14478 7252 14530
rect 7084 14476 7252 14478
rect 6972 14450 6974 14476
rect 7026 14450 7028 14476
rect 5292 13748 5348 13758
rect 6076 13738 6078 13790
rect 6130 13738 6132 13790
rect 6748 14420 6804 14430
rect 6076 13726 6132 13738
rect 6412 13748 6468 13758
rect 5292 13654 5348 13692
rect 6412 13654 6468 13692
rect 5964 13634 6020 13646
rect 5964 13582 5966 13634
rect 6018 13582 6020 13634
rect 5628 12964 5684 12974
rect 5180 12962 5684 12964
rect 5180 12910 5630 12962
rect 5682 12910 5684 12962
rect 5180 12908 5684 12910
rect 5628 12898 5684 12908
rect 5740 12964 5796 12974
rect 5740 12794 5796 12908
rect 5964 12935 6020 13582
rect 5964 12883 5966 12935
rect 6018 12883 6020 12935
rect 5964 12871 6020 12883
rect 6076 13188 6132 13198
rect 5740 12742 5742 12794
rect 5794 12742 5796 12794
rect 5740 12730 5796 12742
rect 5068 12114 5124 12124
rect 5180 12292 5236 12302
rect 4956 11890 5012 11900
rect 5180 11844 5236 12236
rect 4844 11732 5124 11788
rect 5180 11778 5236 11788
rect 5628 12180 5684 12190
rect 4476 11722 4740 11732
rect 4284 11303 4286 11355
rect 4338 11303 4340 11355
rect 4284 11291 4340 11303
rect 4620 11394 4676 11406
rect 4620 11342 4622 11394
rect 4674 11342 4676 11394
rect 4284 10836 4340 10846
rect 4284 10722 4340 10780
rect 4284 10670 4286 10722
rect 4338 10670 4340 10722
rect 4284 10658 4340 10670
rect 4620 10388 4676 11342
rect 4788 10612 4844 10622
rect 4788 10518 4844 10556
rect 5068 10610 5124 11732
rect 5628 11394 5684 12124
rect 5628 11342 5630 11394
rect 5682 11342 5684 11394
rect 5404 10836 5460 10846
rect 5068 10558 5070 10610
rect 5122 10558 5124 10610
rect 5068 10546 5124 10558
rect 5292 10724 5348 10734
rect 5292 10610 5348 10668
rect 5292 10558 5294 10610
rect 5346 10558 5348 10610
rect 5292 10546 5348 10558
rect 4340 10332 4676 10388
rect 4340 10276 4396 10332
rect 4172 10220 4396 10276
rect 4476 10220 4740 10230
rect 4284 9828 4340 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 3948 9735 3950 9787
rect 4002 9735 4004 9787
rect 3948 9723 4004 9735
rect 4172 9826 4340 9828
rect 4172 9774 4286 9826
rect 4338 9774 4340 9826
rect 4172 9772 4340 9774
rect 3724 8642 3780 8652
rect 3388 8178 3390 8230
rect 3442 8178 3444 8230
rect 3612 8484 3668 8494
rect 4172 8428 4228 9772
rect 4284 9762 4340 9772
rect 4732 9940 4788 9950
rect 4284 9044 4340 9054
rect 4732 9044 4788 9884
rect 5404 9828 5460 10780
rect 5628 10724 5684 11342
rect 5628 10658 5684 10668
rect 5740 11506 5796 11518
rect 5740 11454 5742 11506
rect 5794 11454 5796 11506
rect 5572 10386 5628 10398
rect 5572 10334 5574 10386
rect 5626 10334 5628 10386
rect 5572 10052 5628 10334
rect 5572 9986 5628 9996
rect 5628 9828 5684 9838
rect 5404 9826 5684 9828
rect 5404 9774 5630 9826
rect 5682 9774 5684 9826
rect 5404 9772 5684 9774
rect 5628 9762 5684 9772
rect 5740 9716 5796 11454
rect 5964 11338 6020 11350
rect 5964 11286 5966 11338
rect 6018 11286 6020 11338
rect 5964 10836 6020 11286
rect 5852 10612 5908 10622
rect 5852 10518 5908 10556
rect 5964 10610 6020 10780
rect 5964 10558 5966 10610
rect 6018 10558 6020 10610
rect 5964 10546 6020 10558
rect 6076 9940 6132 13132
rect 6300 12962 6356 12974
rect 6300 12910 6302 12962
rect 6354 12910 6356 12962
rect 6300 12852 6356 12910
rect 6300 12786 6356 12796
rect 6636 12852 6692 12862
rect 6412 12404 6468 12414
rect 6412 12310 6468 12348
rect 6300 11396 6356 11406
rect 6300 11302 6356 11340
rect 6636 11396 6692 12796
rect 6748 11732 6804 14364
rect 6972 13746 7028 14450
rect 6972 13694 6974 13746
rect 7026 13694 7028 13746
rect 7196 13802 7252 14476
rect 7196 13750 7198 13802
rect 7250 13750 7252 13802
rect 7196 13738 7252 13750
rect 6972 13682 7028 13694
rect 7308 13636 7364 15922
rect 8036 15316 8092 15326
rect 8036 15222 8092 15260
rect 8764 15148 8820 16716
rect 9772 16660 9828 16670
rect 9772 16566 9828 16604
rect 9716 15540 9772 15550
rect 7476 15092 7532 15102
rect 8652 15092 8820 15148
rect 9548 15538 9772 15540
rect 9548 15486 9718 15538
rect 9770 15486 9772 15538
rect 9548 15484 9772 15486
rect 7476 15090 7644 15092
rect 7476 15038 7478 15090
rect 7530 15038 7644 15090
rect 7476 15036 7644 15038
rect 7476 15026 7532 15036
rect 7420 14644 7476 14654
rect 7420 14550 7476 14588
rect 7588 14586 7644 15036
rect 7588 14534 7590 14586
rect 7642 14534 7644 14586
rect 8540 14644 8596 14654
rect 8540 14550 8596 14588
rect 7588 14522 7644 14534
rect 7756 14532 7812 14542
rect 7756 14438 7812 14476
rect 8036 13972 8092 13982
rect 7756 13970 8092 13972
rect 7196 13580 7364 13636
rect 7420 13914 7476 13926
rect 7420 13862 7422 13914
rect 7474 13862 7476 13914
rect 6972 12964 7028 12974
rect 6972 12870 7028 12908
rect 7196 12962 7252 13580
rect 7196 12910 7198 12962
rect 7250 12910 7252 12962
rect 7196 12898 7252 12910
rect 7308 13130 7364 13142
rect 7308 13078 7310 13130
rect 7362 13078 7364 13130
rect 6748 11666 6804 11676
rect 7196 11562 7252 11574
rect 7196 11510 7198 11562
rect 7250 11510 7252 11562
rect 6636 11394 7140 11396
rect 6636 11342 6638 11394
rect 6690 11342 7140 11394
rect 6636 11340 7140 11342
rect 6636 11330 6692 11340
rect 6188 10724 6244 10734
rect 6188 10610 6244 10668
rect 6188 10558 6190 10610
rect 6242 10558 6244 10610
rect 6188 10546 6244 10558
rect 6412 10610 6468 10622
rect 6412 10558 6414 10610
rect 6466 10558 6468 10610
rect 6300 10388 6356 10398
rect 6076 9884 6244 9940
rect 6076 9770 6132 9782
rect 6076 9718 6078 9770
rect 6130 9718 6132 9770
rect 5740 9660 6020 9716
rect 5818 9268 5874 9278
rect 4284 9042 4788 9044
rect 4284 8990 4286 9042
rect 4338 8990 4734 9042
rect 4786 8990 4788 9042
rect 4284 8988 4788 8990
rect 4284 8978 4340 8988
rect 4732 8820 4788 8988
rect 4900 9210 4956 9222
rect 4900 9158 4902 9210
rect 4954 9158 4956 9210
rect 4900 9044 4956 9158
rect 5818 9080 5874 9212
rect 4900 8978 4956 8988
rect 5628 9044 5684 9054
rect 5818 9028 5820 9080
rect 5872 9028 5874 9080
rect 5818 9016 5874 9028
rect 5964 9042 6020 9660
rect 6076 9268 6132 9718
rect 6188 9492 6244 9884
rect 6300 9826 6356 10332
rect 6412 9940 6468 10558
rect 6692 10388 6748 10398
rect 7084 10388 7140 11340
rect 7196 10612 7252 11510
rect 7308 11394 7364 13078
rect 7420 12404 7476 13862
rect 7756 13918 8038 13970
rect 8090 13918 8092 13970
rect 7756 13916 8092 13918
rect 7532 13748 7588 13758
rect 7756 13748 7812 13916
rect 8036 13906 8092 13916
rect 7532 13746 7812 13748
rect 7532 13694 7534 13746
rect 7586 13694 7812 13746
rect 7532 13692 7812 13694
rect 7868 13748 7924 13758
rect 7532 12964 7588 13692
rect 7868 13654 7924 13692
rect 7812 13524 7868 13534
rect 7812 13186 7868 13468
rect 8652 13300 8708 15092
rect 9548 14868 9604 15484
rect 9716 15474 9772 15484
rect 9884 15334 9940 15346
rect 9548 14802 9604 14812
rect 9772 15316 9828 15326
rect 9660 13914 9716 13926
rect 9660 13862 9662 13914
rect 9714 13862 9716 13914
rect 9100 13748 9156 13758
rect 9548 13748 9604 13758
rect 9100 13654 9156 13692
rect 9324 13746 9604 13748
rect 9324 13694 9550 13746
rect 9602 13694 9604 13746
rect 9324 13692 9604 13694
rect 8764 13524 8820 13534
rect 8764 13522 9268 13524
rect 8764 13470 8766 13522
rect 8818 13470 9268 13522
rect 8764 13468 9268 13470
rect 8764 13458 8820 13468
rect 8988 13300 9044 13310
rect 8652 13244 8820 13300
rect 7812 13134 7814 13186
rect 7866 13134 7868 13186
rect 7812 13122 7868 13134
rect 7532 12898 7588 12908
rect 8092 12962 8148 12974
rect 8092 12910 8094 12962
rect 8146 12910 8148 12962
rect 8092 12852 8148 12910
rect 8092 12786 8148 12796
rect 8316 12962 8372 12974
rect 8316 12910 8318 12962
rect 8370 12910 8372 12962
rect 7420 12348 7700 12404
rect 7532 12180 7588 12190
rect 7308 11342 7310 11394
rect 7362 11342 7364 11394
rect 7308 11330 7364 11342
rect 7420 11956 7476 11966
rect 7196 10556 7364 10612
rect 7196 10388 7252 10398
rect 7084 10386 7252 10388
rect 7084 10334 7198 10386
rect 7250 10334 7252 10386
rect 7084 10332 7252 10334
rect 6692 10294 6748 10332
rect 7196 10322 7252 10332
rect 6412 9874 6468 9884
rect 6300 9774 6302 9826
rect 6354 9774 6356 9826
rect 6300 9762 6356 9774
rect 7308 9793 7364 10556
rect 7308 9741 7310 9793
rect 7362 9741 7364 9793
rect 7308 9729 7364 9741
rect 6412 9716 6468 9726
rect 6412 9658 6468 9660
rect 6412 9606 6414 9658
rect 6466 9606 6468 9658
rect 6412 9594 6468 9606
rect 6188 9436 6636 9492
rect 6580 9268 6636 9436
rect 6076 9212 6468 9268
rect 4732 8764 4900 8820
rect 3612 8258 3668 8428
rect 3612 8206 3614 8258
rect 3666 8206 3668 8258
rect 3612 8194 3668 8206
rect 3724 8372 4228 8428
rect 4284 8708 4340 8718
rect 4284 8428 4340 8652
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4732 8484 4788 8494
rect 4844 8428 4900 8764
rect 5404 8818 5460 8830
rect 5404 8766 5406 8818
rect 5458 8766 5460 8818
rect 5404 8428 5460 8766
rect 4284 8372 4452 8428
rect 3388 8166 3444 8178
rect 3724 7924 3780 8372
rect 4396 8220 4452 8372
rect 4004 8202 4060 8214
rect 3612 7868 3780 7924
rect 3836 8146 3892 8158
rect 3836 8094 3838 8146
rect 3890 8094 3892 8146
rect 1596 7474 1652 7644
rect 1596 7422 1598 7474
rect 1650 7422 1652 7474
rect 1596 7410 1652 7422
rect 2268 7700 2324 7710
rect 2268 5122 2324 7644
rect 2380 7362 2436 7374
rect 2380 7310 2382 7362
rect 2434 7310 2436 7362
rect 2380 6916 2436 7310
rect 2492 6916 2548 6926
rect 2380 6914 2548 6916
rect 2380 6862 2494 6914
rect 2546 6862 2548 6914
rect 2380 6860 2548 6862
rect 2492 6850 2548 6860
rect 2828 6692 2884 6702
rect 2828 6598 2884 6636
rect 3612 6468 3668 7868
rect 3724 7700 3780 7710
rect 3724 6690 3780 7644
rect 3724 6638 3726 6690
rect 3778 6638 3780 6690
rect 3724 6626 3780 6638
rect 3836 6580 3892 8094
rect 4004 8150 4006 8202
rect 4058 8150 4060 8202
rect 4396 8168 4398 8220
rect 4450 8168 4452 8220
rect 4732 8372 4900 8428
rect 4956 8372 5012 8382
rect 4732 8258 4788 8372
rect 4956 8278 5012 8316
rect 5124 8372 5460 8428
rect 5124 8314 5180 8372
rect 4732 8206 4734 8258
rect 4786 8206 4788 8258
rect 5124 8262 5126 8314
rect 5178 8262 5180 8314
rect 5124 8250 5180 8262
rect 5628 8258 5684 8988
rect 5964 8990 5966 9042
rect 6018 8990 6020 9042
rect 5964 8428 6020 8990
rect 6076 9044 6132 9054
rect 6076 8950 6132 8988
rect 5964 8372 6356 8428
rect 4732 8194 4788 8206
rect 5628 8206 5630 8258
rect 5682 8206 5684 8258
rect 6300 8258 6356 8372
rect 5628 8194 5684 8206
rect 6076 8202 6132 8214
rect 4396 8156 4452 8168
rect 4004 8036 4060 8150
rect 6076 8150 6078 8202
rect 6130 8150 6132 8202
rect 6300 8206 6302 8258
rect 6354 8206 6356 8258
rect 6300 8194 6356 8206
rect 4004 7970 4060 7980
rect 4284 8036 4340 8046
rect 4284 7362 4340 7980
rect 4284 7310 4286 7362
rect 4338 7310 4340 7362
rect 4284 6916 4340 7310
rect 5852 7700 5908 7710
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4284 6850 4340 6860
rect 4956 6804 5012 6814
rect 3836 6514 3892 6524
rect 4620 6690 4676 6702
rect 4620 6638 4622 6690
rect 4674 6638 4676 6690
rect 3612 6402 3668 6412
rect 4620 5796 4676 6638
rect 4956 6675 5012 6748
rect 4956 6623 4958 6675
rect 5010 6623 5012 6675
rect 4956 6611 5012 6623
rect 5068 6802 5124 6814
rect 5068 6750 5070 6802
rect 5122 6750 5124 6802
rect 5068 6580 5124 6750
rect 5628 6690 5684 6702
rect 5628 6638 5630 6690
rect 5682 6638 5684 6690
rect 5068 6524 5236 6580
rect 4732 6076 5124 6132
rect 4732 5906 4788 6076
rect 5068 6074 5124 6076
rect 5068 6022 5070 6074
rect 5122 6022 5124 6074
rect 5068 6010 5124 6022
rect 5180 6020 5236 6524
rect 5628 6468 5684 6638
rect 5740 6692 5796 6702
rect 5740 6522 5796 6636
rect 5740 6470 5742 6522
rect 5794 6470 5796 6522
rect 5740 6458 5796 6470
rect 5628 6402 5684 6412
rect 5740 6244 5796 6254
rect 5628 6132 5684 6142
rect 5180 5964 5292 6020
rect 5236 5962 5292 5964
rect 4732 5854 4734 5906
rect 4786 5854 4788 5906
rect 4732 5842 4788 5854
rect 4956 5908 5012 5918
rect 5236 5910 5238 5962
rect 5290 5910 5292 5962
rect 5236 5898 5292 5910
rect 5628 5906 5684 6076
rect 4956 5814 5012 5852
rect 5628 5854 5630 5906
rect 5682 5854 5684 5906
rect 5628 5842 5684 5854
rect 4620 5730 4676 5740
rect 3052 5684 3108 5694
rect 3052 5234 3108 5628
rect 4396 5684 4452 5722
rect 4396 5618 4452 5628
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 3052 5182 3054 5234
rect 3106 5182 3108 5234
rect 3052 5170 3108 5182
rect 4956 5236 5012 5246
rect 4956 5142 5012 5180
rect 5740 5236 5796 6188
rect 5852 5348 5908 7644
rect 6076 6692 6132 8150
rect 5964 6634 6020 6646
rect 5964 6582 5966 6634
rect 6018 6582 6020 6634
rect 6076 6626 6132 6636
rect 6188 8090 6244 8102
rect 6188 8038 6190 8090
rect 6242 8038 6244 8090
rect 5964 6580 6020 6582
rect 5964 6514 6020 6524
rect 6076 5906 6132 5918
rect 6076 5854 6078 5906
rect 6130 5854 6132 5906
rect 6076 5796 6132 5854
rect 6188 5908 6244 8038
rect 6300 6804 6356 6814
rect 6300 6690 6356 6748
rect 6300 6638 6302 6690
rect 6354 6638 6356 6690
rect 6300 6356 6356 6638
rect 6300 6290 6356 6300
rect 6412 6244 6468 9212
rect 6580 9174 6636 9212
rect 7084 9268 7140 9278
rect 7420 9268 7476 11900
rect 7532 11396 7588 12124
rect 7532 11302 7588 11340
rect 7644 12178 7700 12348
rect 7644 12126 7646 12178
rect 7698 12126 7700 12178
rect 7532 10612 7588 10622
rect 7644 10612 7700 12126
rect 8316 12180 8372 12910
rect 8316 12114 8372 12124
rect 8428 12962 8484 12974
rect 8428 12910 8430 12962
rect 8482 12910 8484 12962
rect 8428 12404 8484 12910
rect 7924 12068 7980 12078
rect 7924 11974 7980 12012
rect 8428 11844 8484 12348
rect 8652 12178 8708 12190
rect 8652 12126 8654 12178
rect 8706 12126 8708 12178
rect 8652 12068 8708 12126
rect 8652 12002 8708 12012
rect 8540 11844 8596 11854
rect 8428 11788 8540 11844
rect 7868 11732 7924 11742
rect 7868 11394 7924 11676
rect 7868 11342 7870 11394
rect 7922 11342 7924 11394
rect 7868 11172 7924 11342
rect 8540 11394 8596 11788
rect 8540 11342 8542 11394
rect 8594 11342 8596 11394
rect 8540 11330 8596 11342
rect 8204 11284 8260 11294
rect 8204 11190 8260 11228
rect 7868 11106 7924 11116
rect 8092 10836 8148 10846
rect 8092 10742 8148 10780
rect 7532 10610 7700 10612
rect 7532 10558 7534 10610
rect 7586 10558 7700 10610
rect 7532 10556 7700 10558
rect 8428 10612 8484 10622
rect 7532 10546 7588 10556
rect 8428 10518 8484 10556
rect 8540 10610 8596 10622
rect 8540 10558 8542 10610
rect 8594 10558 8596 10610
rect 8402 9828 8458 9838
rect 7084 9174 7140 9212
rect 7196 9212 7476 9268
rect 7756 9770 7812 9782
rect 7756 9718 7758 9770
rect 7810 9718 7812 9770
rect 7196 8428 7252 9212
rect 7420 9044 7476 9054
rect 7420 8950 7476 8988
rect 7196 8370 7308 8428
rect 7196 8318 7254 8370
rect 7306 8318 7308 8370
rect 7196 8278 7308 8318
rect 7196 7501 7252 8278
rect 7420 8258 7476 8270
rect 7420 8206 7422 8258
rect 7474 8206 7476 8258
rect 7420 7700 7476 8206
rect 7756 8260 7812 9718
rect 8092 9770 8148 9782
rect 8092 9718 8094 9770
rect 8146 9718 8148 9770
rect 8402 9741 8404 9772
rect 8456 9741 8458 9772
rect 8402 9729 8458 9741
rect 8092 9716 8148 9718
rect 8092 9650 8148 9660
rect 8540 9714 8596 10558
rect 8540 9662 8542 9714
rect 8594 9662 8596 9714
rect 8540 9604 8596 9662
rect 8204 9548 8596 9604
rect 7868 9044 7924 9054
rect 7868 8820 7924 8988
rect 8204 9042 8260 9548
rect 8204 8990 8206 9042
rect 8258 8990 8260 9042
rect 8204 8978 8260 8990
rect 8316 9042 8372 9054
rect 8316 8990 8318 9042
rect 8370 8990 8372 9042
rect 8316 8820 8372 8990
rect 7868 8818 8372 8820
rect 7868 8766 7870 8818
rect 7922 8766 8372 8818
rect 7868 8764 8372 8766
rect 7868 8754 7924 8764
rect 7756 8194 7812 8204
rect 8204 8258 8260 8270
rect 8204 8206 8206 8258
rect 8258 8206 8260 8258
rect 7420 7634 7476 7644
rect 7588 7700 7644 7710
rect 7588 7698 8036 7700
rect 7588 7646 7590 7698
rect 7642 7646 8036 7698
rect 7588 7644 8036 7646
rect 7588 7634 7644 7644
rect 7196 7449 7198 7501
rect 7250 7449 7252 7501
rect 7980 7530 8036 7644
rect 7196 7437 7252 7449
rect 7756 7476 7812 7486
rect 7980 7478 7982 7530
rect 8034 7478 8036 7530
rect 8204 7588 8260 8206
rect 7756 7474 7924 7476
rect 7756 7422 7758 7474
rect 7810 7422 7924 7474
rect 7980 7466 8036 7478
rect 8092 7512 8148 7524
rect 8204 7522 8260 7532
rect 8092 7476 8094 7512
rect 8146 7476 8148 7512
rect 7756 7420 7924 7422
rect 7756 7410 7812 7420
rect 7756 7028 7812 7038
rect 7084 6916 7140 6926
rect 6916 6692 6972 6702
rect 6916 6522 6972 6636
rect 7084 6690 7140 6860
rect 7756 6802 7812 6972
rect 7756 6750 7758 6802
rect 7810 6750 7812 6802
rect 7756 6738 7812 6750
rect 7084 6638 7086 6690
rect 7138 6638 7140 6690
rect 7084 6626 7140 6638
rect 7420 6690 7476 6702
rect 7420 6638 7422 6690
rect 7474 6638 7476 6690
rect 7868 6692 7924 7420
rect 8092 7028 8148 7420
rect 8092 6962 8148 6972
rect 8092 6692 8148 6702
rect 6916 6470 6918 6522
rect 6970 6470 6972 6522
rect 6916 6458 6972 6470
rect 6412 6178 6468 6188
rect 6860 6356 6916 6366
rect 6580 6132 6636 6142
rect 6580 6018 6636 6076
rect 6580 5966 6582 6018
rect 6634 5966 6636 6018
rect 6580 5954 6636 5966
rect 6300 5908 6356 5918
rect 6188 5906 6468 5908
rect 6188 5854 6302 5906
rect 6354 5854 6468 5906
rect 6188 5852 6468 5854
rect 6300 5842 6356 5852
rect 6132 5740 6244 5796
rect 6076 5730 6132 5740
rect 5852 5292 6132 5348
rect 2268 5070 2270 5122
rect 2322 5070 2324 5122
rect 2268 5058 2324 5070
rect 5740 5124 5796 5180
rect 5852 5124 5908 5134
rect 5740 5122 5908 5124
rect 5740 5070 5854 5122
rect 5906 5070 5908 5122
rect 5740 5068 5908 5070
rect 5852 5058 5908 5068
rect 6076 4340 6132 5292
rect 6188 5346 6244 5740
rect 6188 5294 6190 5346
rect 6242 5294 6244 5346
rect 6188 5282 6244 5294
rect 6412 5124 6468 5852
rect 6860 5346 6916 6300
rect 7420 6132 7476 6638
rect 7756 6634 7812 6646
rect 7756 6582 7758 6634
rect 7810 6582 7812 6634
rect 7868 6626 7924 6636
rect 7980 6690 8148 6692
rect 7980 6638 8094 6690
rect 8146 6638 8148 6690
rect 7980 6636 8148 6638
rect 7140 6076 7476 6132
rect 7532 6356 7588 6366
rect 6972 5908 7028 5918
rect 6972 5814 7028 5852
rect 7140 5850 7196 6076
rect 7532 6020 7588 6300
rect 7420 5964 7588 6020
rect 7756 6020 7812 6582
rect 7980 6356 8036 6636
rect 8092 6626 8148 6636
rect 8316 6468 8372 8764
rect 8652 8820 8708 8830
rect 8764 8820 8820 13244
rect 8876 12852 8932 12862
rect 8876 12222 8932 12796
rect 8876 12170 8878 12222
rect 8930 12170 8932 12222
rect 8876 12158 8932 12170
rect 8988 12066 9044 13244
rect 9212 13074 9268 13468
rect 9212 13022 9214 13074
rect 9266 13022 9268 13074
rect 9212 13010 9268 13022
rect 9324 12852 9380 13692
rect 9548 13682 9604 13692
rect 9660 13748 9716 13862
rect 9660 13682 9716 13692
rect 9772 13412 9828 15260
rect 9884 15282 9886 15334
rect 9938 15282 9940 15334
rect 9884 14644 9940 15282
rect 9884 14578 9940 14588
rect 9996 15316 10052 15326
rect 10220 15316 10276 16828
rect 10892 16770 10948 16782
rect 10892 16718 10894 16770
rect 10946 16718 10948 16770
rect 10444 16660 10500 16670
rect 10444 16210 10500 16604
rect 10892 16324 10948 16718
rect 10892 16258 10948 16268
rect 11004 16772 11060 16782
rect 10444 16158 10446 16210
rect 10498 16158 10500 16210
rect 10444 16146 10500 16158
rect 9996 15314 10276 15316
rect 9996 15262 9998 15314
rect 10050 15262 10276 15314
rect 9996 15260 10276 15262
rect 11004 15876 11060 16716
rect 11676 16324 11732 16334
rect 11676 16230 11732 16268
rect 11004 15341 11060 15820
rect 11004 15316 11006 15341
rect 11058 15316 11060 15341
rect 9996 15092 10052 15260
rect 11004 15211 11060 15260
rect 11228 16098 11284 16110
rect 11228 16046 11230 16098
rect 11282 16046 11284 16098
rect 11228 15092 11284 16046
rect 12012 16098 12068 17446
rect 12796 17108 12852 18060
rect 13132 17668 13188 18396
rect 13356 17892 13412 18396
rect 13468 18450 13580 18462
rect 13468 18398 13470 18450
rect 13522 18398 13580 18450
rect 13468 18396 13580 18398
rect 13748 18450 13804 19068
rect 13916 18900 13972 19182
rect 14028 19234 14084 20860
rect 14476 20804 14532 20814
rect 14028 19182 14030 19234
rect 14082 19182 14084 19234
rect 14028 19170 14084 19182
rect 14194 19796 14250 19806
rect 14194 19234 14250 19740
rect 14194 19182 14196 19234
rect 14248 19182 14250 19234
rect 14194 19170 14250 19182
rect 14476 19794 14532 20748
rect 14588 20802 14644 21644
rect 14588 20750 14590 20802
rect 14642 20750 14644 20802
rect 14588 20738 14644 20750
rect 14700 20970 14756 20982
rect 14700 20918 14702 20970
rect 14754 20918 14756 20970
rect 14700 20244 14756 20918
rect 14924 20804 14980 22318
rect 15148 21924 15204 21934
rect 15148 21698 15204 21868
rect 15148 21646 15150 21698
rect 15202 21646 15204 21698
rect 15148 21634 15204 21646
rect 15484 21700 15540 23100
rect 16156 23156 16212 24444
rect 16604 23940 16660 24670
rect 16604 23874 16660 23884
rect 16716 24500 16772 24510
rect 16716 23938 16772 24444
rect 16996 24164 17052 24174
rect 16996 24070 17052 24108
rect 17164 23940 17220 26460
rect 17276 26290 17332 26852
rect 17276 26238 17278 26290
rect 17330 26238 17332 26290
rect 17276 26226 17332 26238
rect 17388 27300 17444 27310
rect 17388 26964 17444 27244
rect 17500 27188 17556 27806
rect 17612 28026 17668 28038
rect 17612 27974 17614 28026
rect 17666 27974 17668 28026
rect 17612 27524 17668 27974
rect 17836 27914 17892 28028
rect 17836 27862 17838 27914
rect 17890 27862 17892 27914
rect 17836 27850 17892 27862
rect 17948 27636 18004 30492
rect 18284 30436 18340 30986
rect 18396 30940 18564 30996
rect 18956 31108 19012 31118
rect 18956 30994 19012 31052
rect 19124 31110 19126 31162
rect 19178 31110 19180 31162
rect 19124 31108 19180 31110
rect 19124 31042 19180 31052
rect 18956 30942 18958 30994
rect 19010 30942 19012 30994
rect 18396 30548 18452 30940
rect 18620 30884 18676 30894
rect 18508 30772 18564 30782
rect 18620 30772 18676 30828
rect 18508 30770 18676 30772
rect 18508 30718 18510 30770
rect 18562 30718 18676 30770
rect 18508 30716 18676 30718
rect 18844 30884 18900 30894
rect 18956 30884 19012 30942
rect 19404 30996 19460 31006
rect 19404 30902 19460 30940
rect 19628 30996 19684 31006
rect 19628 30902 19684 30940
rect 20188 30996 20244 31500
rect 20300 31890 20580 31892
rect 20300 31838 20526 31890
rect 20578 31838 20580 31890
rect 20300 31836 20580 31838
rect 20300 31050 20356 31836
rect 20524 31826 20580 31836
rect 20636 31668 20692 32274
rect 20860 32004 20916 32510
rect 20860 31938 20916 31948
rect 20748 31668 20804 31678
rect 20636 31612 20748 31668
rect 20300 30998 20302 31050
rect 20354 30998 20356 31050
rect 20300 30986 20356 30998
rect 20412 31108 20468 31118
rect 20412 31050 20468 31052
rect 20412 30998 20414 31050
rect 20466 30998 20468 31050
rect 20412 30986 20468 30998
rect 20636 31022 20692 31034
rect 20188 30930 20244 30940
rect 20636 30970 20638 31022
rect 20690 30970 20692 31022
rect 20636 30884 20692 30970
rect 18956 30828 19124 30884
rect 18508 30706 18564 30716
rect 18396 30492 18676 30548
rect 18284 30380 18452 30436
rect 18172 30322 18228 30334
rect 18172 30270 18174 30322
rect 18226 30270 18228 30322
rect 18172 30212 18228 30270
rect 18396 30212 18452 30380
rect 18172 30146 18228 30156
rect 18284 30166 18340 30178
rect 18284 30114 18286 30166
rect 18338 30114 18340 30166
rect 18396 30146 18452 30156
rect 18620 30210 18676 30492
rect 18844 30380 18900 30828
rect 19068 30548 19124 30828
rect 20636 30818 20692 30828
rect 19908 30772 19964 30782
rect 19908 30770 20132 30772
rect 19908 30718 19910 30770
rect 19962 30718 20132 30770
rect 19908 30716 20132 30718
rect 19908 30706 19964 30716
rect 19068 30482 19124 30492
rect 19348 30436 19404 30446
rect 18844 30324 19124 30380
rect 18620 30158 18622 30210
rect 18674 30158 18676 30210
rect 18284 30100 18340 30114
rect 18060 29314 18116 29326
rect 18060 29262 18062 29314
rect 18114 29262 18116 29314
rect 18060 28980 18116 29262
rect 18060 28914 18116 28924
rect 18060 28644 18116 28654
rect 18060 28550 18116 28588
rect 18284 28084 18340 30044
rect 18620 29988 18676 30158
rect 18620 29922 18676 29932
rect 18844 30210 18900 30222
rect 18844 30158 18846 30210
rect 18898 30158 18900 30210
rect 18844 29876 18900 30158
rect 19068 30210 19124 30324
rect 19068 30158 19070 30210
rect 19122 30158 19124 30210
rect 19068 30146 19124 30158
rect 19348 30210 19404 30380
rect 19348 30158 19350 30210
rect 19402 30158 19404 30210
rect 19348 30146 19404 30158
rect 19908 30212 19964 30222
rect 19908 30118 19964 30156
rect 18844 29810 18900 29820
rect 19292 29988 19348 29998
rect 18396 28980 18452 28990
rect 18396 28866 18452 28924
rect 18396 28814 18398 28866
rect 18450 28814 18452 28866
rect 18396 28802 18452 28814
rect 18508 28868 18564 28878
rect 18284 28018 18340 28028
rect 18060 27860 18116 27898
rect 18060 27794 18116 27804
rect 18060 27636 18116 27646
rect 17948 27580 18060 27636
rect 17612 27468 18004 27524
rect 17612 27300 17668 27310
rect 17836 27300 17892 27310
rect 17668 27244 17780 27300
rect 17612 27234 17668 27244
rect 17500 27122 17556 27132
rect 17724 27074 17780 27244
rect 17556 27018 17612 27030
rect 17556 26966 17558 27018
rect 17610 26966 17612 27018
rect 17724 27022 17726 27074
rect 17778 27022 17780 27074
rect 17724 27010 17780 27022
rect 17836 27074 17892 27244
rect 17836 27022 17838 27074
rect 17890 27022 17892 27074
rect 17556 26908 17612 26966
rect 17388 24948 17444 26908
rect 17500 26852 17612 26908
rect 17500 26516 17556 26852
rect 17500 26450 17556 26460
rect 17612 26740 17668 26750
rect 17612 26514 17668 26684
rect 17612 26462 17614 26514
rect 17666 26462 17668 26514
rect 17612 26450 17668 26462
rect 17836 26292 17892 27022
rect 16716 23886 16718 23938
rect 16770 23886 16772 23938
rect 16380 23828 16436 23838
rect 16380 23734 16436 23772
rect 16716 23716 16772 23886
rect 17052 23884 17220 23940
rect 17276 24892 17444 24948
rect 17500 26236 17892 26292
rect 17948 26290 18004 27468
rect 17948 26238 17950 26290
rect 18002 26238 18004 26290
rect 17276 23938 17332 24892
rect 17276 23886 17278 23938
rect 17330 23886 17332 23938
rect 16716 23660 16996 23716
rect 16156 23090 16212 23100
rect 16492 23154 16548 23166
rect 16492 23102 16494 23154
rect 16546 23102 16548 23154
rect 15596 22930 15652 22942
rect 16156 22932 16212 22942
rect 15596 22878 15598 22930
rect 15650 22878 15652 22930
rect 15596 22372 15652 22878
rect 15708 22930 16212 22932
rect 15708 22878 16158 22930
rect 16210 22878 16212 22930
rect 15708 22876 16212 22878
rect 15708 22482 15764 22876
rect 16156 22866 16212 22876
rect 16492 22708 16548 23102
rect 16940 23064 16996 23660
rect 16884 23042 16996 23064
rect 16884 22990 16886 23042
rect 16938 22990 16996 23042
rect 16884 22978 16996 22990
rect 16492 22652 16884 22708
rect 15708 22430 15710 22482
rect 15762 22430 15764 22482
rect 15708 22418 15764 22430
rect 15596 22260 15652 22316
rect 15596 22204 15876 22260
rect 15484 21644 15689 21700
rect 15633 21642 15689 21644
rect 15633 21590 15635 21642
rect 15687 21590 15689 21642
rect 15633 21578 15689 21590
rect 15820 21642 15876 22204
rect 15820 21590 15822 21642
rect 15874 21590 15876 21642
rect 15820 21578 15876 21590
rect 16044 22148 16100 22158
rect 16828 22148 16884 22652
rect 16044 21642 16100 22092
rect 16548 22092 16884 22148
rect 16044 21590 16046 21642
rect 16098 21590 16100 21642
rect 16044 21578 16100 21590
rect 16268 21700 16324 21710
rect 16268 21642 16324 21644
rect 16268 21590 16270 21642
rect 16322 21590 16324 21642
rect 16548 21698 16604 22092
rect 16548 21646 16550 21698
rect 16602 21646 16604 21698
rect 16548 21634 16604 21646
rect 16268 21578 16324 21590
rect 15932 20804 15988 20814
rect 14924 20738 14980 20748
rect 15328 20764 15384 20776
rect 15328 20712 15330 20764
rect 15382 20712 15384 20764
rect 15328 20356 15384 20712
rect 15932 20722 15934 20748
rect 15986 20722 15988 20748
rect 15932 20710 15988 20722
rect 15328 20290 15384 20300
rect 16828 20356 16884 20366
rect 14700 20178 14756 20188
rect 16716 20020 16772 20030
rect 16716 19926 16772 19964
rect 16828 20018 16884 20300
rect 16828 19966 16830 20018
rect 16882 19966 16884 20018
rect 16828 19954 16884 19966
rect 16940 20020 16996 22978
rect 17052 21476 17108 23884
rect 17276 23268 17332 23886
rect 17276 23202 17332 23212
rect 17388 24722 17444 24734
rect 17388 24670 17390 24722
rect 17442 24670 17444 24722
rect 17388 23828 17444 24670
rect 17500 24500 17556 26236
rect 17948 26226 18004 26238
rect 17724 26068 17780 26078
rect 17724 25618 17780 26012
rect 18060 25844 18116 27580
rect 18340 27300 18396 27310
rect 18340 27186 18396 27244
rect 18340 27134 18342 27186
rect 18394 27134 18396 27186
rect 18340 27122 18396 27134
rect 18508 27076 18564 28812
rect 19292 28866 19348 29932
rect 20076 29988 20132 30716
rect 20412 30548 20468 30558
rect 20076 29922 20132 29932
rect 20300 30378 20356 30390
rect 20300 30326 20302 30378
rect 20354 30326 20356 30378
rect 19292 28814 19294 28866
rect 19346 28814 19348 28866
rect 19292 28802 19348 28814
rect 19404 29876 19460 29886
rect 19404 28196 19460 29820
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19628 29428 19684 29438
rect 19628 28642 19684 29372
rect 19964 29428 20020 29438
rect 19964 29334 20020 29372
rect 20300 28756 20356 30326
rect 20412 30210 20468 30492
rect 20412 30158 20414 30210
rect 20466 30158 20468 30210
rect 20412 30146 20468 30158
rect 20524 30324 20580 30334
rect 20300 28690 20356 28700
rect 19628 28590 19630 28642
rect 19682 28590 19684 28642
rect 19628 28578 19684 28590
rect 19068 28140 19460 28196
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 18900 27898 18956 27899
rect 18900 27887 19012 27898
rect 18732 27860 18788 27870
rect 18900 27835 18902 27887
rect 18954 27835 19012 27887
rect 18900 27823 19012 27835
rect 18732 27746 18788 27804
rect 18732 27694 18734 27746
rect 18786 27694 18788 27746
rect 18732 27682 18788 27694
rect 18956 27412 19012 27823
rect 18620 27076 18676 27086
rect 18508 27074 18676 27076
rect 18508 27022 18622 27074
rect 18674 27022 18676 27074
rect 18508 27020 18676 27022
rect 18620 27010 18676 27020
rect 18956 27047 19012 27356
rect 18956 26995 18958 27047
rect 19010 26995 19012 27047
rect 18956 26983 19012 26995
rect 19068 26908 19124 28140
rect 20412 28084 20468 28094
rect 20412 28026 20468 28028
rect 19628 27972 19684 27982
rect 20412 27974 20414 28026
rect 20466 27974 20468 28026
rect 20412 27962 20468 27974
rect 20524 27972 20580 30268
rect 20748 30210 20804 31612
rect 20860 31108 20916 31118
rect 20972 31108 21028 33292
rect 21084 32340 21140 34117
rect 21308 35140 21364 35150
rect 21532 35140 21588 35646
rect 21308 34130 21364 35084
rect 21308 34078 21310 34130
rect 21362 34078 21364 34130
rect 21308 34066 21364 34078
rect 21420 35084 21588 35140
rect 21644 35252 21700 35262
rect 21420 34804 21476 35084
rect 21420 34132 21476 34748
rect 21420 34066 21476 34076
rect 21532 34802 21588 34814
rect 21532 34750 21534 34802
rect 21586 34750 21588 34802
rect 21532 33572 21588 34750
rect 21644 34130 21700 35196
rect 21756 34692 21812 36530
rect 21980 38050 22036 40012
rect 22092 40012 22484 40068
rect 22092 38834 22148 40012
rect 22540 38892 22596 41132
rect 22876 41122 22932 41132
rect 22652 40964 22708 40974
rect 22652 40290 22708 40908
rect 22652 40238 22654 40290
rect 22706 40238 22708 40290
rect 22652 40226 22708 40238
rect 23100 39060 23156 42476
rect 23772 41970 23828 41982
rect 23772 41918 23774 41970
rect 23826 41918 23828 41970
rect 23212 41860 23268 41870
rect 23212 41130 23268 41804
rect 23772 41412 23828 41918
rect 23940 41748 23996 41758
rect 23940 41654 23996 41692
rect 23772 41356 23940 41412
rect 23548 41300 23604 41310
rect 23212 41078 23214 41130
rect 23266 41078 23268 41130
rect 23212 41076 23268 41078
rect 23212 41010 23268 41020
rect 23324 41188 23380 41198
rect 23324 40404 23380 41132
rect 23548 41186 23604 41244
rect 23548 41134 23550 41186
rect 23602 41134 23604 41186
rect 23548 41122 23604 41134
rect 23772 41186 23828 41198
rect 23772 41134 23774 41186
rect 23826 41134 23828 41186
rect 23436 41018 23492 41030
rect 23436 40966 23438 41018
rect 23490 40966 23492 41018
rect 23436 40964 23492 40966
rect 23772 40964 23828 41134
rect 23436 40908 23828 40964
rect 23884 40628 23940 41356
rect 24220 41076 24276 42812
rect 24332 42644 24388 42654
rect 24556 42644 24612 43484
rect 24780 42754 24836 43652
rect 24780 42702 24782 42754
rect 24834 42702 24836 42754
rect 24780 42690 24836 42702
rect 24332 42642 24612 42644
rect 24332 42590 24334 42642
rect 24386 42590 24612 42642
rect 24332 42588 24612 42590
rect 24948 42644 25004 42654
rect 24332 41972 24388 42588
rect 24948 42586 25004 42588
rect 24948 42534 24950 42586
rect 25002 42534 25004 42586
rect 24948 42522 25004 42534
rect 24332 41906 24388 41916
rect 24556 41748 24612 41758
rect 24108 40964 24164 40974
rect 24108 40870 24164 40908
rect 24220 40740 24276 41020
rect 23884 40562 23940 40572
rect 24108 40684 24276 40740
rect 24444 41186 24500 41198
rect 24444 41134 24446 41186
rect 24498 41134 24500 41186
rect 24108 40570 24164 40684
rect 24108 40518 24110 40570
rect 24162 40518 24164 40570
rect 24108 40506 24164 40518
rect 24332 40516 24388 40526
rect 24332 40429 24388 40460
rect 23436 40404 23492 40414
rect 23996 40404 24052 40414
rect 23324 40348 23436 40404
rect 23324 39618 23380 40348
rect 23436 40310 23492 40348
rect 23884 40402 24052 40404
rect 23884 40350 23998 40402
rect 24050 40350 24052 40402
rect 24332 40377 24334 40429
rect 24386 40377 24388 40429
rect 24332 40365 24388 40377
rect 24444 40404 24500 41134
rect 23884 40348 24052 40350
rect 23324 39566 23326 39618
rect 23378 39566 23380 39618
rect 23324 39554 23380 39566
rect 22092 38782 22094 38834
rect 22146 38782 22148 38834
rect 22092 38770 22148 38782
rect 22316 38849 22372 38861
rect 22316 38797 22318 38849
rect 22370 38797 22372 38849
rect 22316 38724 22372 38797
rect 22316 38658 22372 38668
rect 22428 38836 22596 38892
rect 22932 38892 22988 38902
rect 22932 38890 23044 38892
rect 22932 38838 22934 38890
rect 22986 38838 23044 38890
rect 22428 38722 22484 38836
rect 22932 38826 23044 38838
rect 22764 38724 22820 38734
rect 22428 38670 22430 38722
rect 22482 38670 22484 38722
rect 22428 38658 22484 38670
rect 22540 38722 22820 38724
rect 22540 38670 22766 38722
rect 22818 38670 22820 38722
rect 22540 38668 22820 38670
rect 22316 38500 22372 38510
rect 22204 38276 22260 38286
rect 21980 37998 21982 38050
rect 22034 37998 22036 38050
rect 21980 37940 22036 37998
rect 21980 36596 22036 37884
rect 22092 38052 22148 38062
rect 22092 36932 22148 37996
rect 22204 37268 22260 38220
rect 22316 38052 22372 38444
rect 22316 37958 22372 37996
rect 22204 37044 22260 37212
rect 22316 37268 22372 37278
rect 22540 37268 22596 38668
rect 22764 38658 22820 38668
rect 22988 38668 23044 38826
rect 23100 38834 23156 39004
rect 23436 39508 23492 39518
rect 23100 38782 23102 38834
rect 23154 38782 23156 38834
rect 23100 38770 23156 38782
rect 23324 38836 23380 38846
rect 22988 38612 23268 38668
rect 23212 38218 23268 38612
rect 23212 38166 23214 38218
rect 23266 38166 23268 38218
rect 23324 38276 23380 38780
rect 23436 38668 23492 39452
rect 23884 38849 23940 40348
rect 23996 40338 24052 40348
rect 24444 40338 24500 40348
rect 24556 40740 24612 41692
rect 24556 40402 24612 40684
rect 24556 40350 24558 40402
rect 24610 40350 24612 40402
rect 24556 40338 24612 40350
rect 24668 40516 24724 40526
rect 24668 39844 24724 40460
rect 24444 39788 24724 39844
rect 24948 40404 25004 40414
rect 24948 39842 25004 40348
rect 24948 39790 24950 39842
rect 25002 39790 25004 39842
rect 24276 39732 24332 39742
rect 23884 38797 23886 38849
rect 23938 38797 23940 38849
rect 23772 38724 23828 38734
rect 23436 38612 23604 38668
rect 23772 38630 23828 38668
rect 23324 38210 23380 38220
rect 23212 38154 23268 38166
rect 23324 38052 23380 38062
rect 23324 38050 23492 38052
rect 23324 37998 23326 38050
rect 23378 37998 23492 38050
rect 23324 37996 23492 37998
rect 23324 37986 23380 37996
rect 22316 37266 22596 37268
rect 22316 37214 22318 37266
rect 22370 37214 22596 37266
rect 22316 37212 22596 37214
rect 22316 37202 22372 37212
rect 22204 36988 22596 37044
rect 22092 36876 22372 36932
rect 22148 36596 22204 36606
rect 21980 36594 22204 36596
rect 21980 36542 22150 36594
rect 22202 36542 22204 36594
rect 21980 36540 22204 36542
rect 21980 35140 22036 36540
rect 22148 36530 22204 36540
rect 22316 35598 22372 36876
rect 22540 36650 22596 36988
rect 23436 36718 23492 37996
rect 22540 36598 22542 36650
rect 22594 36598 22596 36650
rect 22540 36586 22596 36598
rect 22652 36708 22708 36718
rect 22652 36482 22708 36652
rect 23380 36706 23492 36718
rect 23380 36654 23382 36706
rect 23434 36654 23492 36706
rect 23380 36652 23492 36654
rect 23380 36642 23436 36652
rect 22652 36430 22654 36482
rect 22706 36430 22708 36482
rect 22652 36418 22708 36430
rect 22876 36482 22932 36494
rect 22876 36430 22878 36482
rect 22930 36430 22932 36482
rect 22764 35700 22820 35710
rect 22540 35698 22820 35700
rect 22540 35646 22766 35698
rect 22818 35646 22820 35698
rect 22540 35644 22820 35646
rect 22316 35586 22428 35598
rect 22316 35534 22374 35586
rect 22426 35534 22428 35586
rect 22316 35476 22428 35534
rect 22204 35420 22428 35476
rect 22204 35252 22260 35420
rect 22540 35252 22596 35644
rect 22764 35634 22820 35644
rect 22876 35700 22932 36430
rect 22876 35364 22932 35644
rect 23436 35698 23492 35710
rect 23436 35646 23438 35698
rect 23490 35646 23492 35698
rect 23100 35588 23156 35598
rect 23100 35586 23380 35588
rect 23100 35534 23102 35586
rect 23154 35534 23380 35586
rect 23100 35532 23380 35534
rect 23100 35522 23156 35532
rect 22876 35298 22932 35308
rect 23212 35364 23268 35374
rect 22204 35186 22260 35196
rect 22316 35196 22596 35252
rect 21980 35074 22036 35084
rect 21756 34244 21812 34636
rect 21756 34188 22260 34244
rect 21644 34078 21646 34130
rect 21698 34078 21700 34130
rect 22204 34157 22260 34188
rect 22204 34105 22206 34157
rect 22258 34105 22260 34157
rect 22204 34093 22260 34105
rect 21644 34066 21700 34078
rect 21532 33506 21588 33516
rect 21644 33908 21700 33918
rect 21644 32564 21700 33852
rect 22316 33582 22372 35196
rect 23212 33906 23268 35308
rect 23324 35028 23380 35532
rect 23436 35364 23492 35646
rect 23436 35298 23492 35308
rect 23436 35028 23492 35038
rect 23324 35026 23492 35028
rect 23324 34974 23438 35026
rect 23490 34974 23492 35026
rect 23324 34972 23492 34974
rect 23436 34962 23492 34972
rect 23212 33854 23214 33906
rect 23266 33854 23268 33906
rect 23212 33796 23268 33854
rect 22764 33740 23268 33796
rect 22316 33570 22428 33582
rect 22316 33518 22374 33570
rect 22426 33518 22428 33570
rect 22316 33516 22428 33518
rect 22372 33506 22428 33516
rect 22652 33572 22708 33582
rect 22092 33348 22148 33358
rect 22092 33346 22372 33348
rect 22092 33294 22094 33346
rect 22146 33294 22372 33346
rect 22092 33292 22372 33294
rect 22092 33282 22148 33292
rect 21756 33124 21812 33134
rect 21756 33030 21812 33068
rect 21756 32564 21812 32574
rect 21644 32562 21812 32564
rect 21644 32510 21758 32562
rect 21810 32510 21812 32562
rect 21644 32508 21812 32510
rect 21756 32452 21812 32508
rect 21756 32396 22260 32452
rect 21196 32340 21252 32350
rect 21084 32338 21252 32340
rect 21084 32286 21198 32338
rect 21250 32286 21252 32338
rect 21084 32284 21252 32286
rect 21196 31220 21252 32284
rect 21532 32116 21588 32126
rect 21420 31892 21476 31902
rect 21420 31798 21476 31836
rect 21308 31780 21364 31790
rect 21308 31444 21364 31724
rect 21308 31388 21476 31444
rect 21196 31154 21252 31164
rect 20916 31052 21028 31108
rect 20860 31050 20916 31052
rect 20860 30998 20862 31050
rect 20914 30998 20916 31050
rect 20860 30986 20916 30998
rect 21140 30996 21196 31006
rect 21140 30902 21196 30940
rect 20748 30158 20750 30210
rect 20802 30158 20804 30210
rect 20748 30146 20804 30158
rect 21196 30212 21252 30222
rect 21420 30182 21476 31388
rect 21084 29540 21140 29550
rect 21084 29470 21140 29484
rect 21084 29418 21086 29470
rect 21138 29418 21140 29470
rect 21084 29406 21140 29418
rect 21196 29428 21252 30156
rect 21308 30154 21364 30166
rect 21308 30102 21310 30154
rect 21362 30102 21364 30154
rect 21420 30130 21422 30182
rect 21474 30130 21476 30182
rect 21420 30118 21476 30130
rect 21308 29652 21364 30102
rect 21532 29988 21588 32060
rect 21980 31778 22036 31790
rect 21812 31722 21868 31734
rect 21812 31670 21814 31722
rect 21866 31670 21868 31722
rect 21812 31556 21868 31670
rect 21812 31490 21868 31500
rect 21980 31726 21982 31778
rect 22034 31726 22036 31778
rect 21868 30770 21924 30782
rect 21868 30718 21870 30770
rect 21922 30718 21924 30770
rect 21868 30324 21924 30718
rect 21980 30436 22036 31726
rect 22092 31778 22148 31790
rect 22092 31726 22094 31778
rect 22146 31726 22148 31778
rect 22092 31668 22148 31726
rect 22092 31602 22148 31612
rect 22204 31444 22260 32396
rect 22316 32004 22372 33292
rect 22652 33318 22708 33516
rect 22652 33266 22654 33318
rect 22706 33266 22708 33318
rect 22652 33254 22708 33266
rect 22540 33124 22596 33134
rect 22540 32562 22596 33068
rect 22540 32510 22542 32562
rect 22594 32510 22596 32562
rect 22540 32498 22596 32510
rect 22316 31938 22372 31948
rect 22652 32116 22708 32126
rect 22484 31780 22540 31790
rect 22484 31610 22540 31724
rect 22652 31778 22708 32060
rect 22652 31726 22654 31778
rect 22706 31726 22708 31778
rect 22652 31714 22708 31726
rect 22484 31558 22486 31610
rect 22538 31558 22540 31610
rect 22484 31546 22540 31558
rect 22764 31444 22820 33740
rect 22876 33572 22932 33582
rect 22876 33318 22932 33516
rect 22876 33266 22878 33318
rect 22930 33266 22932 33318
rect 23212 33348 23268 33358
rect 22876 33254 22932 33266
rect 23100 33290 23156 33302
rect 23100 33238 23102 33290
rect 23154 33238 23156 33290
rect 23212 33259 23214 33292
rect 23266 33259 23268 33292
rect 23212 33247 23268 33259
rect 23100 32788 23156 33238
rect 23548 33012 23604 38612
rect 23884 38276 23940 38797
rect 23996 39730 24332 39732
rect 23996 39678 24278 39730
rect 24330 39678 24332 39730
rect 23996 39676 24332 39678
rect 23996 38500 24052 39676
rect 24276 39666 24332 39676
rect 24444 39618 24500 39788
rect 24948 39778 25004 39790
rect 24668 39620 24724 39630
rect 24444 39566 24446 39618
rect 24498 39566 24500 39618
rect 24220 38836 24276 38846
rect 24444 38836 24500 39566
rect 24220 38834 24500 38836
rect 24220 38782 24222 38834
rect 24274 38782 24500 38834
rect 24220 38780 24500 38782
rect 24556 39618 24724 39620
rect 24556 39566 24670 39618
rect 24722 39566 24724 39618
rect 24556 39564 24724 39566
rect 24220 38770 24276 38780
rect 24556 38668 24612 39564
rect 24668 39554 24724 39564
rect 25116 39172 25172 43596
rect 25228 43538 25284 44268
rect 25228 43486 25230 43538
rect 25282 43486 25284 43538
rect 25228 43474 25284 43486
rect 25452 42980 25508 42990
rect 25452 42886 25508 42924
rect 25788 42756 25844 42766
rect 25788 42662 25844 42700
rect 25900 42754 25956 45054
rect 26236 45108 26292 45118
rect 26012 43426 26068 43438
rect 26012 43374 26014 43426
rect 26066 43374 26068 43426
rect 26012 42980 26068 43374
rect 26012 42914 26068 42924
rect 25900 42702 25902 42754
rect 25954 42702 25956 42754
rect 25228 41972 25284 41982
rect 25228 41878 25284 41916
rect 25900 41972 25956 42702
rect 25900 41906 25956 41916
rect 25396 41748 25452 41758
rect 25396 41654 25452 41692
rect 26236 41524 26292 45052
rect 26684 45106 26740 45612
rect 27356 45668 27412 45678
rect 27972 45668 28028 45678
rect 27356 45574 27412 45612
rect 27916 45666 28028 45668
rect 27916 45614 27974 45666
rect 28026 45614 28028 45666
rect 27916 45602 28028 45614
rect 26684 45054 26686 45106
rect 26738 45054 26740 45106
rect 26684 45042 26740 45054
rect 27692 44266 27748 44278
rect 27692 44214 27694 44266
rect 27746 44214 27748 44266
rect 27412 44100 27468 44110
rect 27692 44100 27748 44214
rect 27412 44098 27524 44100
rect 27412 44046 27414 44098
rect 27466 44046 27524 44098
rect 27412 44034 27524 44046
rect 27692 44034 27748 44044
rect 27804 44266 27860 44278
rect 27804 44214 27806 44266
rect 27858 44214 27860 44266
rect 27468 43316 27524 44034
rect 27804 43428 27860 44214
rect 27916 44100 27972 45602
rect 28252 44996 28308 45006
rect 28028 44772 28084 44782
rect 28028 44294 28084 44716
rect 28028 44242 28030 44294
rect 28082 44242 28084 44294
rect 28028 44230 28084 44242
rect 28252 44324 28308 44940
rect 28252 44242 28254 44268
rect 28306 44242 28308 44268
rect 28252 44230 28308 44242
rect 27916 44034 27972 44044
rect 28028 43988 28084 43998
rect 27916 43428 27972 43438
rect 27468 43250 27524 43260
rect 27692 43426 27972 43428
rect 27692 43374 27918 43426
rect 27970 43374 27972 43426
rect 27692 43372 27972 43374
rect 27412 42756 27468 42766
rect 27412 42662 27468 42700
rect 27692 42756 27748 43372
rect 27916 43362 27972 43372
rect 27692 42674 27694 42700
rect 27746 42674 27748 42700
rect 27692 42662 27748 42674
rect 27916 43204 27972 43214
rect 27916 42726 27972 43148
rect 27916 42674 27918 42726
rect 27970 42674 27972 42726
rect 27916 42662 27972 42674
rect 26460 41972 26516 41982
rect 26292 41468 26404 41524
rect 26236 41458 26292 41468
rect 25228 41186 25284 41198
rect 25228 41134 25230 41186
rect 25282 41134 25284 41186
rect 25228 39844 25284 41134
rect 25900 40964 25956 40974
rect 25564 40628 25620 40638
rect 25452 40404 25508 40414
rect 25452 40310 25508 40348
rect 25452 39844 25508 39854
rect 25228 39842 25508 39844
rect 25228 39790 25454 39842
rect 25506 39790 25508 39842
rect 25228 39788 25508 39790
rect 25452 39778 25508 39788
rect 25116 39060 25172 39116
rect 24892 39004 25172 39060
rect 25452 39060 25508 39070
rect 25564 39060 25620 40572
rect 25788 40570 25844 40582
rect 25788 40518 25790 40570
rect 25842 40518 25844 40570
rect 25452 39058 25620 39060
rect 25452 39006 25454 39058
rect 25506 39006 25620 39058
rect 25452 39004 25620 39006
rect 25676 40441 25732 40453
rect 25676 40389 25678 40441
rect 25730 40389 25732 40441
rect 24724 38724 24780 38734
rect 23996 38434 24052 38444
rect 24108 38612 24612 38668
rect 24668 38722 24780 38724
rect 24668 38670 24726 38722
rect 24778 38670 24780 38722
rect 24668 38658 24780 38670
rect 24108 38276 24164 38612
rect 23884 38220 24164 38276
rect 23660 38052 23716 38062
rect 23884 38052 23940 38220
rect 24108 38162 24164 38220
rect 24108 38110 24110 38162
rect 24162 38110 24164 38162
rect 24108 38098 24164 38110
rect 24444 38388 24500 38398
rect 23660 38050 23940 38052
rect 23660 37998 23662 38050
rect 23714 37998 23940 38050
rect 23660 37996 23940 37998
rect 23996 38050 24052 38062
rect 23996 37998 23998 38050
rect 24050 37998 24052 38050
rect 23660 37986 23716 37996
rect 23996 37828 24052 37998
rect 24444 38011 24500 38332
rect 24444 37959 24446 38011
rect 24498 37959 24500 38011
rect 23996 37762 24052 37772
rect 24220 37828 24276 37838
rect 24220 37380 24276 37772
rect 24108 37378 24276 37380
rect 24108 37326 24222 37378
rect 24274 37326 24276 37378
rect 24108 37324 24276 37326
rect 23940 37044 23996 37054
rect 23940 36538 23996 36988
rect 23660 36484 23716 36494
rect 23940 36486 23942 36538
rect 23994 36486 23996 36538
rect 23940 36474 23996 36486
rect 24108 36482 24164 37324
rect 24220 37314 24276 37324
rect 24444 37044 24500 37959
rect 24444 36978 24500 36988
rect 24668 38050 24724 38658
rect 24668 37998 24670 38050
rect 24722 37998 24724 38050
rect 24668 37940 24724 37998
rect 24668 36932 24724 37884
rect 24668 36866 24724 36876
rect 24892 36708 24948 39004
rect 25452 38994 25508 39004
rect 25116 38836 25172 38846
rect 25116 38742 25172 38780
rect 25676 38724 25732 40389
rect 25788 39618 25844 40518
rect 25788 39566 25790 39618
rect 25842 39566 25844 39618
rect 25788 39554 25844 39566
rect 25788 38836 25844 38846
rect 25788 38742 25844 38780
rect 25900 38668 25956 40908
rect 26348 40740 26404 41468
rect 26460 40964 26516 41916
rect 27916 41748 27972 41758
rect 27916 41188 27972 41692
rect 27916 41106 27918 41132
rect 27970 41106 27972 41132
rect 27916 41094 27972 41106
rect 26460 40898 26516 40908
rect 27132 41074 27188 41086
rect 27132 41022 27134 41074
rect 27186 41022 27188 41074
rect 26348 40684 26516 40740
rect 26124 40628 26180 40638
rect 26124 40404 26180 40572
rect 26124 40402 26404 40404
rect 26124 40350 26126 40402
rect 26178 40350 26404 40402
rect 26124 40348 26404 40350
rect 26124 40338 26180 40348
rect 26348 39742 26404 40348
rect 26460 40180 26516 40684
rect 26628 40570 26684 40582
rect 26628 40518 26630 40570
rect 26682 40518 26684 40570
rect 26628 40404 26684 40518
rect 26628 40338 26684 40348
rect 26796 40404 26852 40414
rect 27020 40404 27076 40414
rect 27132 40404 27188 41022
rect 27636 41074 27692 41086
rect 27636 41022 27638 41074
rect 27690 41022 27692 41074
rect 27636 40852 27692 41022
rect 27636 40786 27692 40796
rect 28028 40628 28084 43932
rect 28364 43662 28420 46060
rect 28644 45892 28700 45902
rect 29148 45892 29204 45902
rect 29260 45892 29316 47180
rect 28644 45890 29316 45892
rect 28644 45838 28646 45890
rect 28698 45838 29150 45890
rect 29202 45838 29316 45890
rect 28644 45836 29316 45838
rect 29372 45892 29428 47292
rect 29484 47282 29540 47292
rect 30212 47236 30268 47246
rect 30212 47142 30268 47180
rect 30268 46674 30324 46686
rect 30268 46622 30270 46674
rect 30322 46622 30324 46674
rect 29484 46562 29540 46574
rect 29484 46510 29486 46562
rect 29538 46510 29540 46562
rect 29484 46004 29540 46510
rect 29596 46004 29652 46014
rect 29484 46002 29652 46004
rect 29484 45950 29598 46002
rect 29650 45950 29652 46002
rect 29484 45948 29652 45950
rect 29596 45938 29652 45948
rect 30044 45892 30100 45902
rect 29372 45860 29484 45892
rect 29372 45836 29430 45860
rect 28644 45826 28700 45836
rect 28588 44994 28644 45006
rect 28588 44942 28590 44994
rect 28642 44942 28644 44994
rect 28588 44772 28644 44942
rect 28644 44716 28756 44772
rect 28588 44706 28644 44716
rect 28532 44436 28588 44446
rect 28476 44434 28588 44436
rect 28476 44382 28534 44434
rect 28586 44382 28588 44434
rect 28476 44370 28588 44382
rect 28476 44212 28532 44370
rect 28476 44156 28588 44212
rect 28364 43650 28476 43662
rect 28364 43598 28422 43650
rect 28474 43598 28476 43650
rect 28364 43596 28476 43598
rect 28532 43652 28588 44156
rect 28532 43596 28644 43652
rect 28420 43586 28476 43596
rect 28588 43540 28644 43596
rect 28700 43594 28756 44716
rect 29036 44324 29092 44334
rect 29036 44230 29092 44268
rect 28700 43542 28702 43594
rect 28754 43542 28756 43594
rect 29036 44100 29092 44110
rect 28700 43530 28756 43542
rect 28924 43566 28980 43578
rect 28588 43474 28644 43484
rect 28924 43514 28926 43566
rect 28978 43514 28980 43566
rect 28140 43428 28196 43438
rect 28140 42726 28196 43372
rect 28812 43428 28868 43438
rect 28140 42674 28142 42726
rect 28194 42674 28196 42726
rect 28140 42662 28196 42674
rect 28252 43316 28308 43326
rect 28252 42698 28308 43260
rect 28252 42646 28254 42698
rect 28306 42646 28308 42698
rect 28252 41412 28308 42646
rect 28700 43204 28756 43214
rect 28476 41997 28532 42009
rect 28476 41945 28478 41997
rect 28530 41945 28532 41997
rect 28476 41860 28532 41945
rect 28476 41794 28532 41804
rect 28252 41346 28308 41356
rect 28140 41130 28196 41142
rect 28140 41078 28142 41130
rect 28194 41078 28196 41130
rect 28140 41076 28196 41078
rect 28140 41010 28196 41020
rect 28364 41130 28420 41142
rect 28364 41078 28366 41130
rect 28418 41078 28420 41130
rect 28028 40562 28084 40572
rect 28252 40628 28308 40638
rect 28140 40516 28196 40526
rect 28140 40422 28196 40460
rect 26796 40402 27188 40404
rect 26796 40350 26798 40402
rect 26850 40350 27022 40402
rect 27074 40350 27188 40402
rect 26796 40348 27188 40350
rect 27692 40404 27748 40414
rect 26796 40338 26852 40348
rect 27020 40338 27076 40348
rect 27692 40180 27748 40348
rect 27896 40404 27952 40414
rect 27896 40402 28084 40404
rect 27896 40350 27898 40402
rect 27950 40350 28084 40402
rect 27896 40348 28084 40350
rect 27896 40338 27952 40348
rect 26460 40124 26628 40180
rect 27692 40124 27916 40180
rect 26348 39730 26460 39742
rect 26348 39678 26406 39730
rect 26458 39678 26460 39730
rect 26348 39676 26460 39678
rect 26404 39666 26460 39676
rect 26124 39060 26180 39070
rect 26124 38966 26180 39004
rect 26572 38892 26628 40124
rect 26460 38836 26628 38892
rect 26796 40068 26852 40078
rect 26460 38834 26516 38836
rect 26460 38782 26462 38834
rect 26514 38782 26516 38834
rect 26460 38770 26516 38782
rect 26684 38834 26740 38846
rect 26684 38782 26686 38834
rect 26738 38782 26740 38834
rect 25676 38658 25732 38668
rect 25788 38612 25956 38668
rect 26572 38724 26628 38734
rect 25004 38500 25060 38510
rect 25004 38050 25060 38444
rect 25004 37998 25006 38050
rect 25058 37998 25060 38050
rect 25004 37492 25060 37998
rect 25788 38050 25844 38612
rect 25788 37998 25790 38050
rect 25842 37998 25844 38050
rect 25788 37986 25844 37998
rect 26012 38388 26068 38398
rect 25004 37426 25060 37436
rect 25732 37716 25788 37726
rect 25732 37492 25788 37660
rect 25732 37398 25788 37436
rect 26012 37266 26068 38332
rect 26572 38162 26628 38668
rect 26572 38110 26574 38162
rect 26626 38110 26628 38162
rect 26572 38098 26628 38110
rect 26684 37604 26740 38782
rect 26684 37538 26740 37548
rect 26796 37380 26852 40012
rect 27692 39956 27748 39966
rect 27580 39844 27636 39854
rect 27580 39396 27636 39788
rect 27692 39618 27748 39900
rect 27692 39566 27694 39618
rect 27746 39566 27748 39618
rect 27860 39674 27916 40124
rect 27860 39622 27862 39674
rect 27914 39622 27916 39674
rect 27860 39610 27916 39622
rect 27692 39554 27748 39566
rect 28028 39506 28084 40348
rect 28140 39620 28196 39630
rect 28252 39620 28308 40572
rect 28364 40180 28420 41078
rect 28476 41130 28532 41142
rect 28476 41078 28478 41130
rect 28530 41078 28532 41130
rect 28476 40740 28532 41078
rect 28476 40402 28532 40684
rect 28700 40740 28756 43148
rect 28700 40674 28756 40684
rect 28700 40404 28756 40414
rect 28476 40350 28478 40402
rect 28530 40350 28532 40402
rect 28476 40338 28532 40350
rect 28588 40402 28756 40404
rect 28588 40350 28702 40402
rect 28754 40350 28756 40402
rect 28588 40348 28756 40350
rect 28588 40180 28644 40348
rect 28700 40338 28756 40348
rect 28364 40124 28644 40180
rect 28476 39844 28532 40124
rect 28476 39778 28532 39788
rect 28140 39618 28308 39620
rect 28140 39566 28142 39618
rect 28194 39566 28308 39618
rect 28140 39564 28308 39566
rect 28420 39620 28476 39630
rect 28140 39554 28196 39564
rect 28420 39526 28476 39564
rect 28028 39454 28030 39506
rect 28082 39454 28084 39506
rect 27580 39340 27748 39396
rect 26964 38836 27020 38846
rect 27244 38836 27300 38846
rect 26964 38834 27300 38836
rect 26964 38782 26966 38834
rect 27018 38782 27246 38834
rect 27298 38782 27300 38834
rect 26964 38780 27300 38782
rect 26964 38770 27020 38780
rect 27244 38770 27300 38780
rect 27580 38724 27636 38762
rect 27580 38658 27636 38668
rect 26012 37214 26014 37266
rect 26066 37214 26068 37266
rect 26012 37202 26068 37214
rect 26684 37324 26852 37380
rect 27132 37604 27188 37614
rect 27132 37378 27188 37548
rect 27692 37380 27748 39340
rect 28028 38668 28084 39454
rect 28364 39284 28420 39294
rect 28028 38612 28196 38668
rect 27132 37326 27134 37378
rect 27186 37326 27188 37378
rect 23660 35476 23716 36428
rect 24108 36430 24110 36482
rect 24162 36430 24164 36482
rect 24108 36418 24164 36430
rect 24220 36652 24948 36708
rect 23772 36370 23828 36382
rect 23772 36318 23774 36370
rect 23826 36318 23828 36370
rect 23772 36148 23828 36318
rect 23772 36082 23828 36092
rect 24220 35934 24276 36652
rect 24164 35924 24276 35934
rect 23660 35410 23716 35420
rect 24108 35922 24276 35924
rect 24108 35870 24166 35922
rect 24218 35870 24276 35922
rect 24108 35868 24276 35870
rect 24332 36482 24388 36494
rect 24332 36430 24334 36482
rect 24386 36430 24388 36482
rect 24108 35858 24220 35868
rect 23884 33684 23940 33694
rect 23772 33572 23828 33582
rect 23772 33458 23828 33516
rect 23772 33406 23774 33458
rect 23826 33406 23828 33458
rect 23772 33236 23828 33406
rect 23772 33170 23828 33180
rect 23548 32956 23828 33012
rect 23100 32722 23156 32732
rect 23660 32788 23716 32798
rect 23212 32116 23268 32126
rect 22932 32004 22988 32014
rect 22932 31910 22988 31948
rect 22204 31388 22820 31444
rect 22876 31780 22932 31790
rect 22282 31031 22338 31043
rect 22282 30979 22284 31031
rect 22336 30996 22338 31031
rect 22428 30996 22484 31006
rect 22336 30979 22372 30996
rect 22282 30940 22372 30979
rect 22148 30436 22204 30446
rect 21980 30434 22204 30436
rect 21980 30382 22150 30434
rect 22202 30382 22204 30434
rect 21980 30380 22204 30382
rect 22148 30370 22204 30380
rect 21756 30268 21924 30324
rect 22316 30324 22372 30940
rect 21756 30187 21812 30268
rect 22316 30258 22372 30268
rect 22428 30212 22484 30940
rect 22540 30994 22596 31006
rect 22540 30942 22542 30994
rect 22594 30942 22596 30994
rect 22540 30548 22596 30942
rect 22540 30482 22596 30492
rect 22652 30212 22708 31388
rect 22764 31108 22820 31118
rect 22764 30994 22820 31052
rect 22764 30942 22766 30994
rect 22818 30942 22820 30994
rect 22764 30930 22820 30942
rect 22876 30660 22932 31724
rect 23212 31750 23268 32060
rect 23212 31698 23214 31750
rect 23266 31698 23268 31750
rect 23212 31686 23268 31698
rect 23436 31780 23492 31790
rect 23436 31698 23438 31724
rect 23490 31698 23492 31724
rect 23436 31686 23492 31698
rect 23660 31750 23716 32732
rect 23660 31698 23662 31750
rect 23714 31698 23716 31750
rect 23660 31686 23716 31698
rect 23772 31743 23828 32956
rect 23772 31691 23774 31743
rect 23826 31691 23828 31743
rect 22988 30994 23044 31006
rect 23772 30996 23828 31691
rect 22988 30942 22990 30994
rect 23042 30942 23044 30994
rect 22988 30884 23044 30942
rect 22988 30818 23044 30828
rect 23660 30940 23828 30996
rect 23884 31780 23940 33628
rect 24108 33348 24164 35858
rect 24220 35364 24276 35374
rect 24332 35364 24388 36430
rect 25116 36482 25172 36494
rect 25116 36430 25118 36482
rect 25170 36430 25172 36482
rect 25116 35924 25172 36430
rect 26124 36036 26180 36046
rect 25116 35858 25172 35868
rect 25788 35924 25844 35934
rect 25788 35830 25844 35868
rect 25396 35700 25452 35710
rect 25396 35606 25452 35644
rect 26124 35698 26180 35980
rect 26124 35646 26126 35698
rect 26178 35646 26180 35698
rect 26124 35634 26180 35646
rect 24612 35586 24668 35598
rect 24612 35534 24614 35586
rect 24666 35534 24668 35586
rect 24612 35476 24668 35534
rect 24612 35410 24668 35420
rect 25564 35588 25620 35598
rect 24276 35308 24388 35364
rect 24220 34914 24276 35308
rect 24220 34862 24222 34914
rect 24274 34862 24276 34914
rect 24220 34850 24276 34862
rect 24444 34858 24500 34870
rect 24444 34806 24446 34858
rect 24498 34806 24500 34858
rect 24444 34132 24500 34806
rect 24444 34066 24500 34076
rect 24556 34858 24612 34870
rect 24556 34806 24558 34858
rect 24610 34806 24612 34858
rect 24108 33282 24164 33292
rect 24556 32788 24612 34806
rect 24780 34858 24836 34870
rect 24780 34806 24782 34858
rect 24834 34806 24836 34858
rect 24780 33684 24836 34806
rect 24780 33618 24836 33628
rect 25004 34858 25060 34870
rect 25004 34806 25006 34858
rect 25058 34806 25060 34858
rect 25004 33684 25060 34806
rect 25284 34804 25340 34814
rect 25116 34802 25340 34804
rect 25116 34750 25286 34802
rect 25338 34750 25340 34802
rect 25116 34748 25340 34750
rect 25116 34130 25172 34748
rect 25284 34738 25340 34748
rect 25564 34692 25620 35532
rect 26516 35586 26572 35598
rect 26516 35534 26518 35586
rect 26570 35534 26572 35586
rect 26516 35476 26572 35534
rect 26516 35410 26572 35420
rect 25564 34626 25620 34636
rect 25788 34914 25844 34926
rect 25788 34862 25790 34914
rect 25842 34862 25844 34914
rect 25116 34078 25118 34130
rect 25170 34078 25172 34130
rect 25116 34066 25172 34078
rect 25452 33908 25508 33918
rect 25452 33906 25732 33908
rect 25452 33854 25454 33906
rect 25506 33854 25732 33906
rect 25452 33852 25732 33854
rect 25452 33842 25508 33852
rect 25004 33618 25060 33628
rect 25676 33458 25732 33852
rect 25676 33406 25678 33458
rect 25730 33406 25732 33458
rect 25676 33394 25732 33406
rect 25788 33348 25844 34862
rect 26572 34914 26628 34926
rect 26572 34862 26574 34914
rect 26626 34862 26628 34914
rect 26460 34580 26516 34590
rect 26460 34142 26516 34524
rect 26572 34356 26628 34862
rect 26572 34290 26628 34300
rect 26460 34132 26572 34142
rect 26460 34076 26516 34132
rect 26516 34038 26572 34076
rect 26068 34020 26124 34030
rect 25788 33282 25844 33292
rect 26012 34018 26124 34020
rect 26012 33966 26070 34018
rect 26122 33966 26124 34018
rect 26012 33954 26124 33966
rect 24556 32722 24612 32732
rect 25116 33124 25172 33134
rect 26012 33124 26068 33954
rect 26460 33348 26516 33358
rect 26460 33254 26516 33292
rect 24444 32450 24500 32462
rect 24444 32398 24446 32450
rect 24498 32398 24500 32450
rect 24444 32116 24500 32398
rect 24444 32050 24500 32060
rect 23268 30770 23324 30782
rect 23268 30718 23270 30770
rect 23322 30718 23324 30770
rect 22876 30604 23044 30660
rect 22764 30212 22820 30222
rect 21700 30175 21812 30187
rect 21700 30123 21702 30175
rect 21754 30128 21812 30175
rect 21924 30184 21980 30187
rect 21924 30175 22036 30184
rect 21754 30123 21756 30128
rect 21700 30111 21756 30123
rect 21924 30123 21926 30175
rect 21978 30123 22036 30175
rect 22428 30156 22596 30212
rect 22652 30210 22820 30212
rect 22652 30158 22766 30210
rect 22818 30158 22820 30210
rect 22652 30156 22820 30158
rect 21924 30111 22036 30123
rect 21980 30100 22036 30111
rect 21980 30044 22484 30100
rect 21868 29988 21924 29998
rect 21532 29932 21700 29988
rect 21308 29596 21476 29652
rect 21308 29428 21364 29438
rect 21196 29426 21364 29428
rect 21196 29374 21310 29426
rect 21362 29374 21364 29426
rect 21196 29372 21364 29374
rect 20972 29316 21028 29326
rect 20972 29222 21028 29260
rect 21308 28980 21364 29372
rect 21308 28914 21364 28924
rect 21420 29428 21476 29596
rect 21420 28756 21476 29372
rect 21420 28690 21476 28700
rect 21532 28868 21588 28878
rect 21252 28588 21308 28598
rect 19628 27902 19684 27916
rect 18956 26852 19124 26908
rect 19180 27858 19236 27870
rect 19180 27806 19182 27858
rect 19234 27806 19236 27858
rect 19628 27850 19630 27902
rect 19682 27850 19684 27902
rect 19628 27838 19684 27850
rect 19964 27860 20020 27870
rect 19180 26852 19236 27806
rect 19964 27766 20020 27804
rect 20524 27858 20580 27916
rect 21196 28586 21308 28588
rect 21196 28534 21254 28586
rect 21306 28534 21308 28586
rect 21196 28522 21308 28534
rect 21420 28588 21476 28598
rect 21532 28588 21588 28812
rect 21420 28586 21588 28588
rect 21420 28534 21422 28586
rect 21474 28534 21588 28586
rect 21644 28614 21700 29932
rect 21868 29428 21924 29932
rect 22204 29465 22260 29477
rect 21980 29428 22036 29438
rect 21868 29426 22036 29428
rect 21868 29374 21982 29426
rect 22034 29374 22036 29426
rect 21868 29372 22036 29374
rect 21980 29362 22036 29372
rect 22204 29413 22206 29465
rect 22258 29413 22260 29465
rect 21644 28562 21646 28614
rect 21698 28562 21700 28614
rect 21644 28550 21700 28562
rect 21868 29092 21924 29102
rect 21868 28614 21924 29036
rect 22204 28980 22260 29413
rect 22428 29204 22484 30044
rect 22540 29764 22596 30156
rect 22764 30146 22820 30156
rect 22540 29708 22708 29764
rect 22540 29594 22596 29606
rect 22540 29542 22542 29594
rect 22594 29542 22596 29594
rect 22540 29428 22596 29542
rect 22540 29362 22596 29372
rect 22652 29426 22708 29708
rect 22652 29374 22654 29426
rect 22706 29374 22708 29426
rect 22652 29362 22708 29374
rect 22876 29428 22932 29438
rect 22876 29334 22932 29372
rect 22988 29204 23044 30604
rect 23268 30548 23324 30718
rect 23268 30482 23324 30492
rect 23548 30210 23604 30222
rect 23548 30158 23550 30210
rect 23602 30158 23604 30210
rect 23548 29652 23604 30158
rect 23660 29652 23716 30940
rect 23772 30772 23828 30782
rect 23884 30772 23940 31724
rect 24332 31890 24388 31902
rect 24332 31838 24334 31890
rect 24386 31838 24388 31890
rect 24108 30996 24164 31006
rect 24220 30996 24276 31006
rect 24332 30996 24388 31838
rect 24780 31778 24836 31790
rect 24444 31734 24500 31746
rect 24444 31682 24446 31734
rect 24498 31682 24500 31734
rect 24444 31668 24500 31682
rect 24444 31602 24500 31612
rect 24780 31726 24782 31778
rect 24834 31726 24836 31778
rect 24780 31220 24836 31726
rect 25116 31743 25172 33068
rect 25788 33068 26068 33124
rect 25340 32788 25396 32798
rect 25340 31780 25396 32732
rect 25676 32564 25732 32574
rect 25564 32562 25732 32564
rect 25564 32510 25678 32562
rect 25730 32510 25732 32562
rect 25564 32508 25732 32510
rect 25116 31691 25118 31743
rect 25170 31691 25172 31743
rect 25116 31679 25172 31691
rect 25284 31743 25396 31780
rect 25284 31691 25286 31743
rect 25338 31724 25396 31743
rect 25452 31780 25508 31790
rect 25338 31691 25340 31724
rect 25284 31679 25340 31691
rect 25452 31698 25454 31724
rect 25506 31698 25508 31724
rect 25452 31686 25508 31698
rect 25564 31668 25620 32508
rect 25676 32498 25732 32508
rect 25676 31892 25732 31902
rect 25676 31750 25732 31836
rect 25676 31698 25678 31750
rect 25730 31698 25732 31750
rect 25676 31686 25732 31698
rect 25564 31556 25620 31612
rect 25564 31500 25732 31556
rect 24780 31154 24836 31164
rect 25508 31029 25564 31041
rect 24108 30994 24388 30996
rect 24108 30942 24110 30994
rect 24162 30942 24222 30994
rect 24274 30942 24388 30994
rect 24108 30940 24388 30942
rect 24556 30996 24612 31006
rect 25508 30996 25510 31029
rect 24108 30930 24164 30940
rect 24220 30930 24276 30940
rect 24556 30902 24612 30940
rect 25452 30977 25510 30996
rect 25562 30977 25564 31029
rect 25452 30940 25564 30977
rect 23772 30770 23940 30772
rect 23772 30718 23774 30770
rect 23826 30718 23940 30770
rect 23772 30716 23940 30718
rect 24668 30884 24724 30894
rect 23772 30706 23828 30716
rect 24444 29652 24500 29662
rect 23660 29596 24108 29652
rect 23548 29586 23604 29596
rect 24052 29540 24108 29596
rect 24444 29558 24500 29596
rect 24052 29538 24164 29540
rect 24052 29486 24054 29538
rect 24106 29486 24164 29538
rect 24052 29474 24164 29486
rect 23100 29426 23156 29438
rect 23100 29374 23102 29426
rect 23154 29374 23156 29426
rect 23100 29316 23156 29374
rect 23100 29250 23156 29260
rect 22428 29148 22820 29204
rect 22316 29092 22372 29102
rect 22372 29036 22652 29092
rect 22316 29026 22372 29036
rect 21868 28562 21870 28614
rect 21922 28562 21924 28614
rect 21868 28550 21924 28562
rect 22092 28924 22260 28980
rect 21420 28532 21588 28534
rect 22092 28542 22148 28924
rect 22596 28866 22652 29036
rect 22596 28814 22598 28866
rect 22650 28814 22652 28866
rect 22596 28802 22652 28814
rect 22428 28644 22484 28654
rect 22428 28550 22484 28588
rect 21420 28522 21476 28532
rect 22092 28530 22204 28542
rect 20860 27885 20916 27898
rect 20860 27860 20862 27885
rect 20914 27860 20916 27885
rect 20524 27806 20526 27858
rect 20578 27806 20580 27858
rect 19516 27746 19572 27758
rect 19516 27694 19518 27746
rect 19570 27694 19572 27746
rect 19516 27412 19572 27694
rect 19516 27346 19572 27356
rect 19292 27076 19348 27086
rect 20132 27076 20188 27086
rect 19292 27074 20188 27076
rect 19292 27022 19294 27074
rect 19346 27022 20134 27074
rect 20186 27022 20188 27074
rect 19292 27020 20188 27022
rect 19292 27010 19348 27020
rect 20132 27010 20188 27020
rect 20412 27076 20468 27086
rect 20524 27076 20580 27806
rect 20412 27074 20580 27076
rect 20412 27022 20414 27074
rect 20466 27022 20580 27074
rect 20412 27020 20580 27022
rect 20636 27804 20860 27860
rect 20636 27074 20692 27804
rect 20860 27794 20916 27804
rect 21196 27858 21252 28522
rect 22092 28478 22150 28530
rect 22202 28478 22204 28530
rect 22092 28476 22204 28478
rect 22148 28420 22204 28476
rect 22148 28364 22640 28420
rect 21196 27806 21198 27858
rect 21250 27806 21252 27858
rect 21196 27300 21252 27806
rect 21644 27891 21700 27903
rect 21644 27860 21646 27891
rect 21698 27860 21700 27891
rect 21364 27300 21420 27310
rect 21196 27298 21420 27300
rect 21196 27246 21366 27298
rect 21418 27246 21420 27298
rect 21196 27244 21420 27246
rect 21364 27234 21420 27244
rect 20636 27022 20638 27074
rect 20690 27022 20692 27074
rect 20412 27010 20468 27020
rect 20636 27010 20692 27022
rect 21532 27074 21588 27086
rect 21532 27022 21534 27074
rect 21586 27022 21588 27074
rect 18956 26404 19012 26852
rect 18844 26348 19012 26404
rect 18284 26068 18340 26078
rect 18284 25974 18340 26012
rect 17724 25566 17726 25618
rect 17778 25566 17780 25618
rect 17724 25554 17780 25566
rect 17948 25788 18116 25844
rect 17500 24434 17556 24444
rect 17612 25172 17668 25182
rect 17612 24554 17668 25116
rect 17612 24502 17614 24554
rect 17666 24502 17668 24554
rect 17612 24052 17668 24502
rect 17724 24722 17780 24734
rect 17724 24670 17726 24722
rect 17778 24670 17780 24722
rect 17724 24276 17780 24670
rect 17724 24210 17780 24220
rect 17948 24164 18004 25788
rect 18172 24722 18228 24734
rect 18172 24670 18174 24722
rect 18226 24670 18228 24722
rect 17948 24108 18116 24164
rect 17612 23986 17668 23996
rect 17724 23938 17780 23950
rect 17388 23044 17444 23772
rect 17556 23882 17612 23894
rect 17556 23830 17558 23882
rect 17610 23830 17612 23882
rect 17556 23828 17612 23830
rect 17556 23762 17612 23772
rect 17724 23886 17726 23938
rect 17778 23886 17780 23938
rect 17612 23268 17668 23278
rect 17612 23210 17668 23212
rect 17612 23158 17614 23210
rect 17666 23158 17668 23210
rect 17612 23146 17668 23158
rect 17500 23098 17556 23110
rect 17500 23046 17502 23098
rect 17554 23046 17556 23098
rect 17500 23044 17556 23046
rect 17052 21410 17108 21420
rect 17164 22988 17556 23044
rect 17724 23044 17780 23886
rect 17948 23940 18004 23950
rect 17948 23846 18004 23884
rect 17164 20020 17220 22988
rect 17724 22978 17780 22988
rect 17612 22260 17668 22270
rect 17500 22258 17668 22260
rect 17500 22206 17614 22258
rect 17666 22206 17668 22258
rect 17500 22204 17668 22206
rect 17276 21924 17332 21934
rect 17276 21586 17332 21868
rect 17500 21700 17556 22204
rect 17612 22194 17668 22204
rect 17500 21634 17556 21644
rect 17612 21812 17668 21822
rect 17276 21534 17278 21586
rect 17330 21534 17332 21586
rect 17276 21522 17332 21534
rect 17444 21362 17500 21374
rect 17444 21310 17446 21362
rect 17498 21310 17500 21362
rect 17444 20916 17500 21310
rect 17444 20850 17500 20860
rect 17612 20802 17668 21756
rect 17612 20750 17614 20802
rect 17666 20750 17668 20802
rect 17612 20132 17668 20750
rect 17948 21474 18004 21486
rect 17948 21422 17950 21474
rect 18002 21422 18004 21474
rect 17948 20356 18004 21422
rect 17948 20290 18004 20300
rect 18060 20804 18116 24108
rect 18172 23266 18228 24670
rect 18284 24722 18340 24734
rect 18844 24724 18900 26348
rect 19068 26292 19124 26302
rect 18284 24670 18286 24722
rect 18338 24670 18340 24722
rect 18284 24164 18340 24670
rect 18732 24668 18900 24724
rect 18956 26290 19124 26292
rect 18956 26238 19070 26290
rect 19122 26238 19124 26290
rect 18956 26236 19124 26238
rect 18564 24500 18620 24510
rect 18564 24406 18620 24444
rect 18732 24164 18788 24668
rect 18284 24098 18340 24108
rect 18620 24108 18788 24164
rect 18844 24500 18900 24510
rect 18172 23214 18174 23266
rect 18226 23214 18228 23266
rect 18172 23202 18228 23214
rect 18284 23828 18340 23838
rect 18284 23278 18340 23772
rect 18284 23268 18396 23278
rect 18284 23212 18340 23268
rect 18340 23210 18396 23212
rect 18340 23158 18342 23210
rect 18394 23158 18396 23210
rect 18340 23146 18396 23158
rect 18060 20188 18116 20748
rect 17612 20066 17668 20076
rect 17836 20132 18116 20188
rect 18172 23044 18228 23054
rect 18172 22158 18228 22988
rect 18508 22370 18564 22382
rect 18508 22318 18510 22370
rect 18562 22318 18564 22370
rect 18172 22146 18284 22158
rect 18172 22094 18230 22146
rect 18282 22094 18284 22146
rect 18172 22082 18284 22094
rect 17724 20045 17780 20057
rect 17388 20020 17444 20030
rect 17164 20018 17444 20020
rect 17164 19966 17390 20018
rect 17442 19966 17444 20018
rect 17164 19964 17444 19966
rect 16940 19954 16996 19964
rect 17388 19954 17444 19964
rect 17724 19993 17726 20045
rect 17778 19993 17780 20045
rect 17612 19908 17668 19918
rect 17612 19814 17668 19852
rect 16436 19796 16492 19806
rect 14476 19742 14478 19794
rect 14530 19742 14532 19794
rect 13916 18564 13972 18844
rect 13916 18498 13972 18508
rect 13748 18398 13750 18450
rect 13802 18398 13804 18450
rect 13468 18386 13524 18396
rect 13748 18386 13804 18398
rect 14028 18452 14084 18462
rect 14476 18452 14532 19742
rect 16268 19794 16492 19796
rect 16268 19742 16438 19794
rect 16490 19742 16492 19794
rect 16268 19740 16492 19742
rect 16268 19460 16324 19740
rect 16436 19730 16492 19740
rect 16156 19404 16324 19460
rect 16716 19684 16772 19694
rect 14588 19348 14644 19358
rect 14588 19254 14644 19292
rect 15092 19236 15148 19246
rect 15092 19142 15148 19180
rect 15316 19178 15372 19190
rect 15316 19126 15318 19178
rect 15370 19126 15372 19178
rect 15316 19124 15372 19126
rect 15260 19068 15372 19124
rect 15596 19178 15652 19190
rect 15596 19126 15598 19178
rect 15650 19126 15652 19178
rect 15260 18676 15316 19068
rect 15596 19012 15652 19126
rect 15596 18946 15652 18956
rect 15820 19178 15876 19190
rect 15820 19126 15822 19178
rect 15874 19126 15876 19178
rect 14028 18450 14532 18452
rect 14028 18398 14030 18450
rect 14082 18398 14532 18450
rect 14028 18396 14532 18398
rect 15036 18620 15316 18676
rect 15820 18676 15876 19126
rect 15036 18452 15092 18620
rect 15820 18610 15876 18620
rect 15932 19178 15988 19190
rect 15932 19126 15934 19178
rect 15986 19126 15988 19178
rect 13580 18004 13636 18014
rect 13356 17836 13524 17892
rect 13356 17668 13412 17678
rect 13132 17666 13412 17668
rect 13132 17614 13358 17666
rect 13410 17614 13412 17666
rect 13132 17612 13412 17614
rect 13356 17602 13412 17612
rect 12796 16994 12852 17052
rect 12796 16942 12798 16994
rect 12850 16942 12852 16994
rect 12796 16930 12852 16942
rect 13356 16996 13412 17006
rect 13468 16996 13524 17836
rect 13580 17666 13636 17948
rect 13580 17614 13582 17666
rect 13634 17614 13636 17666
rect 13580 17602 13636 17614
rect 13860 17668 13916 17678
rect 13860 17574 13916 17612
rect 13356 16994 13524 16996
rect 13356 16942 13358 16994
rect 13410 16942 13524 16994
rect 13356 16940 13524 16942
rect 13356 16930 13412 16940
rect 12012 16046 12014 16098
rect 12066 16046 12068 16098
rect 12012 16034 12068 16046
rect 13468 16100 13524 16940
rect 13692 16884 13748 16894
rect 13692 16100 13748 16828
rect 14028 16884 14084 18396
rect 14812 18338 14868 18350
rect 14812 18286 14814 18338
rect 14866 18286 14868 18338
rect 14812 17780 14868 18286
rect 14812 17714 14868 17724
rect 15036 17668 15092 18396
rect 15540 18116 15596 18126
rect 15540 17722 15596 18060
rect 15932 18116 15988 19126
rect 15932 18050 15988 18060
rect 16156 17892 16212 19404
rect 16436 19348 16492 19358
rect 16436 19290 16492 19292
rect 16268 19236 16324 19246
rect 16436 19238 16438 19290
rect 16490 19238 16492 19290
rect 16436 19226 16492 19238
rect 16716 19234 16772 19628
rect 17724 19572 17780 19993
rect 16996 19516 17780 19572
rect 16996 19458 17052 19516
rect 16996 19406 16998 19458
rect 17050 19406 17052 19458
rect 16996 19394 17052 19406
rect 17836 19358 17892 20132
rect 18060 20020 18116 20030
rect 17780 19346 17892 19358
rect 17780 19294 17782 19346
rect 17834 19294 17892 19346
rect 17780 19292 17892 19294
rect 17948 20018 18116 20020
rect 17948 19966 18062 20018
rect 18114 19966 18116 20018
rect 17948 19964 18116 19966
rect 17780 19282 17836 19292
rect 16268 19142 16324 19180
rect 16716 19182 16718 19234
rect 16770 19182 16772 19234
rect 16716 19170 16772 19182
rect 16604 19124 16660 19134
rect 17948 19124 18004 19964
rect 18060 19954 18116 19964
rect 18172 19796 18228 22082
rect 18508 21252 18564 22318
rect 18620 21364 18676 24108
rect 18732 23938 18788 23950
rect 18732 23886 18734 23938
rect 18786 23886 18788 23938
rect 18732 23604 18788 23886
rect 18844 23716 18900 24444
rect 18956 23940 19012 26236
rect 19068 26226 19124 26236
rect 19180 25620 19236 26796
rect 19404 26906 19460 26918
rect 19404 26854 19406 26906
rect 19458 26854 19460 26906
rect 19404 26180 19460 26854
rect 21532 26852 21588 27022
rect 21532 26786 21588 26796
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19404 26124 19796 26180
rect 19180 25554 19236 25564
rect 19628 25620 19684 25630
rect 19628 25526 19684 25564
rect 19740 25508 19796 26124
rect 19852 26178 19908 26190
rect 19852 26126 19854 26178
rect 19906 26126 19908 26178
rect 19852 25732 19908 26126
rect 19852 25666 19908 25676
rect 20188 25956 20244 25966
rect 19964 25508 20020 25518
rect 19740 25506 20020 25508
rect 19740 25454 19966 25506
rect 20018 25454 20020 25506
rect 19740 25452 20020 25454
rect 19964 25442 20020 25452
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 18956 23874 19012 23884
rect 18844 23660 19012 23716
rect 18732 23538 18788 23548
rect 18788 23380 18844 23390
rect 18844 23324 18900 23380
rect 18788 23286 18900 23324
rect 18620 21298 18676 21308
rect 18732 22370 18788 22382
rect 18732 22318 18734 22370
rect 18786 22318 18788 22370
rect 18732 21252 18788 22318
rect 18844 21812 18900 23286
rect 18956 23154 19012 23660
rect 19292 23604 19348 23614
rect 19292 23378 19348 23548
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20188 23380 20244 25900
rect 21644 25742 21700 27804
rect 21980 27894 22036 27906
rect 21980 27842 21982 27894
rect 22034 27842 22036 27894
rect 21980 27524 22036 27842
rect 22428 27894 22484 27906
rect 22428 27860 22430 27894
rect 22482 27860 22484 27894
rect 22584 27898 22640 28364
rect 22764 27970 22820 29148
rect 22764 27918 22766 27970
rect 22818 27918 22820 27970
rect 22764 27906 22820 27918
rect 22876 29148 23044 29204
rect 23380 29204 23436 29214
rect 22584 27846 22586 27898
rect 22638 27846 22640 27898
rect 22584 27834 22640 27846
rect 22428 27636 22484 27804
rect 22428 27580 22596 27636
rect 21980 27458 22036 27468
rect 21868 27074 21924 27086
rect 21868 27022 21870 27074
rect 21922 27022 21924 27074
rect 21756 26404 21812 26414
rect 21868 26404 21924 27022
rect 21756 26402 21924 26404
rect 21756 26350 21758 26402
rect 21810 26350 21924 26402
rect 21756 26348 21924 26350
rect 21756 26338 21812 26348
rect 20300 25732 20356 25742
rect 21644 25730 21756 25742
rect 21644 25678 21702 25730
rect 21754 25678 21756 25730
rect 21644 25676 21756 25678
rect 20300 25638 20356 25676
rect 21700 25666 21756 25676
rect 21868 25506 21924 26348
rect 22316 26740 22372 26750
rect 22316 26290 22372 26684
rect 22316 26238 22318 26290
rect 22370 26238 22372 26290
rect 22316 26226 22372 26238
rect 22540 26122 22596 27580
rect 22744 27524 22800 27534
rect 22744 27074 22800 27468
rect 22744 27022 22746 27074
rect 22798 27022 22800 27074
rect 22744 26908 22800 27022
rect 22744 26852 22820 26908
rect 22540 26070 22542 26122
rect 22594 26070 22596 26122
rect 22540 26058 22596 26070
rect 22764 26404 22820 26852
rect 22764 25620 22820 26348
rect 22764 25554 22820 25564
rect 21868 25454 21870 25506
rect 21922 25454 21924 25506
rect 21868 25442 21924 25454
rect 22764 25284 22820 25294
rect 22540 25282 22820 25284
rect 22540 25230 22766 25282
rect 22818 25230 22820 25282
rect 22540 25228 22820 25230
rect 21084 24749 21140 24761
rect 19292 23326 19294 23378
rect 19346 23326 19348 23378
rect 19292 23314 19348 23326
rect 20076 23324 20244 23380
rect 20412 24724 20468 24734
rect 20412 24498 20468 24668
rect 20412 24446 20414 24498
rect 20466 24446 20468 24498
rect 20412 23940 20468 24446
rect 18956 23102 18958 23154
rect 19010 23102 19012 23154
rect 18956 23090 19012 23102
rect 19908 23156 19964 23166
rect 19908 23062 19964 23100
rect 19012 22372 19068 22382
rect 19292 22372 19348 22382
rect 19012 22370 19348 22372
rect 19012 22318 19014 22370
rect 19066 22318 19294 22370
rect 19346 22318 19348 22370
rect 19012 22316 19348 22318
rect 19012 22306 19068 22316
rect 19292 22306 19348 22316
rect 18844 21746 18900 21756
rect 19628 22146 19684 22158
rect 19628 22094 19630 22146
rect 19682 22094 19684 22146
rect 19628 21588 19684 22094
rect 20076 22148 20132 23324
rect 20076 22092 20244 22148
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19852 21588 19908 21598
rect 19628 21586 19908 21588
rect 19628 21534 19854 21586
rect 19906 21534 19908 21586
rect 19628 21532 19908 21534
rect 19852 21522 19908 21532
rect 20188 21252 20244 22092
rect 20412 21588 20468 23884
rect 21084 24697 21086 24749
rect 21138 24697 21140 24749
rect 20636 23826 20692 23838
rect 20636 23774 20638 23826
rect 20690 23774 20692 23826
rect 20636 23044 20692 23774
rect 21084 23380 21140 24697
rect 21756 24724 21812 24734
rect 21756 24630 21812 24668
rect 22540 24722 22596 25228
rect 22764 25218 22820 25228
rect 22876 24948 22932 29148
rect 23380 29110 23436 29148
rect 23324 28980 23380 28990
rect 23212 27860 23268 27870
rect 22988 27858 23268 27860
rect 22988 27806 23214 27858
rect 23266 27806 23268 27858
rect 22988 27804 23268 27806
rect 22988 27298 23044 27804
rect 23212 27794 23268 27804
rect 23324 27690 23380 28924
rect 23436 27860 23492 27870
rect 23436 27766 23492 27804
rect 23324 27638 23326 27690
rect 23378 27638 23380 27690
rect 23324 27626 23380 27638
rect 22988 27246 22990 27298
rect 23042 27246 23044 27298
rect 22988 27234 23044 27246
rect 23100 27188 23156 27198
rect 23100 26628 23156 27132
rect 23056 26572 23156 26628
rect 23056 26328 23112 26572
rect 23056 26276 23058 26328
rect 23110 26276 23112 26328
rect 23056 26264 23112 26276
rect 23436 25620 23492 25630
rect 23436 25526 23492 25564
rect 22540 24670 22542 24722
rect 22594 24670 22596 24722
rect 22540 24658 22596 24670
rect 22764 24892 22932 24948
rect 23100 25506 23156 25518
rect 23100 25454 23102 25506
rect 23154 25454 23156 25506
rect 23100 24948 23156 25454
rect 22764 24164 22820 24892
rect 23100 24882 23156 24892
rect 23884 24948 23940 24958
rect 23772 24612 23828 24622
rect 22764 24108 22932 24164
rect 22671 24052 22727 24062
rect 21756 23940 21812 23950
rect 22428 23940 22484 23950
rect 21756 23938 21924 23940
rect 21756 23886 21758 23938
rect 21810 23886 21924 23938
rect 21756 23884 21924 23886
rect 21756 23874 21812 23884
rect 21420 23716 21476 23726
rect 21420 23622 21476 23660
rect 20916 23322 20972 23334
rect 20916 23270 20918 23322
rect 20970 23270 20972 23322
rect 21084 23314 21140 23324
rect 20916 23268 20972 23270
rect 20916 23202 20972 23212
rect 20636 22978 20692 22988
rect 21084 23154 21140 23166
rect 21084 23102 21086 23154
rect 21138 23102 21140 23154
rect 21084 23044 21140 23102
rect 21084 22978 21140 22988
rect 21868 23064 21924 23884
rect 22428 23846 22484 23884
rect 22671 23938 22727 23996
rect 22671 23886 22673 23938
rect 22725 23886 22727 23938
rect 22671 23874 22727 23886
rect 21868 23042 21980 23064
rect 21868 22990 21926 23042
rect 21978 22990 21980 23042
rect 21868 22978 21980 22990
rect 20860 22372 20916 22382
rect 20860 22278 20916 22316
rect 21420 22370 21476 22382
rect 21420 22318 21422 22370
rect 21474 22318 21476 22370
rect 20524 22148 20580 22158
rect 20524 22054 20580 22092
rect 20636 21588 20692 21598
rect 20412 21586 20692 21588
rect 20412 21534 20638 21586
rect 20690 21534 20692 21586
rect 20412 21532 20692 21534
rect 20636 21522 20692 21532
rect 20972 21474 21028 21486
rect 20972 21422 20974 21474
rect 21026 21422 21028 21474
rect 18732 21196 19572 21252
rect 18508 21186 18564 21196
rect 19272 21028 19328 21038
rect 18396 20802 18452 20814
rect 18396 20750 18398 20802
rect 18450 20750 18452 20802
rect 18396 20356 18452 20750
rect 18396 20290 18452 20300
rect 18508 20804 18564 20814
rect 18508 19908 18564 20748
rect 19272 20802 19328 20972
rect 19516 21026 19572 21196
rect 20188 21186 20244 21196
rect 20356 21252 20412 21262
rect 19516 20974 19518 21026
rect 19570 20974 19572 21026
rect 19516 20962 19572 20974
rect 20188 21028 20244 21038
rect 19272 20750 19274 20802
rect 19326 20750 19328 20802
rect 19272 20738 19328 20750
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 18620 20132 18900 20188
rect 20188 20142 20244 20972
rect 20356 20914 20412 21196
rect 20356 20862 20358 20914
rect 20410 20862 20412 20914
rect 20356 20850 20412 20862
rect 20860 20804 20916 20814
rect 20972 20804 21028 21422
rect 21420 21038 21476 22318
rect 21644 22372 21700 22382
rect 21644 21252 21700 22316
rect 21756 22146 21812 22158
rect 21756 22094 21758 22146
rect 21810 22094 21812 22146
rect 21756 21588 21812 22094
rect 21868 22036 21924 22978
rect 21868 21970 21924 21980
rect 22484 22708 22540 22718
rect 22484 22146 22540 22652
rect 22484 22094 22486 22146
rect 22538 22094 22540 22146
rect 22484 21812 22540 22094
rect 22484 21746 22540 21756
rect 22652 21812 22708 21822
rect 22876 21812 22932 24108
rect 23548 23940 23604 23950
rect 23772 23940 23828 24556
rect 23884 24174 23940 24892
rect 23884 24162 23996 24174
rect 23884 24110 23942 24162
rect 23994 24110 23996 24162
rect 23884 24108 23996 24110
rect 23940 24098 23996 24108
rect 23548 23938 23828 23940
rect 23548 23886 23550 23938
rect 23602 23886 23828 23938
rect 23548 23884 23828 23886
rect 23548 23874 23604 23884
rect 24108 23044 24164 29474
rect 24444 29092 24500 29102
rect 24220 28644 24276 28654
rect 24220 27188 24276 28588
rect 24220 27094 24276 27132
rect 24276 26180 24332 26190
rect 24276 26086 24332 26124
rect 24444 25844 24500 29036
rect 24668 28868 24724 30828
rect 24780 30772 24836 30782
rect 24780 29426 24836 30716
rect 25284 30772 25340 30782
rect 25284 30678 25340 30716
rect 25452 30100 25508 30940
rect 24780 29374 24782 29426
rect 24834 29374 24836 29426
rect 24780 29362 24836 29374
rect 25116 30098 25508 30100
rect 25116 30046 25454 30098
rect 25506 30046 25508 30098
rect 25116 30044 25508 30046
rect 24948 28868 25004 28878
rect 24668 28866 25004 28868
rect 24668 28814 24950 28866
rect 25002 28814 25004 28866
rect 24668 28812 25004 28814
rect 24948 28802 25004 28812
rect 25116 28642 25172 30044
rect 25452 30034 25508 30044
rect 25340 29428 25396 29438
rect 25340 29334 25396 29372
rect 25676 29428 25732 31500
rect 25788 31220 25844 33068
rect 26684 32788 26740 37324
rect 27132 37314 27188 37326
rect 27580 37324 27748 37380
rect 26888 37266 26944 37278
rect 26888 37214 26890 37266
rect 26942 37214 26944 37266
rect 26888 37044 26944 37214
rect 26888 36978 26944 36988
rect 27020 36596 27076 36606
rect 27580 36596 27636 37324
rect 27748 37154 27804 37166
rect 27748 37102 27750 37154
rect 27802 37102 27804 37154
rect 27748 37044 27804 37102
rect 27748 36978 27804 36988
rect 28140 36596 28196 38612
rect 28364 38612 28420 39228
rect 28812 39060 28868 43372
rect 28924 43204 28980 43514
rect 28924 43138 28980 43148
rect 29036 42754 29092 44044
rect 29148 43988 29204 45836
rect 29428 45808 29430 45836
rect 29482 45808 29484 45860
rect 29428 45796 29484 45808
rect 30044 45798 30100 45836
rect 30268 45892 30324 46622
rect 30380 46676 30436 46686
rect 30492 46676 30548 47404
rect 30828 47458 30884 47470
rect 30828 47406 30830 47458
rect 30882 47406 30884 47458
rect 30828 47012 30884 47406
rect 30716 46956 30884 47012
rect 31164 47234 31220 47246
rect 31164 47182 31166 47234
rect 31218 47182 31220 47234
rect 31164 47012 31220 47182
rect 30604 46676 30660 46686
rect 30492 46674 30660 46676
rect 30492 46622 30606 46674
rect 30658 46622 30660 46674
rect 30492 46620 30660 46622
rect 30380 46582 30436 46620
rect 30604 46610 30660 46620
rect 30268 45826 30324 45836
rect 30716 45274 30772 46956
rect 31164 46946 31220 46956
rect 31444 46705 31500 46715
rect 31444 46703 31556 46705
rect 31444 46651 31446 46703
rect 31498 46651 31556 46703
rect 31444 46639 31556 46651
rect 31276 46564 31332 46574
rect 31052 46562 31332 46564
rect 31052 46510 31278 46562
rect 31330 46510 31332 46562
rect 31052 46508 31332 46510
rect 30884 46452 30940 46462
rect 30884 46358 30940 46396
rect 30828 46004 30884 46014
rect 30828 45910 30884 45948
rect 31052 45444 31108 46508
rect 31276 46498 31332 46508
rect 31500 46452 31556 46639
rect 31500 46228 31556 46396
rect 31724 46674 31780 46686
rect 31724 46622 31726 46674
rect 31778 46622 31780 46674
rect 31724 46340 31780 46622
rect 31836 46676 31892 47966
rect 39284 48132 39340 48142
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 38836 47684 38892 47694
rect 32620 47572 32676 47582
rect 32620 47478 32676 47516
rect 33852 47572 33908 47582
rect 32172 47458 32228 47470
rect 32172 47406 32174 47458
rect 32226 47406 32228 47458
rect 32172 47236 32228 47406
rect 32172 47170 32228 47180
rect 32508 47414 32564 47426
rect 32508 47362 32510 47414
rect 32562 47362 32564 47414
rect 32508 47124 32564 47362
rect 32508 47058 32564 47068
rect 33740 47234 33796 47246
rect 33740 47182 33742 47234
rect 33794 47182 33796 47234
rect 32060 46676 32116 46686
rect 31836 46674 32116 46676
rect 31836 46622 32062 46674
rect 32114 46622 32116 46674
rect 31836 46620 32116 46622
rect 32060 46610 32116 46620
rect 32956 46676 33012 46686
rect 32956 46582 33012 46620
rect 33628 46562 33684 46574
rect 33628 46510 33630 46562
rect 33682 46510 33684 46562
rect 32396 46450 32452 46462
rect 33124 46452 33180 46462
rect 32396 46398 32398 46450
rect 32450 46398 32452 46450
rect 31724 46284 32116 46340
rect 31500 46172 32004 46228
rect 31724 45668 31780 45678
rect 31052 45388 31332 45444
rect 30716 45222 30718 45274
rect 30770 45222 30772 45274
rect 30716 45210 30772 45222
rect 31052 45145 31108 45157
rect 30604 45108 30660 45118
rect 30604 45014 30660 45052
rect 31052 45108 31054 45145
rect 31106 45108 31108 45145
rect 31052 45042 31108 45052
rect 31276 45106 31332 45388
rect 31276 45054 31278 45106
rect 31330 45054 31332 45106
rect 31276 45042 31332 45054
rect 31724 45106 31780 45612
rect 31724 45054 31726 45106
rect 31778 45054 31780 45106
rect 29540 44994 29596 45006
rect 29540 44942 29542 44994
rect 29594 44942 29596 44994
rect 29260 44772 29316 44782
rect 29260 44322 29316 44716
rect 29260 44270 29262 44322
rect 29314 44270 29316 44322
rect 29260 44258 29316 44270
rect 29372 44660 29428 44670
rect 29372 44548 29428 44604
rect 29540 44548 29596 44942
rect 31724 44884 31780 45054
rect 31948 45106 32004 46172
rect 32060 45668 32116 46284
rect 32060 45602 32116 45612
rect 31948 45054 31950 45106
rect 32002 45054 32004 45106
rect 31948 45042 32004 45054
rect 32228 45108 32284 45118
rect 29372 44492 29596 44548
rect 31276 44828 31780 44884
rect 29372 44100 29428 44492
rect 30604 44490 30660 44502
rect 30604 44438 30606 44490
rect 30658 44438 30660 44490
rect 29540 44324 29596 44334
rect 29540 44230 29596 44268
rect 30156 44322 30212 44334
rect 30156 44270 30158 44322
rect 30210 44270 30212 44322
rect 29148 43922 29204 43932
rect 29260 44044 29428 44100
rect 29148 43566 29204 43578
rect 29148 43514 29150 43566
rect 29202 43514 29204 43566
rect 29148 43428 29204 43514
rect 29148 43362 29204 43372
rect 29260 43573 29316 44044
rect 29260 43521 29262 43573
rect 29314 43521 29316 43573
rect 29260 42980 29316 43521
rect 29036 42702 29038 42754
rect 29090 42702 29092 42754
rect 29036 42690 29092 42702
rect 29148 42924 29316 42980
rect 29372 43540 29428 43550
rect 29148 42308 29204 42924
rect 29260 42756 29316 42766
rect 29260 42662 29316 42700
rect 29148 42242 29204 42252
rect 28980 41860 29036 41870
rect 28980 41412 29036 41804
rect 28980 41356 29204 41412
rect 29036 41188 29092 41198
rect 29036 41094 29092 41132
rect 28980 40628 29036 40638
rect 28980 40514 29036 40572
rect 28980 40462 28982 40514
rect 29034 40462 29036 40514
rect 28980 40450 29036 40462
rect 28812 38994 28868 39004
rect 28812 38834 28868 38846
rect 28812 38782 28814 38834
rect 28866 38782 28868 38834
rect 28364 37502 28420 38556
rect 28476 38722 28532 38734
rect 28476 38670 28478 38722
rect 28530 38670 28532 38722
rect 28476 38388 28532 38670
rect 28812 38668 28868 38782
rect 28924 38836 28980 38846
rect 28924 38834 29092 38836
rect 28924 38782 28926 38834
rect 28978 38782 29092 38834
rect 28924 38780 29092 38782
rect 28924 38770 28980 38780
rect 28476 38322 28532 38332
rect 28588 38612 28868 38668
rect 28476 38164 28532 38174
rect 28588 38164 28644 38612
rect 28476 38162 28588 38164
rect 28476 38110 28478 38162
rect 28530 38110 28588 38162
rect 28476 38108 28588 38110
rect 28476 38098 28532 38108
rect 28588 38070 28644 38108
rect 28924 38276 28980 38286
rect 28308 37492 28420 37502
rect 28308 37490 28644 37492
rect 28308 37438 28310 37490
rect 28362 37438 28644 37490
rect 28308 37436 28644 37438
rect 28308 37426 28364 37436
rect 28588 37266 28644 37436
rect 28588 37214 28590 37266
rect 28642 37214 28644 37266
rect 28588 37202 28644 37214
rect 28924 37281 28980 38220
rect 28924 37229 28926 37281
rect 28978 37229 28980 37281
rect 27020 36594 27748 36596
rect 27020 36542 27022 36594
rect 27074 36542 27748 36594
rect 27020 36540 27748 36542
rect 28140 36540 28532 36596
rect 27020 36530 27076 36540
rect 27692 36484 27748 36540
rect 28028 36484 28084 36494
rect 27692 36447 27804 36484
rect 27692 36428 27750 36447
rect 27748 36395 27750 36428
rect 27802 36395 27804 36447
rect 27748 36383 27804 36395
rect 28028 36402 28030 36428
rect 28082 36402 28084 36428
rect 28028 36390 28084 36402
rect 28252 36426 28308 36438
rect 27356 36372 27412 36382
rect 27356 35754 27412 36316
rect 27524 36370 27580 36382
rect 27524 36318 27526 36370
rect 27578 36318 27580 36370
rect 27524 36036 27580 36318
rect 28252 36374 28254 36426
rect 28306 36374 28308 36426
rect 27524 35970 27580 35980
rect 28028 36260 28084 36270
rect 27132 35726 27188 35738
rect 27132 35700 27134 35726
rect 27186 35700 27188 35726
rect 27356 35702 27358 35754
rect 27410 35702 27412 35754
rect 27692 35812 27748 35822
rect 27692 35754 27748 35756
rect 27356 35690 27412 35702
rect 27580 35726 27636 35738
rect 27132 35634 27188 35644
rect 27580 35674 27582 35726
rect 27634 35674 27636 35726
rect 27692 35702 27694 35754
rect 27746 35702 27748 35754
rect 27692 35690 27748 35702
rect 26852 35474 26908 35486
rect 26852 35422 26854 35474
rect 26906 35422 26908 35474
rect 26852 35252 26908 35422
rect 27580 35476 27636 35674
rect 27580 35410 27636 35420
rect 26796 35196 26908 35252
rect 26796 34692 26852 35196
rect 27020 34692 27076 34702
rect 26796 34636 26964 34692
rect 26908 34130 26964 34636
rect 26908 34078 26910 34130
rect 26962 34078 26964 34130
rect 26908 34066 26964 34078
rect 26852 33236 26908 33246
rect 26852 33142 26908 33180
rect 27020 32788 27076 34636
rect 27244 34356 27300 34366
rect 27244 34262 27300 34300
rect 26348 32732 26740 32788
rect 26796 32732 27076 32788
rect 27692 34244 27748 34254
rect 26012 32450 26068 32462
rect 26012 32398 26014 32450
rect 26066 32398 26068 32450
rect 26012 32004 26068 32398
rect 26012 31938 26068 31948
rect 25956 31780 26012 31790
rect 26236 31780 26292 31790
rect 25956 31778 26292 31780
rect 25956 31726 25958 31778
rect 26010 31726 26238 31778
rect 26290 31726 26292 31778
rect 25956 31724 26292 31726
rect 25956 31714 26012 31724
rect 26236 31714 26292 31724
rect 25788 31154 25844 31164
rect 26124 31332 26180 31342
rect 26124 31050 26180 31276
rect 25788 31022 25844 31034
rect 25788 30996 25790 31022
rect 25842 30996 25844 31022
rect 25956 31029 26012 31041
rect 25956 30996 25958 31029
rect 25788 30930 25844 30940
rect 25900 30977 25958 30996
rect 26010 30977 26012 31029
rect 26124 30998 26126 31050
rect 26178 30998 26180 31050
rect 26124 30986 26180 30998
rect 25900 30940 26012 30977
rect 25676 29362 25732 29372
rect 25676 29204 25732 29214
rect 25900 29204 25956 30940
rect 26012 30212 26068 30222
rect 26012 30118 26068 30156
rect 26124 29652 26180 29662
rect 26124 29482 26180 29596
rect 26124 29430 26126 29482
rect 26178 29430 26180 29482
rect 26124 29418 26180 29430
rect 26236 29454 26292 29466
rect 26236 29402 26238 29454
rect 26290 29402 26292 29454
rect 26236 29204 26292 29402
rect 25676 29202 26292 29204
rect 25676 29150 25678 29202
rect 25730 29150 26292 29202
rect 25676 29148 26292 29150
rect 25676 29138 25732 29148
rect 25732 28756 25788 28766
rect 25732 28662 25788 28700
rect 25116 28590 25118 28642
rect 25170 28590 25172 28642
rect 25116 28578 25172 28590
rect 25676 27885 25732 27897
rect 25676 27833 25678 27885
rect 25730 27833 25732 27885
rect 25396 27748 25452 27758
rect 25396 27654 25452 27692
rect 25676 27748 25732 27833
rect 25676 27682 25732 27692
rect 25452 26852 25508 26862
rect 25340 26628 25396 26638
rect 25340 26346 25396 26572
rect 25228 26325 25284 26337
rect 24724 26292 24780 26302
rect 24724 26198 24780 26236
rect 25228 26292 25230 26325
rect 25282 26292 25284 26325
rect 25340 26294 25342 26346
rect 25394 26294 25396 26346
rect 25340 26282 25396 26294
rect 24220 25788 24500 25844
rect 24220 24836 24276 25788
rect 24220 24770 24276 24780
rect 25116 24722 25172 24734
rect 25116 24670 25118 24722
rect 25170 24670 25172 24722
rect 24444 24612 24500 24622
rect 24444 24518 24500 24556
rect 24220 23940 24276 23950
rect 24220 23846 24276 23884
rect 24444 23940 24500 23950
rect 24500 23884 24612 23940
rect 24444 23846 24500 23884
rect 23548 22988 24164 23044
rect 23212 22370 23268 22382
rect 23212 22318 23214 22370
rect 23266 22318 23268 22370
rect 23212 21924 23268 22318
rect 23212 21858 23268 21868
rect 21756 21522 21812 21532
rect 22428 21252 22484 21262
rect 21644 21196 21924 21252
rect 21364 21026 21476 21038
rect 21364 20974 21366 21026
rect 21418 20974 21476 21026
rect 21364 20972 21476 20974
rect 21364 20962 21420 20972
rect 20860 20802 21644 20804
rect 20860 20750 20862 20802
rect 20914 20767 21644 20802
rect 20914 20750 21590 20767
rect 20860 20748 21590 20750
rect 20860 20738 20916 20748
rect 21588 20715 21590 20748
rect 21642 20715 21644 20767
rect 21588 20703 21644 20715
rect 21868 20774 21924 21196
rect 21868 20722 21870 20774
rect 21922 20722 21924 20774
rect 21868 20710 21924 20722
rect 22092 21140 22148 21150
rect 22092 20774 22148 21084
rect 22092 20722 22094 20774
rect 22146 20722 22148 20774
rect 22428 20802 22484 21196
rect 22652 21252 22708 21756
rect 22652 21186 22708 21196
rect 22764 21756 22932 21812
rect 22764 21028 22820 21756
rect 22876 21588 22932 21598
rect 22876 21494 22932 21532
rect 22092 20710 22148 20722
rect 22204 20746 22260 20758
rect 22204 20694 22206 20746
rect 22258 20694 22260 20746
rect 22204 20692 22260 20694
rect 22204 20626 22260 20636
rect 22428 20750 22430 20802
rect 22482 20750 22484 20802
rect 20692 20580 20748 20590
rect 20524 20578 20748 20580
rect 20524 20526 20694 20578
rect 20746 20526 20748 20578
rect 20524 20524 20748 20526
rect 18620 19908 18676 20132
rect 18508 19852 18676 19908
rect 16604 19030 16660 19068
rect 17780 19068 18004 19124
rect 18060 19740 18228 19796
rect 18620 19850 18676 19852
rect 18620 19798 18622 19850
rect 18674 19798 18676 19850
rect 18620 19786 18676 19798
rect 18732 20018 18788 20030
rect 18732 19966 18734 20018
rect 18786 19966 18788 20018
rect 18732 19908 18788 19966
rect 16156 17826 16212 17836
rect 16492 18900 16548 18910
rect 15148 17668 15204 17678
rect 15036 17666 15204 17668
rect 14812 17610 14868 17622
rect 15036 17614 15150 17666
rect 15202 17614 15204 17666
rect 15540 17670 15542 17722
rect 15594 17670 15596 17722
rect 15820 17780 15876 17790
rect 15820 17686 15876 17724
rect 15540 17658 15596 17670
rect 16156 17666 16212 17678
rect 15036 17612 15204 17614
rect 14812 17558 14814 17610
rect 14866 17558 14868 17610
rect 15148 17602 15204 17612
rect 15932 17622 15988 17634
rect 15932 17570 15934 17622
rect 15986 17570 15988 17622
rect 14812 17556 14868 17558
rect 14868 17500 15092 17556
rect 14812 17490 14868 17500
rect 15036 17220 15092 17500
rect 15372 17554 15428 17566
rect 15372 17502 15374 17554
rect 15426 17502 15428 17554
rect 15372 17444 15428 17502
rect 15932 17444 15988 17570
rect 15372 17388 15988 17444
rect 16156 17614 16158 17666
rect 16210 17614 16212 17666
rect 16156 17444 16212 17614
rect 16492 17666 16548 18844
rect 17500 18564 17556 18574
rect 17276 18450 17332 18462
rect 17276 18398 17278 18450
rect 17330 18398 17332 18450
rect 16716 18338 16772 18350
rect 16716 18286 16718 18338
rect 16770 18286 16772 18338
rect 16716 18116 16772 18286
rect 16716 18050 16772 18060
rect 17276 18116 17332 18398
rect 17500 18450 17556 18508
rect 17780 18562 17836 19068
rect 17780 18510 17782 18562
rect 17834 18510 17836 18562
rect 17780 18498 17836 18510
rect 17500 18398 17502 18450
rect 17554 18398 17556 18450
rect 17500 18386 17556 18398
rect 17276 18050 17332 18060
rect 18060 17892 18116 19740
rect 18732 19460 18788 19852
rect 18620 19404 18788 19460
rect 18172 19122 18228 19134
rect 18172 19070 18174 19122
rect 18226 19070 18228 19122
rect 18172 18900 18228 19070
rect 18172 18844 18452 18900
rect 18396 18485 18452 18844
rect 18620 18564 18676 19404
rect 18844 18564 18900 20132
rect 19852 20132 19908 20142
rect 20188 20130 20300 20142
rect 20188 20078 20246 20130
rect 20298 20078 20300 20130
rect 20188 20076 20300 20078
rect 18956 20018 19012 20030
rect 19292 20020 19348 20030
rect 18956 19966 18958 20018
rect 19010 19966 19012 20018
rect 18956 19908 19012 19966
rect 18956 19842 19012 19852
rect 19068 20018 19348 20020
rect 19068 19966 19294 20018
rect 19346 19966 19348 20018
rect 19068 19964 19348 19966
rect 19068 19572 19124 19964
rect 19292 19954 19348 19964
rect 19628 19796 19684 19806
rect 19628 19702 19684 19740
rect 18956 19516 19124 19572
rect 18956 19012 19012 19516
rect 19852 19012 19908 20076
rect 20244 20066 20300 20076
rect 20412 20020 20468 20030
rect 20188 19908 20244 19918
rect 20076 19796 20132 19806
rect 20076 19346 20132 19740
rect 20076 19294 20078 19346
rect 20130 19294 20132 19346
rect 20076 19282 20132 19294
rect 18956 18956 19292 19012
rect 18396 18433 18398 18485
rect 18450 18433 18452 18485
rect 18564 18508 18676 18564
rect 18564 18506 18620 18508
rect 18564 18454 18566 18506
rect 18618 18454 18620 18506
rect 18564 18442 18620 18454
rect 18788 18506 18900 18564
rect 18788 18454 18790 18506
rect 18842 18454 18900 18506
rect 19236 18562 19292 18956
rect 19236 18510 19238 18562
rect 19290 18510 19292 18562
rect 19236 18498 19292 18510
rect 19628 18956 19908 19012
rect 18788 18442 18900 18454
rect 18396 18340 18452 18433
rect 18396 18274 18452 18284
rect 18060 17826 18116 17836
rect 18396 17892 18452 17902
rect 16492 17614 16494 17666
rect 16546 17614 16548 17666
rect 16492 17602 16548 17614
rect 16716 17668 16772 17678
rect 16716 17574 16772 17612
rect 17948 17668 18004 17678
rect 17948 17574 18004 17612
rect 18396 17666 18452 17836
rect 18396 17614 18398 17666
rect 18450 17614 18452 17666
rect 18396 17602 18452 17614
rect 18844 17668 18900 18442
rect 18956 18478 19012 18490
rect 18956 18452 18958 18478
rect 19010 18452 19012 18478
rect 18956 18386 19012 18396
rect 19348 17892 19404 17902
rect 19348 17778 19404 17836
rect 19348 17726 19350 17778
rect 19402 17726 19404 17778
rect 19348 17714 19404 17726
rect 18844 17602 18900 17612
rect 16996 17556 17052 17566
rect 16996 17462 17052 17500
rect 16156 17378 16212 17388
rect 16604 17444 16660 17454
rect 15036 17164 15204 17220
rect 14028 16818 14084 16828
rect 15036 16996 15092 17006
rect 15036 16322 15092 16940
rect 15036 16270 15038 16322
rect 15090 16270 15092 16322
rect 15036 16258 15092 16270
rect 13916 16100 13972 16110
rect 13692 16044 13860 16100
rect 13468 16034 13524 16044
rect 13636 15876 13692 15886
rect 13636 15782 13692 15820
rect 12236 15316 12292 15326
rect 9996 14532 10052 15036
rect 11116 15036 11228 15092
rect 10444 14644 10500 14654
rect 10444 14550 10500 14588
rect 9996 14466 10052 14476
rect 10220 14532 10276 14542
rect 8988 12014 8990 12066
rect 9042 12014 9044 12066
rect 8988 12002 9044 12014
rect 9212 12796 9380 12852
rect 9436 13356 9828 13412
rect 9884 13773 9940 13785
rect 9884 13721 9886 13773
rect 9938 13721 9940 13773
rect 9212 11284 9268 12796
rect 9436 12740 9492 13356
rect 9884 13300 9940 13721
rect 10220 13746 10276 14476
rect 10220 13694 10222 13746
rect 10274 13694 10276 13746
rect 10220 13524 10276 13694
rect 11116 13746 11172 15036
rect 11228 15026 11284 15036
rect 11900 15314 12292 15316
rect 11900 15262 12238 15314
rect 12290 15262 12292 15314
rect 11900 15260 12292 15262
rect 11900 15092 11956 15260
rect 12236 15250 12292 15260
rect 13804 15314 13860 16044
rect 13916 16006 13972 16044
rect 14792 16100 14848 16110
rect 15148 16100 15204 17164
rect 16380 16996 16436 17006
rect 16380 16926 16436 16940
rect 16044 16884 16100 16894
rect 16380 16874 16382 16926
rect 16434 16874 16436 16926
rect 16380 16862 16436 16874
rect 16604 16882 16660 17388
rect 17612 17444 17668 17454
rect 17612 17350 17668 17388
rect 18732 17444 18788 17454
rect 18732 17442 19158 17444
rect 18732 17390 18734 17442
rect 18786 17390 19158 17442
rect 18732 17388 19158 17390
rect 18732 17378 18788 17388
rect 16044 16790 16100 16828
rect 16604 16830 16606 16882
rect 16658 16830 16660 16882
rect 16604 16818 16660 16830
rect 17836 16920 17892 16932
rect 17836 16868 17838 16920
rect 17890 16868 17892 16920
rect 19102 16920 19158 17388
rect 15260 16770 15316 16782
rect 15260 16718 15262 16770
rect 15314 16718 15316 16770
rect 15260 16660 15316 16718
rect 16268 16770 16324 16782
rect 16268 16718 16270 16770
rect 16322 16718 16324 16770
rect 16268 16660 16324 16718
rect 15260 16604 16324 16660
rect 16660 16660 16716 16670
rect 16660 16322 16716 16604
rect 16660 16270 16662 16322
rect 16714 16270 16716 16322
rect 16660 16258 16716 16270
rect 14792 16098 15204 16100
rect 14792 16046 14794 16098
rect 14846 16046 15204 16098
rect 14792 16044 15204 16046
rect 16492 16098 16548 16110
rect 16492 16046 16494 16098
rect 16546 16046 16548 16098
rect 14792 16034 14848 16044
rect 13804 15262 13806 15314
rect 13858 15262 13860 15314
rect 13804 15250 13860 15262
rect 15932 15876 15988 15886
rect 14588 15204 14644 15242
rect 14588 15138 14644 15148
rect 11900 15026 11956 15036
rect 13468 15092 13524 15102
rect 12124 14644 12180 14654
rect 11788 14532 11844 14542
rect 11788 14530 12068 14532
rect 11788 14478 11790 14530
rect 11842 14478 12068 14530
rect 11788 14476 12068 14478
rect 11788 14466 11844 14476
rect 11452 14308 11508 14318
rect 11452 14306 11956 14308
rect 11452 14254 11454 14306
rect 11506 14254 11956 14306
rect 11452 14252 11956 14254
rect 11452 14242 11508 14252
rect 11116 13694 11118 13746
rect 11170 13694 11172 13746
rect 11116 13682 11172 13694
rect 11900 13746 11956 14252
rect 11900 13694 11902 13746
rect 11954 13694 11956 13746
rect 11900 13682 11956 13694
rect 10220 13458 10276 13468
rect 9884 13234 9940 13244
rect 11900 12962 11956 12974
rect 11900 12910 11902 12962
rect 11954 12910 11956 12962
rect 11116 12850 11172 12862
rect 11116 12798 11118 12850
rect 11170 12798 11172 12850
rect 9436 12684 9772 12740
rect 9716 12402 9772 12684
rect 9716 12350 9718 12402
rect 9770 12350 9772 12402
rect 9716 11956 9772 12350
rect 10220 12346 10276 12358
rect 10220 12294 10222 12346
rect 10274 12294 10276 12346
rect 10220 12292 10276 12294
rect 10220 12226 10276 12236
rect 10444 12180 10500 12190
rect 10444 12086 10500 12124
rect 11004 12180 11060 12190
rect 11116 12180 11172 12798
rect 11900 12404 11956 12910
rect 12012 12794 12068 14476
rect 12124 14515 12180 14588
rect 13132 14644 13188 14654
rect 12124 14463 12126 14515
rect 12178 14463 12180 14515
rect 12124 14451 12180 14463
rect 12460 14532 12516 14542
rect 12460 14438 12516 14476
rect 13020 14532 13076 14542
rect 12124 14362 12180 14374
rect 12124 14310 12126 14362
rect 12178 14310 12180 14362
rect 12124 12935 12180 14310
rect 13020 13076 13076 14476
rect 12796 13020 13076 13076
rect 12124 12883 12126 12935
rect 12178 12883 12180 12935
rect 12124 12871 12180 12883
rect 12460 12962 12516 12974
rect 12460 12910 12462 12962
rect 12514 12910 12516 12962
rect 12012 12742 12014 12794
rect 12066 12742 12068 12794
rect 12012 12730 12068 12742
rect 12460 12404 12516 12910
rect 11900 12348 12068 12404
rect 11900 12205 11956 12217
rect 11004 12178 11172 12180
rect 11004 12126 11006 12178
rect 11058 12126 11172 12178
rect 11004 12124 11172 12126
rect 11564 12178 11620 12190
rect 11564 12126 11566 12178
rect 11618 12126 11620 12178
rect 11004 12068 11060 12124
rect 11004 12002 11060 12012
rect 9716 11890 9772 11900
rect 9548 11844 9604 11854
rect 9212 11218 9268 11228
rect 9324 11394 9380 11406
rect 9324 11342 9326 11394
rect 9378 11342 9380 11394
rect 8876 11172 8932 11182
rect 8876 10834 8932 11116
rect 8876 10782 8878 10834
rect 8930 10782 8932 10834
rect 8876 10770 8932 10782
rect 9324 10836 9380 11342
rect 9548 11172 9604 11788
rect 10444 11284 10500 11294
rect 9548 11116 9828 11172
rect 9324 10770 9380 10780
rect 9660 10778 9716 10790
rect 9660 10726 9662 10778
rect 9714 10726 9716 10778
rect 9660 10612 9716 10726
rect 9660 10546 9716 10556
rect 9772 10610 9828 11116
rect 9772 10558 9774 10610
rect 9826 10558 9828 10610
rect 9772 10546 9828 10558
rect 10108 10637 10164 10649
rect 10108 10585 10110 10637
rect 10162 10585 10164 10637
rect 10108 9940 10164 10585
rect 10444 10610 10500 11228
rect 11228 11282 11284 11294
rect 11228 11230 11230 11282
rect 11282 11230 11284 11282
rect 11228 11172 11284 11230
rect 11228 11106 11284 11116
rect 11564 11172 11620 12126
rect 11676 12180 11732 12190
rect 11676 12066 11732 12124
rect 11676 12014 11678 12066
rect 11730 12014 11732 12066
rect 11676 12002 11732 12014
rect 11900 12153 11902 12205
rect 11954 12153 11956 12205
rect 11900 11620 11956 12153
rect 11564 11106 11620 11116
rect 11788 11564 11900 11620
rect 11228 10724 11284 10734
rect 11228 10630 11284 10668
rect 11788 10724 11844 11564
rect 11900 11554 11956 11564
rect 11900 11396 11956 11434
rect 12012 11396 12068 12348
rect 12460 12338 12516 12348
rect 12236 12180 12292 12190
rect 12796 12180 12852 13020
rect 13132 12964 13188 14588
rect 13468 14530 13524 15036
rect 13468 14478 13470 14530
rect 13522 14478 13524 14530
rect 13468 14466 13524 14478
rect 13804 14532 13860 14542
rect 13804 13858 13860 14476
rect 13804 13806 13806 13858
rect 13858 13806 13860 13858
rect 13804 13794 13860 13806
rect 14252 14530 14308 14542
rect 14252 14478 14254 14530
rect 14306 14478 14308 14530
rect 14252 13076 14308 14478
rect 14252 13010 14308 13020
rect 13020 12908 13188 12964
rect 13692 12964 13748 12974
rect 13692 12962 14084 12964
rect 13692 12910 13694 12962
rect 13746 12910 14084 12962
rect 13692 12908 14084 12910
rect 12236 12178 12852 12180
rect 12236 12126 12238 12178
rect 12290 12126 12798 12178
rect 12850 12126 12852 12178
rect 12236 12124 12852 12126
rect 12236 12114 12292 12124
rect 12796 12114 12852 12124
rect 12908 12180 12964 12190
rect 13020 12180 13076 12908
rect 12908 12178 13076 12180
rect 12908 12126 12910 12178
rect 12962 12126 13076 12178
rect 12908 12124 13076 12126
rect 13188 12404 13244 12414
rect 13188 12290 13244 12348
rect 13188 12238 13190 12290
rect 13242 12238 13244 12290
rect 12908 12114 12964 12124
rect 11956 11340 12068 11396
rect 12348 11508 12404 11518
rect 12348 11355 12404 11452
rect 11900 11330 11956 11340
rect 12348 11303 12350 11355
rect 12402 11303 12404 11355
rect 12348 11291 12404 11303
rect 12572 11394 12628 11406
rect 12572 11342 12574 11394
rect 12626 11342 12628 11394
rect 12572 11284 12628 11342
rect 13188 11396 13244 12238
rect 13188 11330 13244 11340
rect 12012 11226 12068 11238
rect 11788 10658 11844 10668
rect 11900 11172 11956 11182
rect 10444 10558 10446 10610
rect 10498 10558 10500 10610
rect 10444 10546 10500 10558
rect 10108 9874 10164 9884
rect 10780 9828 10836 9838
rect 10780 9156 10836 9772
rect 11340 9826 11396 9838
rect 11340 9774 11342 9826
rect 11394 9774 11396 9826
rect 10892 9156 10948 9166
rect 10780 9154 10948 9156
rect 10780 9102 10894 9154
rect 10946 9102 10948 9154
rect 10780 9100 10948 9102
rect 10892 9090 10948 9100
rect 9996 9042 10052 9054
rect 9996 8990 9998 9042
rect 10050 8990 10052 9042
rect 8708 8764 8820 8820
rect 9660 8818 9716 8830
rect 9660 8766 9662 8818
rect 9714 8766 9716 8818
rect 8652 8726 8708 8764
rect 9660 8428 9716 8766
rect 9548 8372 9716 8428
rect 9996 8428 10052 8990
rect 10444 8820 10500 8830
rect 9996 8372 10164 8428
rect 8652 7588 8708 7598
rect 8652 7494 8708 7532
rect 8820 7418 8876 7430
rect 8820 7366 8822 7418
rect 8874 7366 8876 7418
rect 8820 6804 8876 7366
rect 8764 6748 8876 6804
rect 7980 6290 8036 6300
rect 8092 6412 8372 6468
rect 8428 6692 8484 6702
rect 8484 6657 8708 6692
rect 8484 6636 8654 6657
rect 7756 5964 7924 6020
rect 7140 5798 7142 5850
rect 7194 5798 7196 5850
rect 7140 5796 7196 5798
rect 7140 5730 7196 5740
rect 7308 5906 7364 5918
rect 7308 5854 7310 5906
rect 7362 5854 7364 5906
rect 7308 5796 7364 5854
rect 7420 5906 7476 5964
rect 7420 5854 7422 5906
rect 7474 5854 7476 5906
rect 7420 5842 7476 5854
rect 7308 5730 7364 5740
rect 7532 5796 7588 5806
rect 6860 5294 6862 5346
rect 6914 5294 6916 5346
rect 6860 5282 6916 5294
rect 6524 5124 6580 5134
rect 6412 5122 6580 5124
rect 6412 5070 6526 5122
rect 6578 5070 6580 5122
rect 6412 5068 6580 5070
rect 6524 5058 6580 5068
rect 7532 5122 7588 5740
rect 7700 5684 7756 5694
rect 7700 5590 7756 5628
rect 7868 5348 7924 5964
rect 8092 5908 8148 6412
rect 8428 6356 8484 6636
rect 8652 6605 8654 6636
rect 8706 6605 8708 6657
rect 8652 6593 8708 6605
rect 8260 6300 8428 6356
rect 8260 5962 8316 6300
rect 8428 6290 8484 6300
rect 8540 6132 8596 6142
rect 8260 5910 8262 5962
rect 8314 5910 8316 5962
rect 8428 6020 8484 6030
rect 8428 5926 8484 5964
rect 8260 5898 8316 5910
rect 8540 5906 8596 6076
rect 8764 6030 8820 6748
rect 8988 6634 9044 6646
rect 8988 6582 8990 6634
rect 9042 6582 9044 6634
rect 8764 6018 8876 6030
rect 8764 5966 8822 6018
rect 8874 5966 8876 6018
rect 8764 5964 8876 5966
rect 8820 5954 8876 5964
rect 8988 6020 9044 6582
rect 9436 6634 9492 6646
rect 9436 6582 9438 6634
rect 9490 6582 9492 6634
rect 9436 6132 9492 6582
rect 9548 6356 9604 8372
rect 10108 8148 10164 8372
rect 10108 8054 10164 8092
rect 9884 7700 9940 7710
rect 9660 7476 9716 7486
rect 9660 7382 9716 7420
rect 9772 6804 9828 6842
rect 9772 6738 9828 6748
rect 9548 6290 9604 6300
rect 9746 6650 9802 6662
rect 9746 6598 9748 6650
rect 9800 6598 9802 6650
rect 9746 6132 9802 6598
rect 9746 6076 9828 6132
rect 9436 6066 9492 6076
rect 8988 5954 9044 5964
rect 8092 5814 8148 5852
rect 8540 5854 8542 5906
rect 8594 5854 8596 5906
rect 7868 5282 7924 5292
rect 8428 5684 8484 5694
rect 7980 5236 8036 5246
rect 7532 5070 7534 5122
rect 7586 5070 7588 5122
rect 7532 5058 7588 5070
rect 7868 5124 7924 5147
rect 7980 5142 8036 5180
rect 8316 5234 8372 5246
rect 8316 5182 8318 5234
rect 8370 5182 8372 5234
rect 7868 5055 7870 5068
rect 7922 5055 7924 5068
rect 7868 5043 7924 5055
rect 6188 4340 6244 4350
rect 6076 4338 6244 4340
rect 6076 4286 6190 4338
rect 6242 4286 6244 4338
rect 6076 4284 6244 4286
rect 6188 4274 6244 4284
rect 6972 4340 7028 4350
rect 6972 4246 7028 4284
rect 8316 4340 8372 5182
rect 8428 5107 8484 5628
rect 8428 5055 8430 5107
rect 8482 5055 8484 5107
rect 8540 5124 8596 5854
rect 9436 5908 9492 5918
rect 8876 5348 8932 5358
rect 8540 5058 8596 5068
rect 8652 5236 8708 5246
rect 8652 5122 8708 5180
rect 8652 5070 8654 5122
rect 8706 5070 8708 5122
rect 8652 5058 8708 5070
rect 8428 5043 8484 5055
rect 8876 4450 8932 5292
rect 9212 5348 9268 5358
rect 9212 5122 9268 5292
rect 9212 5070 9214 5122
rect 9266 5070 9268 5122
rect 9212 5058 9268 5070
rect 9436 5122 9492 5852
rect 9772 5908 9828 6076
rect 9772 5842 9828 5852
rect 9884 5684 9940 7644
rect 10444 7588 10500 8764
rect 9996 7489 10052 7501
rect 9996 7437 9998 7489
rect 10050 7437 10052 7489
rect 9996 6580 10052 7437
rect 10444 7474 10500 7532
rect 10444 7422 10446 7474
rect 10498 7422 10500 7474
rect 10444 7410 10500 7422
rect 10556 8258 10612 8270
rect 10556 8206 10558 8258
rect 10610 8206 10612 8258
rect 10108 7364 10164 7374
rect 10108 7270 10164 7308
rect 10556 6916 10612 8206
rect 10668 8260 10724 8270
rect 11228 8258 11284 8270
rect 10668 8090 10724 8204
rect 10668 8038 10670 8090
rect 10722 8038 10724 8090
rect 10892 8202 10948 8214
rect 10892 8150 10894 8202
rect 10946 8150 10948 8202
rect 10892 8148 10948 8150
rect 10892 8082 10948 8092
rect 11228 8206 11230 8258
rect 11282 8206 11284 8258
rect 10668 8026 10724 8038
rect 11228 7700 11284 8206
rect 11004 7642 11060 7654
rect 11004 7590 11006 7642
rect 11058 7590 11060 7642
rect 11228 7634 11284 7644
rect 10556 6850 10612 6860
rect 10780 7501 10836 7513
rect 10780 7449 10782 7501
rect 10834 7449 10836 7501
rect 10780 6804 10836 7449
rect 10780 6738 10836 6748
rect 9996 6524 10164 6580
rect 9996 6356 10052 6366
rect 9996 5906 10052 6300
rect 9996 5854 9998 5906
rect 10050 5854 10052 5906
rect 9996 5842 10052 5854
rect 9716 5628 9940 5684
rect 10108 5738 10164 6524
rect 10332 6578 10388 6590
rect 10332 6526 10334 6578
rect 10386 6526 10388 6578
rect 10108 5686 10110 5738
rect 10162 5686 10164 5738
rect 10108 5674 10164 5686
rect 10220 6020 10276 6030
rect 9716 5346 9772 5628
rect 9716 5294 9718 5346
rect 9770 5294 9772 5346
rect 9716 5282 9772 5294
rect 9996 5348 10052 5358
rect 10220 5348 10276 5964
rect 10332 5908 10388 6526
rect 11004 5908 11060 7590
rect 11116 7476 11172 7486
rect 11340 7476 11396 9774
rect 11900 9826 11956 11116
rect 11900 9774 11902 9826
rect 11954 9774 11956 9826
rect 11900 9762 11956 9774
rect 12012 11174 12014 11226
rect 12066 11174 12068 11226
rect 11564 9658 11620 9670
rect 11564 9606 11566 9658
rect 11618 9606 11620 9658
rect 11564 9044 11620 9606
rect 12012 9492 12068 11174
rect 12572 10836 12628 11228
rect 13524 11284 13580 11294
rect 13524 11190 13580 11228
rect 12572 10770 12628 10780
rect 13132 10498 13188 10510
rect 13132 10446 13134 10498
rect 13186 10446 13188 10498
rect 12236 10276 12292 10286
rect 12236 9811 12292 10220
rect 12348 9940 12404 9950
rect 12348 9846 12404 9884
rect 12236 9759 12238 9811
rect 12290 9759 12292 9811
rect 12236 9747 12292 9759
rect 12012 9436 12628 9492
rect 11564 8978 11620 8988
rect 12572 8428 12628 9436
rect 12796 9044 12852 9054
rect 12796 8950 12852 8988
rect 13132 8428 13188 10446
rect 12460 8372 12628 8428
rect 12796 8372 12852 8382
rect 12908 8372 13188 8428
rect 13580 9828 13636 9838
rect 13692 9828 13748 12908
rect 14028 12178 14084 12908
rect 14476 12962 14532 12974
rect 14476 12910 14478 12962
rect 14530 12910 14532 12962
rect 14476 12292 14532 12910
rect 14476 12226 14532 12236
rect 14028 12126 14030 12178
rect 14082 12126 14084 12178
rect 14028 12114 14084 12126
rect 14812 12068 14868 12078
rect 14812 11974 14868 12012
rect 13916 11620 13972 11630
rect 13804 11396 13860 11406
rect 13804 11302 13860 11340
rect 13916 11394 13972 11564
rect 14588 11620 14644 11630
rect 14252 11508 14308 11518
rect 14252 11414 14308 11452
rect 13916 11342 13918 11394
rect 13970 11342 13972 11394
rect 13916 11330 13972 11342
rect 14364 11396 14420 11406
rect 14364 11327 14366 11340
rect 14418 11327 14420 11340
rect 14588 11394 14644 11564
rect 15932 11518 15988 15820
rect 16492 15426 16548 16046
rect 17164 16100 17220 16110
rect 17164 16006 17220 16044
rect 17836 15876 17892 16868
rect 16492 15374 16494 15426
rect 16546 15374 16548 15426
rect 16492 14532 16548 15374
rect 17612 15820 17892 15876
rect 17948 16884 18004 16894
rect 17948 15876 18004 16828
rect 18172 16882 18228 16894
rect 18172 16830 18174 16882
rect 18226 16830 18228 16882
rect 18844 16882 18900 16894
rect 18172 16660 18228 16830
rect 18564 16826 18620 16838
rect 18172 16594 18228 16604
rect 18396 16770 18452 16782
rect 18396 16718 18398 16770
rect 18450 16718 18452 16770
rect 18396 16436 18452 16718
rect 18564 16774 18566 16826
rect 18618 16774 18620 16826
rect 18564 16436 18620 16774
rect 18844 16830 18846 16882
rect 18898 16830 18900 16882
rect 18844 16660 18900 16830
rect 18844 16594 18900 16604
rect 18956 16882 19012 16894
rect 18956 16830 18958 16882
rect 19010 16830 19012 16882
rect 18564 16380 18900 16436
rect 18396 16370 18452 16380
rect 17948 15820 18284 15876
rect 17612 15370 17668 15820
rect 17612 15318 17614 15370
rect 17666 15318 17668 15370
rect 18228 15370 18284 15820
rect 16492 14466 16548 14476
rect 16604 14530 16660 14542
rect 16604 14478 16606 14530
rect 16658 14478 16660 14530
rect 17276 14532 17332 14542
rect 17500 14532 17556 14542
rect 16156 14420 16212 14430
rect 16156 14326 16212 14364
rect 16604 13972 16660 14478
rect 16940 14474 16996 14486
rect 16492 13916 16660 13972
rect 16716 14420 16772 14430
rect 16492 13802 16548 13916
rect 16492 13750 16494 13802
rect 16546 13750 16548 13802
rect 16324 13524 16380 13534
rect 16324 13430 16380 13468
rect 16380 13076 16436 13086
rect 16492 13076 16548 13750
rect 16604 13748 16660 13758
rect 16716 13748 16772 14364
rect 16940 14422 16942 14474
rect 16994 14422 16996 14474
rect 17276 14438 17332 14476
rect 17388 14476 17500 14532
rect 16940 14420 16996 14422
rect 16940 14354 16996 14364
rect 17388 14362 17444 14476
rect 17500 14466 17556 14476
rect 17388 14310 17390 14362
rect 17442 14310 17444 14362
rect 17388 14298 17444 14310
rect 17612 13972 17668 15318
rect 16604 13746 16772 13748
rect 16604 13694 16606 13746
rect 16658 13694 16772 13746
rect 16604 13692 16772 13694
rect 16828 13860 16884 13870
rect 17612 13860 17668 13916
rect 16604 13682 16660 13692
rect 16828 13636 16884 13804
rect 16772 13580 16884 13636
rect 17500 13804 17668 13860
rect 17836 15314 17892 15326
rect 17836 15262 17838 15314
rect 17890 15262 17892 15314
rect 18228 15318 18230 15370
rect 18282 15318 18284 15370
rect 18228 15306 18284 15318
rect 17836 13860 17892 15262
rect 18060 15204 18116 15242
rect 18060 15138 18116 15148
rect 18620 15204 18676 15214
rect 18396 14532 18452 14542
rect 18396 14438 18452 14476
rect 18620 14530 18676 15148
rect 18844 15202 18900 16380
rect 18844 15150 18846 15202
rect 18898 15150 18900 15202
rect 18844 15138 18900 15150
rect 18620 14478 18622 14530
rect 18674 14478 18676 14530
rect 18620 14466 18676 14478
rect 18956 14644 19012 16830
rect 19102 16868 19104 16920
rect 19156 16868 19158 16920
rect 19102 16660 19158 16868
rect 19516 16884 19572 16894
rect 19516 16770 19572 16828
rect 19516 16718 19518 16770
rect 19570 16718 19572 16770
rect 19516 16706 19572 16718
rect 19102 16604 19236 16660
rect 19068 16436 19124 16446
rect 19068 16210 19124 16380
rect 19068 16158 19070 16210
rect 19122 16158 19124 16210
rect 19068 16146 19124 16158
rect 19180 15876 19236 16604
rect 19516 16212 19572 16222
rect 19180 15820 19274 15876
rect 19218 15352 19274 15820
rect 19218 15316 19220 15352
rect 19272 15316 19274 15352
rect 19218 15222 19274 15260
rect 19404 15314 19460 15326
rect 19404 15262 19406 15314
rect 19458 15262 19460 15314
rect 18116 14420 18172 14430
rect 18116 14326 18172 14364
rect 16772 13578 16828 13580
rect 16772 13526 16774 13578
rect 16826 13526 16828 13578
rect 16772 13514 16828 13526
rect 16380 13074 16548 13076
rect 16380 13022 16382 13074
rect 16434 13022 16548 13074
rect 16380 13020 16548 13022
rect 16380 13010 16436 13020
rect 17500 12924 17556 13804
rect 17836 13746 17892 13804
rect 17836 13694 17838 13746
rect 17890 13694 17892 13746
rect 17836 13682 17892 13694
rect 17948 13748 18004 13758
rect 17948 13654 18004 13692
rect 18116 13746 18172 13758
rect 18116 13694 18118 13746
rect 18170 13694 18172 13746
rect 17500 12872 17502 12924
rect 17554 12872 17556 12924
rect 17836 13524 17892 13534
rect 17836 12962 17892 13468
rect 18116 13412 18172 13694
rect 18956 13748 19012 14588
rect 19292 15092 19348 15102
rect 19068 14532 19124 14542
rect 19068 14450 19070 14476
rect 19122 14450 19124 14476
rect 19292 14530 19348 15036
rect 19404 14644 19460 15262
rect 19516 15314 19572 16156
rect 19628 15540 19684 18956
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19796 18676 19852 18686
rect 20188 18676 20244 19852
rect 19796 18674 20244 18676
rect 19796 18622 19798 18674
rect 19850 18622 20244 18674
rect 19796 18620 20244 18622
rect 19796 18610 19852 18620
rect 20244 18452 20300 18462
rect 20412 18452 20468 19964
rect 20524 18564 20580 20524
rect 20692 20514 20748 20524
rect 22428 20356 22484 20750
rect 22428 20290 22484 20300
rect 22540 21026 22820 21028
rect 22540 20974 22766 21026
rect 22818 20974 22820 21026
rect 22540 20972 22820 20974
rect 21028 20020 21084 20030
rect 21028 19926 21084 19964
rect 21868 20020 21924 20058
rect 21868 19954 21924 19964
rect 22204 20018 22260 20030
rect 22204 19966 22206 20018
rect 22258 19966 22260 20018
rect 21476 19908 21532 19918
rect 21476 19814 21532 19852
rect 21868 19850 21924 19862
rect 21868 19798 21870 19850
rect 21922 19798 21924 19850
rect 20860 19236 20916 19246
rect 20860 19142 20916 19180
rect 21196 19236 21252 19246
rect 21196 19142 21252 19180
rect 20524 18498 20580 18508
rect 20916 18788 20972 18798
rect 20244 18450 20468 18452
rect 20244 18398 20246 18450
rect 20298 18398 20468 18450
rect 20244 18396 20468 18398
rect 20748 18452 20804 18462
rect 20244 18386 20300 18396
rect 20748 18358 20804 18396
rect 20916 18282 20972 18732
rect 20916 18230 20918 18282
rect 20970 18230 20972 18282
rect 21532 18450 21588 18462
rect 21532 18398 21534 18450
rect 21586 18398 21588 18450
rect 21532 18340 21588 18398
rect 21868 18452 21924 19798
rect 21980 19234 22036 19246
rect 21980 19182 21982 19234
rect 22034 19182 22036 19234
rect 21980 18788 22036 19182
rect 22204 18900 22260 19966
rect 22540 20018 22596 20972
rect 22764 20962 22820 20972
rect 23100 21476 23156 21486
rect 23100 20916 23156 21420
rect 23100 20802 23156 20860
rect 23100 20750 23102 20802
rect 23154 20750 23156 20802
rect 23100 20738 23156 20750
rect 23436 20804 23492 20814
rect 23436 20580 23492 20748
rect 23324 20578 23492 20580
rect 23324 20526 23438 20578
rect 23490 20526 23492 20578
rect 23324 20524 23492 20526
rect 22540 19966 22542 20018
rect 22594 19966 22596 20018
rect 22540 19908 22596 19966
rect 22540 19842 22596 19852
rect 22876 20020 22932 20030
rect 22876 19794 22932 19964
rect 22876 19742 22878 19794
rect 22930 19742 22932 19794
rect 22876 19572 22932 19742
rect 22876 19516 23156 19572
rect 23100 19012 23156 19516
rect 22652 18956 23156 19012
rect 23212 19124 23268 19134
rect 22204 18844 22596 18900
rect 21980 18722 22036 18732
rect 22272 18564 22328 18574
rect 22272 18488 22328 18508
rect 22272 18436 22274 18488
rect 22326 18436 22328 18488
rect 22272 18424 22328 18436
rect 22540 18450 22596 18844
rect 21868 18386 21924 18396
rect 22540 18398 22542 18450
rect 22594 18398 22596 18450
rect 22540 18340 22596 18398
rect 21532 18274 21588 18284
rect 21756 18282 21812 18294
rect 20916 18218 20972 18230
rect 21756 18230 21758 18282
rect 21810 18230 21812 18282
rect 22540 18274 22596 18284
rect 21420 17780 21476 17790
rect 21308 17612 21364 17622
rect 20972 17610 21364 17612
rect 20860 17556 20916 17566
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20076 16882 20132 16894
rect 20076 16830 20078 16882
rect 20130 16830 20132 16882
rect 20076 16436 20132 16830
rect 20860 16770 20916 17500
rect 20860 16718 20862 16770
rect 20914 16718 20916 16770
rect 20860 16706 20916 16718
rect 20972 17558 21310 17610
rect 21362 17558 21364 17610
rect 20972 17556 21364 17558
rect 20972 16436 21028 17556
rect 21308 17546 21364 17556
rect 21420 17610 21476 17724
rect 21420 17558 21422 17610
rect 21474 17558 21476 17610
rect 21420 17220 21476 17558
rect 19852 16380 20132 16436
rect 20692 16380 21028 16436
rect 21084 17164 21476 17220
rect 19852 16098 19908 16380
rect 20692 16322 20804 16380
rect 20132 16266 20188 16278
rect 20132 16214 20134 16266
rect 20186 16214 20188 16266
rect 20692 16270 20694 16322
rect 20746 16270 20804 16322
rect 20692 16258 20804 16270
rect 20132 16212 20188 16214
rect 20132 16146 20188 16156
rect 19852 16046 19854 16098
rect 19906 16046 19908 16098
rect 19852 15876 19908 16046
rect 19964 16100 20020 16110
rect 19964 16025 19966 16044
rect 20018 16025 20020 16044
rect 19964 16006 20020 16025
rect 19852 15820 20244 15876
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20020 15540 20076 15550
rect 19628 15484 20020 15540
rect 20020 15446 20076 15484
rect 19516 15262 19518 15314
rect 19570 15262 19572 15314
rect 19516 15204 19572 15262
rect 19516 15138 19572 15148
rect 20076 14644 20132 14654
rect 19404 14578 19460 14588
rect 19684 14642 20132 14644
rect 19684 14590 20078 14642
rect 20130 14590 20132 14642
rect 19684 14588 20132 14590
rect 19292 14478 19294 14530
rect 19346 14478 19348 14530
rect 19292 14466 19348 14478
rect 19684 14530 19740 14588
rect 20076 14578 20132 14588
rect 19684 14478 19686 14530
rect 19738 14478 19740 14530
rect 19684 14466 19740 14478
rect 19068 14438 19124 14450
rect 19516 14418 19572 14430
rect 19516 14366 19518 14418
rect 19570 14366 19572 14418
rect 19068 13972 19124 13982
rect 19068 13878 19124 13916
rect 19516 13860 19572 14366
rect 20188 14308 20244 15820
rect 20300 15540 20356 15550
rect 20300 15341 20356 15484
rect 20300 15289 20302 15341
rect 20354 15289 20356 15341
rect 20300 15277 20356 15289
rect 20524 15316 20580 15326
rect 20524 15148 20580 15260
rect 20470 15092 20580 15148
rect 20470 14530 20526 15092
rect 20470 14478 20472 14530
rect 20524 14478 20526 14530
rect 20470 14466 20526 14478
rect 20636 14644 20692 14654
rect 20636 14530 20692 14588
rect 20636 14478 20638 14530
rect 20690 14478 20692 14530
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19516 13794 19572 13804
rect 18956 13682 19012 13692
rect 19404 13746 19460 13758
rect 19404 13694 19406 13746
rect 19458 13694 19460 13746
rect 18508 13524 18564 13534
rect 18116 13346 18172 13356
rect 18228 13522 18564 13524
rect 18228 13470 18510 13522
rect 18562 13470 18564 13522
rect 18228 13468 18564 13470
rect 18060 13076 18116 13086
rect 18060 12982 18116 13020
rect 18228 13018 18284 13468
rect 18508 13458 18564 13468
rect 18620 13524 18676 13534
rect 18620 13188 18676 13468
rect 19404 13524 19460 13694
rect 19740 13748 19796 13758
rect 19740 13654 19796 13692
rect 20188 13748 20244 14252
rect 20188 13682 20244 13692
rect 20524 13860 20580 13870
rect 20524 13746 20580 13804
rect 20524 13694 20526 13746
rect 20578 13694 20580 13746
rect 20524 13682 20580 13694
rect 20300 13636 20356 13646
rect 19404 13458 19460 13468
rect 19628 13524 19684 13534
rect 17836 12910 17838 12962
rect 17890 12910 17892 12962
rect 18228 12966 18230 13018
rect 18282 12966 18284 13018
rect 18228 12954 18284 12966
rect 18508 13132 18676 13188
rect 18788 13412 18844 13422
rect 18508 12962 18564 13132
rect 17836 12898 17892 12910
rect 18508 12910 18510 12962
rect 18562 12910 18564 12962
rect 18508 12898 18564 12910
rect 18620 12964 18676 12974
rect 17500 12234 17556 12872
rect 17500 12182 17502 12234
rect 17554 12182 17556 12234
rect 18060 12292 18116 12302
rect 18060 12198 18116 12236
rect 18228 12292 18284 12302
rect 18228 12234 18284 12236
rect 17500 12170 17556 12182
rect 17836 12180 17892 12190
rect 17724 12124 17836 12180
rect 18228 12182 18230 12234
rect 18282 12182 18284 12234
rect 18228 12170 18284 12182
rect 18508 12180 18564 12190
rect 16716 12066 16772 12078
rect 16716 12014 16718 12066
rect 16770 12014 16772 12066
rect 15876 11506 15988 11518
rect 15876 11454 15878 11506
rect 15930 11454 15988 11506
rect 15876 11442 15988 11454
rect 14588 11342 14590 11394
rect 14642 11342 14644 11394
rect 14588 11330 14644 11342
rect 14364 11302 14420 11327
rect 13916 10612 13972 10622
rect 14028 10612 14084 10622
rect 13916 10610 14084 10612
rect 13916 10558 13918 10610
rect 13970 10558 14030 10610
rect 14082 10558 14084 10610
rect 13916 10556 14084 10558
rect 13916 10546 13972 10556
rect 13580 9826 13748 9828
rect 13580 9774 13582 9826
rect 13634 9774 13748 9826
rect 13580 9772 13748 9774
rect 13580 9042 13636 9772
rect 13580 8990 13582 9042
rect 13634 8990 13636 9042
rect 13580 8428 13636 8990
rect 14028 9044 14084 10556
rect 14812 10500 14868 10510
rect 14812 10406 14868 10444
rect 15932 10164 15988 11442
rect 16324 11508 16380 11518
rect 16324 11414 16380 11452
rect 16716 11396 16772 12014
rect 16940 11508 16996 11518
rect 16828 11396 16884 11406
rect 16716 11394 16884 11396
rect 16716 11342 16830 11394
rect 16882 11342 16884 11394
rect 16716 11340 16884 11342
rect 16828 11330 16884 11340
rect 16940 11394 16996 11452
rect 16940 11342 16942 11394
rect 16994 11342 16996 11394
rect 16940 11330 16996 11342
rect 17612 11396 17668 11406
rect 17724 11396 17780 12124
rect 17836 12086 17892 12124
rect 18508 12086 18564 12124
rect 18620 12178 18676 12908
rect 18788 12906 18844 13356
rect 19180 13074 19236 13086
rect 19180 13022 19182 13074
rect 19234 13022 19236 13074
rect 18788 12854 18790 12906
rect 18842 12854 18844 12906
rect 18788 12292 18844 12854
rect 19068 12964 19124 12974
rect 18788 12236 18862 12292
rect 18620 12126 18622 12178
rect 18674 12126 18676 12178
rect 18620 12114 18676 12126
rect 18806 12215 18862 12236
rect 18806 12163 18808 12215
rect 18860 12163 18862 12215
rect 18806 12068 18862 12163
rect 18806 12012 18900 12068
rect 18116 11844 18172 11854
rect 18116 11618 18172 11788
rect 18116 11566 18118 11618
rect 18170 11566 18172 11618
rect 18116 11554 18172 11566
rect 18284 11620 18340 11630
rect 17612 11394 17780 11396
rect 17612 11342 17614 11394
rect 17666 11342 17780 11394
rect 17612 11340 17780 11342
rect 17836 11394 17892 11406
rect 17836 11342 17838 11394
rect 17890 11342 17892 11394
rect 16660 11172 16716 11182
rect 16660 11078 16716 11116
rect 17276 11170 17332 11182
rect 17276 11118 17278 11170
rect 17330 11118 17332 11170
rect 17276 10836 17332 11118
rect 17612 11172 17668 11340
rect 17612 11106 17668 11116
rect 17276 10770 17332 10780
rect 17556 10724 17612 10734
rect 17556 10666 17612 10668
rect 17556 10614 17558 10666
rect 17610 10614 17612 10666
rect 17556 10602 17612 10614
rect 16716 10498 16772 10510
rect 16716 10446 16718 10498
rect 16770 10446 16772 10498
rect 15932 10108 16324 10164
rect 14364 9826 14420 9838
rect 14364 9774 14366 9826
rect 14418 9774 14420 9826
rect 14364 9044 14420 9774
rect 15148 9826 15204 9838
rect 15148 9774 15150 9826
rect 15202 9774 15204 9826
rect 14028 9042 14420 9044
rect 14028 8990 14030 9042
rect 14082 8990 14420 9042
rect 14028 8988 14420 8990
rect 14812 9716 14868 9726
rect 14812 9042 14868 9660
rect 15148 9268 15204 9774
rect 16268 9604 16324 10108
rect 16716 9828 16772 10446
rect 17724 10500 17780 10510
rect 17724 10406 17780 10444
rect 16716 9762 16772 9772
rect 17724 9828 17780 9838
rect 15148 9202 15204 9212
rect 16156 9548 16324 9604
rect 17052 9714 17108 9726
rect 17052 9662 17054 9714
rect 17106 9662 17108 9714
rect 17052 9604 17108 9662
rect 14812 8990 14814 9042
rect 14866 8990 14868 9042
rect 13580 8372 13972 8428
rect 12348 8260 12404 8270
rect 12348 8166 12404 8204
rect 12460 8258 12516 8372
rect 12796 8370 12964 8372
rect 12796 8318 12798 8370
rect 12850 8318 12964 8370
rect 12796 8316 12964 8318
rect 12796 8306 12852 8316
rect 12460 8206 12462 8258
rect 12514 8206 12516 8258
rect 12460 8194 12516 8206
rect 12180 8036 12236 8046
rect 12180 8034 12628 8036
rect 12180 7982 12182 8034
rect 12234 7982 12628 8034
rect 12180 7980 12628 7982
rect 12180 7970 12236 7980
rect 11844 7588 11900 7598
rect 11844 7494 11900 7532
rect 12292 7588 12348 7598
rect 12292 7494 12348 7532
rect 11116 7474 11396 7476
rect 11116 7422 11118 7474
rect 11170 7422 11396 7474
rect 11116 7420 11396 7422
rect 12572 7474 12628 7980
rect 12572 7422 12574 7474
rect 12626 7422 12628 7474
rect 13448 7588 13504 7598
rect 13448 7530 13504 7532
rect 13448 7478 13450 7530
rect 13502 7478 13504 7530
rect 13448 7466 13504 7478
rect 11116 7364 11172 7420
rect 12572 7410 12628 7422
rect 11116 7298 11172 7308
rect 13580 7252 13636 8372
rect 13916 8258 13972 8372
rect 13916 8206 13918 8258
rect 13970 8206 13972 8258
rect 13916 8194 13972 8206
rect 14028 7474 14084 8988
rect 14812 8978 14868 8990
rect 14028 7422 14030 7474
rect 14082 7422 14084 7474
rect 13356 7196 13636 7252
rect 13692 7250 13748 7262
rect 13692 7198 13694 7250
rect 13746 7198 13748 7250
rect 12236 6804 12292 6814
rect 12236 6710 12292 6748
rect 13020 6692 13076 6702
rect 13356 6692 13412 7196
rect 13692 6804 13748 7198
rect 13692 6738 13748 6748
rect 13020 6690 13412 6692
rect 13020 6638 13022 6690
rect 13074 6638 13358 6690
rect 13410 6638 13412 6690
rect 13020 6636 13412 6638
rect 13020 6626 13076 6636
rect 13356 6626 13412 6636
rect 11452 6468 11508 6478
rect 11452 6130 11508 6412
rect 11452 6078 11454 6130
rect 11506 6078 11508 6130
rect 11452 6066 11508 6078
rect 11116 5908 11172 5918
rect 11004 5906 11172 5908
rect 11004 5854 11118 5906
rect 11170 5854 11172 5906
rect 11004 5852 11172 5854
rect 10332 5814 10388 5852
rect 11116 5842 11172 5852
rect 10332 5348 10388 5358
rect 10220 5346 10388 5348
rect 10220 5294 10334 5346
rect 10386 5294 10388 5346
rect 10220 5292 10388 5294
rect 9436 5070 9438 5122
rect 9490 5070 9492 5122
rect 9436 5058 9492 5070
rect 9996 5122 10052 5292
rect 10332 5282 10388 5292
rect 9996 5070 9998 5122
rect 10050 5070 10052 5122
rect 9996 5058 10052 5070
rect 14028 5124 14084 7422
rect 14812 8596 14868 8606
rect 14812 7474 14868 8540
rect 16156 8260 16212 9548
rect 17052 9538 17108 9548
rect 17724 9492 17780 9772
rect 17836 9658 17892 11342
rect 18284 10666 18340 11564
rect 17948 10612 18004 10622
rect 17948 10518 18004 10556
rect 18284 10614 18286 10666
rect 18338 10614 18340 10666
rect 18620 11506 18676 11518
rect 18620 11454 18622 11506
rect 18674 11454 18676 11506
rect 18620 10724 18676 11454
rect 18844 11396 18900 12012
rect 19068 11844 19124 12908
rect 19180 12292 19236 13022
rect 19628 12404 19684 13468
rect 19964 12964 20020 12974
rect 19964 12870 20020 12908
rect 20300 12962 20356 13580
rect 20636 13188 20692 14478
rect 20748 14530 20804 16258
rect 20860 16098 20916 16110
rect 20860 16046 20862 16098
rect 20914 16046 20916 16098
rect 20860 15540 20916 16046
rect 20860 15474 20916 15484
rect 20748 14478 20750 14530
rect 20802 14478 20804 14530
rect 20748 14466 20804 14478
rect 21084 14532 21140 17164
rect 21756 17108 21812 18230
rect 22148 17610 22204 17622
rect 21980 17556 22036 17566
rect 21980 17462 22036 17500
rect 22148 17558 22150 17610
rect 22202 17558 22204 17610
rect 22148 17108 22204 17558
rect 21756 17042 21812 17052
rect 21980 17052 22204 17108
rect 21980 16548 22036 17052
rect 21532 16492 22036 16548
rect 22092 16884 22148 16894
rect 21532 16322 21588 16492
rect 21532 16270 21534 16322
rect 21586 16270 21588 16322
rect 21532 16258 21588 16270
rect 22092 16098 22148 16828
rect 21926 16042 21982 16054
rect 21926 15990 21928 16042
rect 21980 15990 21982 16042
rect 22092 16046 22094 16098
rect 22146 16046 22148 16098
rect 22092 16034 22148 16046
rect 22204 16100 22260 16110
rect 22204 16006 22260 16044
rect 21926 15988 21982 15990
rect 21926 15932 22036 15988
rect 21980 15316 22036 15932
rect 21980 15250 22036 15260
rect 22428 15540 22484 15550
rect 22428 15316 22484 15484
rect 21084 14084 21140 14476
rect 21644 14502 21700 14514
rect 21644 14450 21646 14502
rect 21698 14450 21700 14502
rect 21644 14308 21700 14450
rect 21644 14242 21700 14252
rect 21084 14018 21140 14028
rect 22428 13858 22484 15260
rect 22540 15314 22596 15326
rect 22540 15262 22542 15314
rect 22594 15262 22596 15314
rect 22540 14308 22596 15262
rect 22540 14242 22596 14252
rect 22428 13806 22430 13858
rect 22482 13806 22484 13858
rect 22428 13794 22484 13806
rect 21756 13748 21812 13758
rect 21420 13188 21476 13198
rect 20636 13186 21476 13188
rect 20636 13134 21422 13186
rect 21474 13134 21476 13186
rect 20636 13132 21476 13134
rect 21420 13122 21476 13132
rect 21756 12964 21812 13692
rect 20300 12910 20302 12962
rect 20354 12910 20356 12962
rect 20300 12898 20356 12910
rect 21308 12962 21812 12964
rect 21308 12910 21758 12962
rect 21810 12910 21812 12962
rect 21308 12908 21812 12910
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19628 12348 19908 12404
rect 19180 12226 19236 12236
rect 19572 12178 19628 12190
rect 19572 12126 19574 12178
rect 19626 12126 19628 12178
rect 19180 12068 19236 12078
rect 19572 12068 19628 12126
rect 19180 12066 19628 12068
rect 19180 12014 19182 12066
rect 19234 12014 19628 12066
rect 19180 12012 19628 12014
rect 19740 12068 19796 12078
rect 19180 12002 19236 12012
rect 19740 11974 19796 12012
rect 19852 11844 19908 12348
rect 19068 11788 19236 11844
rect 19014 11396 19070 11406
rect 18844 11340 19014 11396
rect 19014 11302 19070 11340
rect 19180 11394 19236 11788
rect 19628 11788 19908 11844
rect 20188 12206 20244 12218
rect 20188 12154 20190 12206
rect 20242 12154 20244 12206
rect 19180 11342 19182 11394
rect 19234 11342 19236 11394
rect 19180 11172 19236 11342
rect 18620 10658 18676 10668
rect 18844 11116 19236 11172
rect 19292 11732 19348 11742
rect 19292 11394 19348 11676
rect 19292 11342 19294 11394
rect 19346 11342 19348 11394
rect 18060 10500 18116 10510
rect 18116 10444 18228 10500
rect 18060 10434 18116 10444
rect 17836 9606 17838 9658
rect 17890 9606 17892 9658
rect 17836 9594 17892 9606
rect 18060 9770 18116 9782
rect 18060 9718 18062 9770
rect 18114 9718 18116 9770
rect 18060 9604 18116 9718
rect 17724 9436 18004 9492
rect 17276 9042 17332 9054
rect 17276 8990 17278 9042
rect 17330 8990 17332 9042
rect 16716 8932 16772 8942
rect 16716 8838 16772 8876
rect 16156 8178 16158 8204
rect 16210 8178 16212 8204
rect 16156 8166 16212 8178
rect 14812 7422 14814 7474
rect 14866 7422 14868 7474
rect 14812 7410 14868 7422
rect 16044 8148 16100 8158
rect 14140 6804 14196 6814
rect 14140 6710 14196 6748
rect 16044 6578 16100 8092
rect 16716 7362 16772 7374
rect 16716 7310 16718 7362
rect 16770 7310 16772 7362
rect 16044 6526 16046 6578
rect 16098 6526 16100 6578
rect 16044 6468 16100 6526
rect 16044 6402 16100 6412
rect 16604 6690 16660 6702
rect 16604 6638 16606 6690
rect 16658 6638 16660 6690
rect 16604 6356 16660 6638
rect 16716 6692 16772 7310
rect 17164 6690 17220 6702
rect 16716 6626 16772 6636
rect 16940 6634 16996 6646
rect 16940 6582 16942 6634
rect 16994 6582 16996 6634
rect 16940 6356 16996 6582
rect 17164 6638 17166 6690
rect 17218 6638 17220 6690
rect 17164 6580 17220 6638
rect 17164 6514 17220 6524
rect 17276 6522 17332 8990
rect 17948 9042 18004 9436
rect 17948 8990 17950 9042
rect 18002 8990 18004 9042
rect 17948 8978 18004 8990
rect 18060 9044 18116 9548
rect 18060 8978 18116 8988
rect 18172 8830 18228 10444
rect 18284 10164 18340 10614
rect 18284 10098 18340 10108
rect 18732 10612 18788 10622
rect 17612 8818 17668 8830
rect 17612 8766 17614 8818
rect 17666 8766 17668 8818
rect 17612 8596 17668 8766
rect 18116 8818 18228 8830
rect 18116 8766 18118 8818
rect 18170 8766 18228 8818
rect 18116 8764 18228 8766
rect 18284 9826 18340 9838
rect 18284 9774 18286 9826
rect 18338 9774 18340 9826
rect 18284 8932 18340 9774
rect 18732 9156 18788 10556
rect 18844 10610 18900 11116
rect 18844 10558 18846 10610
rect 18898 10558 18900 10610
rect 19002 10836 19058 10846
rect 19002 10660 19058 10780
rect 19002 10608 19004 10660
rect 19056 10608 19058 10660
rect 19002 10596 19058 10608
rect 19180 10612 19236 10622
rect 18844 10546 18900 10558
rect 18732 9090 18788 9100
rect 18956 10164 19012 10174
rect 18956 9788 19012 10108
rect 18956 9736 18958 9788
rect 19010 9736 19012 9788
rect 18956 9098 19012 9736
rect 18956 9046 18958 9098
rect 19010 9046 19012 9098
rect 18956 9034 19012 9046
rect 19180 9044 19236 10556
rect 19292 10500 19348 11342
rect 19628 11396 19684 11788
rect 20188 11732 20244 12154
rect 21308 12178 21364 12908
rect 21756 12898 21812 12908
rect 22428 13524 22484 13534
rect 22428 12962 22484 13468
rect 22652 13188 22708 18956
rect 23212 18564 23268 19068
rect 23212 18450 23268 18508
rect 23212 18398 23214 18450
rect 23266 18398 23268 18450
rect 23212 18386 23268 18398
rect 23324 18452 23380 20524
rect 23436 20514 23492 20524
rect 23548 20692 23604 22988
rect 24444 22932 24500 22942
rect 23996 22930 24500 22932
rect 23996 22878 24446 22930
rect 24498 22878 24500 22930
rect 23996 22876 24500 22878
rect 23996 22482 24052 22876
rect 24444 22866 24500 22876
rect 24556 22708 24612 23884
rect 24780 23156 24836 23166
rect 24780 23062 24836 23100
rect 23996 22430 23998 22482
rect 24050 22430 24052 22482
rect 23996 22418 24052 22430
rect 24220 22652 24612 22708
rect 23884 22372 23940 22382
rect 23660 21924 23716 21934
rect 23660 21586 23716 21868
rect 23660 21534 23662 21586
rect 23714 21534 23716 21586
rect 23660 21522 23716 21534
rect 23884 21474 23940 22316
rect 23996 21812 24052 21822
rect 23996 21630 24052 21756
rect 23996 21578 23998 21630
rect 24050 21578 24052 21630
rect 23996 21566 24052 21578
rect 23884 21422 23886 21474
rect 23938 21422 23940 21474
rect 23884 21410 23940 21422
rect 24108 21028 24164 21038
rect 23772 20916 23828 20926
rect 23772 20802 23828 20860
rect 23772 20750 23774 20802
rect 23826 20750 23828 20802
rect 23772 20738 23828 20750
rect 23548 20254 23604 20636
rect 24108 20356 24164 20972
rect 24220 20580 24276 22652
rect 25116 21924 25172 24670
rect 25228 24052 25284 26236
rect 25340 25620 25396 25630
rect 25452 25620 25508 26796
rect 25900 26628 25956 29148
rect 26236 28868 26292 29148
rect 26236 28802 26292 28812
rect 26124 28644 26180 28654
rect 26012 28586 26068 28598
rect 26012 28534 26014 28586
rect 26066 28534 26068 28586
rect 26012 28532 26068 28534
rect 26012 28466 26068 28476
rect 26124 27186 26180 28588
rect 26124 27134 26126 27186
rect 26178 27134 26180 27186
rect 26124 27122 26180 27134
rect 26236 28586 26292 28598
rect 26236 28534 26238 28586
rect 26290 28534 26292 28586
rect 26236 28532 26292 28534
rect 26012 26964 26068 26974
rect 26012 26852 26124 26908
rect 25900 26562 25956 26572
rect 25788 26404 25844 26414
rect 25788 26346 25844 26348
rect 25620 26325 25676 26337
rect 25620 26273 25622 26325
rect 25674 26292 25676 26325
rect 25788 26294 25790 26346
rect 25842 26294 25844 26346
rect 26068 26402 26124 26852
rect 26068 26350 26070 26402
rect 26122 26350 26124 26402
rect 26068 26338 26124 26350
rect 25674 26273 25732 26292
rect 25788 26282 25844 26294
rect 25620 26236 25732 26273
rect 25676 26180 25732 26236
rect 26236 26180 26292 28476
rect 25676 26124 26292 26180
rect 26348 25732 26404 32732
rect 26572 32452 26628 32462
rect 26572 31890 26628 32396
rect 26796 32228 26852 32732
rect 26796 32172 27132 32228
rect 26572 31838 26574 31890
rect 26626 31838 26628 31890
rect 26572 31826 26628 31838
rect 27076 31890 27132 32172
rect 27076 31838 27078 31890
rect 27130 31838 27132 31890
rect 27076 31826 27132 31838
rect 27356 31778 27412 31790
rect 27356 31726 27358 31778
rect 27410 31726 27412 31778
rect 26628 31332 26684 31342
rect 26460 30996 26516 31006
rect 26460 29482 26516 30940
rect 26628 30882 26684 31276
rect 26628 30830 26630 30882
rect 26682 30830 26684 30882
rect 26628 30324 26684 30830
rect 26628 30258 26684 30268
rect 26796 30994 26852 31006
rect 26796 30942 26798 30994
rect 26850 30942 26852 30994
rect 26460 29430 26462 29482
rect 26514 29430 26516 29482
rect 26460 29428 26516 29430
rect 26684 30100 26740 30110
rect 26684 29482 26740 30044
rect 26796 29540 26852 30942
rect 27356 30996 27412 31726
rect 27580 31780 27636 31790
rect 27580 31686 27636 31724
rect 27692 31052 27748 34188
rect 27916 32452 27972 32462
rect 27916 32358 27972 32396
rect 27860 32228 27916 32238
rect 27860 31890 27916 32172
rect 28028 31948 28084 36204
rect 28140 35812 28196 35822
rect 28252 35812 28308 36374
rect 28364 36426 28420 36438
rect 28364 36374 28366 36426
rect 28418 36374 28420 36426
rect 28364 36372 28420 36374
rect 28364 36306 28420 36316
rect 28252 35756 28420 35812
rect 28140 35598 28196 35756
rect 28140 35586 28252 35598
rect 28140 35534 28198 35586
rect 28250 35534 28252 35586
rect 28140 35532 28252 35534
rect 28196 35522 28252 35532
rect 28364 35476 28420 35756
rect 28364 35410 28420 35420
rect 28476 35700 28532 36540
rect 28924 35700 28980 37229
rect 29036 37268 29092 38780
rect 29036 37154 29092 37212
rect 29036 37102 29038 37154
rect 29090 37102 29092 37154
rect 29036 37090 29092 37102
rect 29036 35700 29092 35710
rect 28476 35026 28532 35644
rect 28476 34974 28478 35026
rect 28530 34974 28532 35026
rect 28476 34962 28532 34974
rect 28588 35698 29092 35700
rect 28588 35646 29038 35698
rect 29090 35646 29092 35698
rect 28588 35644 29092 35646
rect 28028 31892 28532 31948
rect 27860 31838 27862 31890
rect 27914 31838 27916 31890
rect 27860 31826 27916 31838
rect 28140 31778 28196 31790
rect 28140 31726 28142 31778
rect 28194 31726 28196 31778
rect 27692 30996 28084 31052
rect 27356 30930 27412 30940
rect 27748 30884 27804 30894
rect 27748 30790 27804 30828
rect 27132 30772 27188 30782
rect 27132 30770 27636 30772
rect 27132 30718 27134 30770
rect 27186 30718 27636 30770
rect 27132 30716 27636 30718
rect 27132 30706 27188 30716
rect 27580 30548 27636 30716
rect 27580 30492 27972 30548
rect 27916 30322 27972 30492
rect 27916 30270 27918 30322
rect 27970 30270 27972 30322
rect 27916 30258 27972 30270
rect 28028 30100 28084 30996
rect 28140 30436 28196 31726
rect 28364 31780 28420 31790
rect 28140 30380 28308 30436
rect 27692 30044 28084 30100
rect 28140 30212 28196 30222
rect 26964 29540 27020 29550
rect 26796 29538 27020 29540
rect 26796 29486 26966 29538
rect 27018 29486 27020 29538
rect 26796 29484 27020 29486
rect 26684 29430 26686 29482
rect 26738 29430 26740 29482
rect 26964 29474 27020 29484
rect 26460 29372 26628 29428
rect 26684 29418 26740 29430
rect 27524 29428 27580 29438
rect 26572 29316 26628 29372
rect 27524 29334 27580 29372
rect 26572 29260 26740 29316
rect 26460 29204 26516 29214
rect 26516 29148 26628 29204
rect 26460 29138 26516 29148
rect 26460 28868 26516 28878
rect 26460 28614 26516 28812
rect 26460 28562 26462 28614
rect 26514 28562 26516 28614
rect 26460 28550 26516 28562
rect 26572 28607 26628 29148
rect 26572 28555 26574 28607
rect 26626 28555 26628 28607
rect 26572 28543 26628 28555
rect 26684 28532 26740 29260
rect 26908 28980 26964 28990
rect 26796 28756 26852 28766
rect 26796 28642 26852 28700
rect 26796 28590 26798 28642
rect 26850 28590 26852 28642
rect 26796 28578 26852 28590
rect 26684 28466 26740 28476
rect 26796 28420 26852 28430
rect 26684 28308 26740 28318
rect 25340 25618 25508 25620
rect 25340 25566 25342 25618
rect 25394 25566 25508 25618
rect 25340 25564 25508 25566
rect 26012 25676 26404 25732
rect 26572 26066 26628 26078
rect 26572 26014 26574 26066
rect 26626 26014 26628 26066
rect 25340 25554 25396 25564
rect 25900 25060 25956 25070
rect 25228 23986 25284 23996
rect 25452 24948 25508 24958
rect 24332 21588 24388 21598
rect 24332 21586 24500 21588
rect 24332 21534 24334 21586
rect 24386 21534 24500 21586
rect 24332 21532 24500 21534
rect 24332 21522 24388 21532
rect 24444 20804 24500 21532
rect 24780 21140 24836 21150
rect 24780 21026 24836 21084
rect 24780 20974 24782 21026
rect 24834 20974 24836 21026
rect 24780 20962 24836 20974
rect 24444 20710 24500 20748
rect 24780 20804 24836 20814
rect 25116 20804 25172 21868
rect 25228 23716 25284 23726
rect 25228 21028 25284 23660
rect 25452 23390 25508 24892
rect 25900 24722 25956 25004
rect 25900 24670 25902 24722
rect 25954 24670 25956 24722
rect 25900 24658 25956 24670
rect 26012 24500 26068 25676
rect 26124 25508 26180 25518
rect 26124 25414 26180 25452
rect 26348 25508 26404 25518
rect 26348 25414 26404 25452
rect 26572 25060 26628 26014
rect 26572 24994 26628 25004
rect 26684 24948 26740 28252
rect 26796 25172 26852 28364
rect 26908 27074 26964 28924
rect 27692 28868 27748 30044
rect 27804 29876 27860 29886
rect 27804 29426 27860 29820
rect 27804 29374 27806 29426
rect 27858 29374 27860 29426
rect 27804 29362 27860 29374
rect 28028 29426 28084 29438
rect 28028 29374 28030 29426
rect 28082 29374 28084 29426
rect 27916 29316 27972 29326
rect 27692 28812 27860 28868
rect 27132 28644 27188 28654
rect 27132 28550 27188 28588
rect 27636 28644 27692 28654
rect 27636 28550 27692 28588
rect 27804 27300 27860 28812
rect 27916 28642 27972 29260
rect 28028 28756 28084 29374
rect 28140 29426 28196 30156
rect 28140 29374 28142 29426
rect 28194 29374 28196 29426
rect 28140 28980 28196 29374
rect 28140 28914 28196 28924
rect 28252 28868 28308 30380
rect 28364 29316 28420 31724
rect 28364 29250 28420 29260
rect 28252 28802 28308 28812
rect 28476 29204 28532 31892
rect 28588 31118 28644 35644
rect 29036 35634 29092 35644
rect 28700 35476 28756 35486
rect 28924 35476 28980 35486
rect 28700 35474 28924 35476
rect 28700 35422 28702 35474
rect 28754 35422 28924 35474
rect 28700 35420 28924 35422
rect 28700 35410 28756 35420
rect 28812 34468 28868 34478
rect 28812 34186 28868 34412
rect 28812 34134 28814 34186
rect 28866 34134 28868 34186
rect 28812 34122 28868 34134
rect 28924 34186 28980 35420
rect 28924 34134 28926 34186
rect 28978 34134 28980 34186
rect 28924 34122 28980 34134
rect 29036 34914 29092 34926
rect 29036 34862 29038 34914
rect 29090 34862 29092 34914
rect 28700 33348 28756 33358
rect 28700 32564 28756 33292
rect 29036 33348 29092 34862
rect 29148 34580 29204 41356
rect 29260 41186 29316 41198
rect 29260 41134 29262 41186
rect 29314 41134 29316 41186
rect 29260 41076 29316 41134
rect 29260 41010 29316 41020
rect 29260 40740 29316 40750
rect 29260 39058 29316 40684
rect 29372 40404 29428 43484
rect 29820 43540 29876 43550
rect 30156 43538 30212 44270
rect 29820 43446 29876 43484
rect 29988 43482 30044 43494
rect 29988 43430 29990 43482
rect 30042 43430 30044 43482
rect 29540 43092 29596 43102
rect 29540 42978 29596 43036
rect 29988 42980 30044 43430
rect 29540 42926 29542 42978
rect 29594 42926 29596 42978
rect 29540 42914 29596 42926
rect 29708 42924 30044 42980
rect 30156 43486 30158 43538
rect 30210 43486 30212 43538
rect 30156 42980 30212 43486
rect 30268 44324 30324 44334
rect 30268 43538 30324 44268
rect 30492 44324 30548 44334
rect 30492 44230 30548 44268
rect 30604 43652 30660 44438
rect 31164 44324 31220 44334
rect 31276 44324 31332 44828
rect 32228 44772 32284 45052
rect 32228 44706 32284 44716
rect 32396 44660 32452 46398
rect 32396 44594 32452 44604
rect 32620 46450 33180 46452
rect 32620 46398 33126 46450
rect 33178 46398 33180 46450
rect 32620 46396 33180 46398
rect 32620 44436 32676 46396
rect 33124 46386 33180 46396
rect 32956 45892 33012 45902
rect 32732 45778 32788 45790
rect 32732 45726 32734 45778
rect 32786 45726 32788 45778
rect 32732 45668 32788 45726
rect 32732 45602 32788 45612
rect 32956 45106 33012 45836
rect 33516 45892 33572 45902
rect 33516 45810 33518 45836
rect 33570 45810 33572 45836
rect 33516 45798 33572 45810
rect 32956 45054 32958 45106
rect 33010 45054 33012 45106
rect 32956 45042 33012 45054
rect 33628 44772 33684 46510
rect 33740 45892 33796 47182
rect 33740 45826 33796 45836
rect 33740 45108 33796 45118
rect 33852 45108 33908 47516
rect 35980 47570 36036 47582
rect 35980 47518 35982 47570
rect 36034 47518 36036 47570
rect 35196 47460 35252 47470
rect 35196 47378 35198 47404
rect 35250 47378 35252 47404
rect 35196 47366 35252 47378
rect 33740 45106 33908 45108
rect 33740 45054 33742 45106
rect 33794 45054 33908 45106
rect 33740 45052 33908 45054
rect 33964 47348 34020 47358
rect 33740 45042 33796 45052
rect 33292 44716 33684 44772
rect 33964 44772 34020 47292
rect 35420 47124 35476 47134
rect 35420 46452 35476 47068
rect 35532 46676 35588 46686
rect 35980 46676 36036 47518
rect 38836 47570 38892 47628
rect 38836 47518 38838 47570
rect 38890 47518 38892 47570
rect 38836 47506 38892 47518
rect 39284 47570 39340 48076
rect 44604 48132 44660 50200
rect 49308 48916 49364 48926
rect 44604 48066 44660 48076
rect 47292 48132 47348 48142
rect 39284 47518 39286 47570
rect 39338 47518 39340 47570
rect 39284 47506 39340 47518
rect 43372 48018 43428 48030
rect 43372 47966 43374 48018
rect 43426 47966 43428 48018
rect 36316 47458 36372 47470
rect 35532 46674 36036 46676
rect 35532 46622 35534 46674
rect 35586 46622 36036 46674
rect 35532 46620 36036 46622
rect 36092 47414 36148 47426
rect 36092 47362 36094 47414
rect 36146 47362 36148 47414
rect 35532 46610 35588 46620
rect 35420 46396 35812 46452
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 34860 45780 34916 45790
rect 34392 44772 34448 44782
rect 33964 44716 34244 44772
rect 32060 44380 32676 44436
rect 31164 44322 31332 44324
rect 31164 44270 31166 44322
rect 31218 44270 31332 44322
rect 31724 44324 31780 44334
rect 32060 44324 32116 44380
rect 31164 44268 31332 44270
rect 31164 44258 31220 44268
rect 31388 44266 31444 44278
rect 31388 44214 31390 44266
rect 31442 44214 31444 44266
rect 30996 44100 31052 44110
rect 31388 44100 31444 44214
rect 31556 44266 31612 44278
rect 31556 44214 31558 44266
rect 31610 44214 31612 44266
rect 31724 44242 31726 44268
rect 31778 44242 31780 44268
rect 31724 44230 31780 44242
rect 32004 44287 32116 44324
rect 32004 44235 32006 44287
rect 32058 44268 32116 44287
rect 32620 44322 32676 44380
rect 32844 44660 32900 44670
rect 32620 44270 32622 44322
rect 32674 44270 32676 44322
rect 32058 44235 32060 44268
rect 32620 44258 32676 44270
rect 32732 44324 32788 44334
rect 32004 44223 32060 44235
rect 31556 44212 31612 44214
rect 31556 44156 31668 44212
rect 30996 44098 31444 44100
rect 30996 44046 30998 44098
rect 31050 44046 31444 44098
rect 30996 44044 31444 44046
rect 30996 44034 31052 44044
rect 30940 43652 30996 43662
rect 30604 43596 30772 43652
rect 30268 43486 30270 43538
rect 30322 43486 30324 43538
rect 30268 43474 30324 43486
rect 30548 43428 30604 43438
rect 30548 43334 30604 43372
rect 30324 42980 30380 42990
rect 30156 42978 30380 42980
rect 30156 42926 30326 42978
rect 30378 42926 30380 42978
rect 30156 42924 30380 42926
rect 29708 42420 29764 42924
rect 30324 42914 30380 42924
rect 30716 42868 30772 43596
rect 30716 42802 30772 42812
rect 29820 42754 29876 42766
rect 29820 42702 29822 42754
rect 29874 42702 29876 42754
rect 29820 42644 29876 42702
rect 30044 42756 30100 42766
rect 30044 42754 30212 42756
rect 30044 42702 30046 42754
rect 30098 42702 30212 42754
rect 30044 42700 30212 42702
rect 30044 42690 30100 42700
rect 29820 42578 29876 42588
rect 29540 42364 29764 42420
rect 29540 42082 29596 42364
rect 29540 42030 29542 42082
rect 29594 42030 29596 42082
rect 29540 42018 29596 42030
rect 30156 42084 30212 42700
rect 30716 42644 30772 42654
rect 30156 42028 30324 42084
rect 29764 42005 29820 42017
rect 29764 41972 29766 42005
rect 29708 41953 29766 41972
rect 29818 41953 29820 42005
rect 29708 41916 29820 41953
rect 30044 41998 30100 42010
rect 30044 41946 30046 41998
rect 30098 41972 30100 41998
rect 30268 41998 30324 42028
rect 30268 41972 30270 41998
rect 30322 41972 30324 41998
rect 30098 41946 30212 41972
rect 30044 41916 30212 41946
rect 29540 41300 29596 41310
rect 29540 41206 29596 41244
rect 29708 40852 29764 41916
rect 30156 41300 30212 41916
rect 30436 41986 30492 41998
rect 30436 41934 30438 41986
rect 30490 41972 30492 41986
rect 30716 41972 30772 42588
rect 30490 41970 30772 41972
rect 30490 41934 30718 41970
rect 30436 41918 30718 41934
rect 30770 41918 30772 41970
rect 30436 41916 30772 41918
rect 30268 41906 30324 41916
rect 30716 41906 30772 41916
rect 30828 41972 30884 41982
rect 30716 41748 30772 41758
rect 30212 41244 30548 41300
rect 30156 41206 30212 41244
rect 29372 40338 29428 40348
rect 29484 40796 29764 40852
rect 29820 41186 29876 41198
rect 29820 41134 29822 41186
rect 29874 41134 29876 41186
rect 29484 39842 29540 40796
rect 29820 40628 29876 41134
rect 30044 41186 30100 41198
rect 30044 41134 30046 41186
rect 30098 41134 30100 41186
rect 29820 40562 29876 40572
rect 29932 40852 29988 40862
rect 29932 40458 29988 40796
rect 29708 40404 29764 40414
rect 29932 40406 29934 40458
rect 29986 40406 29988 40458
rect 30044 40516 30100 41134
rect 30324 41076 30380 41086
rect 30044 40450 30100 40460
rect 30156 41020 30324 41076
rect 29932 40394 29988 40406
rect 29708 40310 29764 40348
rect 29484 39790 29486 39842
rect 29538 39790 29540 39842
rect 29484 39778 29540 39790
rect 29876 39620 29932 39630
rect 29876 39526 29932 39564
rect 30044 39620 30100 39630
rect 30044 39526 30100 39564
rect 30156 39618 30212 41020
rect 30324 40982 30380 41020
rect 30268 40628 30324 40638
rect 30268 40570 30324 40572
rect 30268 40518 30270 40570
rect 30322 40518 30324 40570
rect 30268 40506 30324 40518
rect 30156 39566 30158 39618
rect 30210 39566 30212 39618
rect 30156 39554 30212 39566
rect 30380 40402 30436 40414
rect 30380 40350 30382 40402
rect 30434 40350 30436 40402
rect 30380 39620 30436 40350
rect 30492 40180 30548 41244
rect 30492 40114 30548 40124
rect 30604 39786 30660 39798
rect 30604 39734 30606 39786
rect 30658 39734 30660 39786
rect 30492 39620 30548 39630
rect 30380 39618 30548 39620
rect 30380 39566 30494 39618
rect 30546 39566 30548 39618
rect 30380 39564 30548 39566
rect 29260 39006 29262 39058
rect 29314 39006 29316 39058
rect 29260 38948 29316 39006
rect 29932 39060 29988 39070
rect 29932 38966 29988 39004
rect 29260 38882 29316 38892
rect 29596 38834 29652 38846
rect 29596 38782 29598 38834
rect 29650 38782 29652 38834
rect 29596 38276 29652 38782
rect 30380 38668 30436 39564
rect 30492 39554 30548 39564
rect 30604 39620 30660 39734
rect 30604 39554 30660 39564
rect 30716 39396 30772 41692
rect 30828 40852 30884 41916
rect 30940 41802 30996 43596
rect 31164 43540 31220 43550
rect 31052 43538 31220 43540
rect 31052 43486 31166 43538
rect 31218 43486 31220 43538
rect 31052 43484 31220 43486
rect 31052 43092 31108 43484
rect 31164 43474 31220 43484
rect 31388 43316 31444 44044
rect 31500 43652 31556 43662
rect 31500 43538 31556 43596
rect 31500 43486 31502 43538
rect 31554 43486 31556 43538
rect 31500 43474 31556 43486
rect 31612 43540 31668 44156
rect 32228 44210 32284 44222
rect 32228 44158 32230 44210
rect 32282 44158 32284 44210
rect 31836 43764 31892 43774
rect 32228 43764 32284 44158
rect 31836 43594 31892 43708
rect 31836 43542 31838 43594
rect 31890 43542 31892 43594
rect 31612 43484 31780 43540
rect 31836 43530 31892 43542
rect 32060 43708 32284 43764
rect 31388 43260 31556 43316
rect 31052 43026 31108 43036
rect 31164 42980 31220 42990
rect 31164 42754 31220 42924
rect 31164 42702 31166 42754
rect 31218 42702 31220 42754
rect 31164 42690 31220 42702
rect 31388 42868 31444 42878
rect 31388 42715 31444 42812
rect 31388 42663 31390 42715
rect 31442 42663 31444 42715
rect 31388 42651 31444 42663
rect 31276 42586 31332 42598
rect 31276 42534 31278 42586
rect 31330 42534 31332 42586
rect 31052 41972 31108 41982
rect 31052 41878 31108 41916
rect 30940 41750 30942 41802
rect 30994 41750 30996 41802
rect 30940 41738 30996 41750
rect 31052 41636 31108 41646
rect 31108 41580 31220 41636
rect 31052 41570 31108 41580
rect 30828 40786 30884 40796
rect 30940 41186 30996 41198
rect 30940 41134 30942 41186
rect 30994 41134 30996 41186
rect 30940 40628 30996 41134
rect 30940 40562 30996 40572
rect 31052 41076 31108 41086
rect 31052 40402 31108 41020
rect 31164 40516 31220 41580
rect 31276 41186 31332 42534
rect 31500 41970 31556 43260
rect 31500 41918 31502 41970
rect 31554 41918 31556 41970
rect 31500 41906 31556 41918
rect 31724 41970 31780 43484
rect 31836 43426 31892 43438
rect 31836 43374 31838 43426
rect 31890 43374 31892 43426
rect 31836 42980 31892 43374
rect 31836 42914 31892 42924
rect 32060 43204 32116 43708
rect 32172 43540 32228 43550
rect 32172 43446 32228 43484
rect 31836 42756 31892 42766
rect 32060 42756 32116 43148
rect 32732 43092 32788 44268
rect 32844 43428 32900 44604
rect 33292 44324 33348 44716
rect 33516 44324 33572 44334
rect 33292 44322 33572 44324
rect 33292 44270 33518 44322
rect 33570 44270 33572 44322
rect 33292 44268 33572 44270
rect 33012 44212 33068 44222
rect 32956 44210 33068 44212
rect 32956 44158 33014 44210
rect 33066 44158 33068 44210
rect 32956 44146 33068 44158
rect 33516 44212 33572 44268
rect 33516 44146 33572 44156
rect 32956 43652 33012 44146
rect 32956 43586 33012 43596
rect 33404 43652 33460 43662
rect 33404 43558 33460 43596
rect 33068 43538 33124 43550
rect 33068 43486 33070 43538
rect 33122 43486 33124 43538
rect 33516 43538 33572 43550
rect 32844 43372 33012 43428
rect 32620 43036 32788 43092
rect 32620 42980 32676 43036
rect 32956 42980 33012 43372
rect 33068 43204 33124 43486
rect 33236 43482 33292 43494
rect 33236 43430 33238 43482
rect 33290 43430 33292 43482
rect 33236 43428 33292 43430
rect 33236 43362 33292 43372
rect 33516 43486 33518 43538
rect 33570 43486 33572 43538
rect 33068 43138 33124 43148
rect 33516 43092 33572 43486
rect 33516 43026 33572 43036
rect 33796 43314 33852 43326
rect 33796 43262 33798 43314
rect 33850 43262 33852 43314
rect 33180 42980 33236 42990
rect 32956 42924 33124 42980
rect 32620 42914 32676 42924
rect 32788 42868 32844 42878
rect 32788 42810 32844 42812
rect 31836 42754 32116 42756
rect 31836 42702 31838 42754
rect 31890 42702 32116 42754
rect 31836 42700 32116 42702
rect 32508 42754 32564 42766
rect 32508 42702 32510 42754
rect 32562 42702 32564 42754
rect 32788 42758 32790 42810
rect 32842 42758 32844 42810
rect 32788 42746 32844 42758
rect 32956 42756 33012 42766
rect 31836 42690 31892 42700
rect 32228 42644 32284 42654
rect 32228 42642 32452 42644
rect 32228 42590 32230 42642
rect 32282 42590 32452 42642
rect 32228 42588 32452 42590
rect 32228 42578 32284 42588
rect 31724 41918 31726 41970
rect 31778 41918 31780 41970
rect 31724 41748 31780 41918
rect 31724 41682 31780 41692
rect 31836 42532 31892 42542
rect 31836 41412 31892 42476
rect 32004 41746 32060 41758
rect 32004 41694 32006 41746
rect 32058 41694 32060 41746
rect 32004 41636 32060 41694
rect 32004 41570 32060 41580
rect 31388 41356 31780 41412
rect 31836 41356 32004 41412
rect 31388 41354 31444 41356
rect 31388 41302 31390 41354
rect 31442 41302 31444 41354
rect 31388 41290 31444 41302
rect 31612 41188 31668 41198
rect 31276 41134 31278 41186
rect 31330 41134 31332 41186
rect 31276 41122 31332 41134
rect 31388 41186 31668 41188
rect 31388 41134 31614 41186
rect 31666 41134 31668 41186
rect 31388 41132 31668 41134
rect 31724 41188 31780 41356
rect 31836 41188 31892 41198
rect 31724 41186 31892 41188
rect 31724 41134 31838 41186
rect 31890 41134 31892 41186
rect 31724 41132 31892 41134
rect 31164 40460 31276 40516
rect 31052 40350 31054 40402
rect 31106 40350 31108 40402
rect 31220 40458 31276 40460
rect 31220 40406 31222 40458
rect 31274 40406 31276 40458
rect 31220 40394 31276 40406
rect 31052 40338 31108 40350
rect 31276 40292 31332 40302
rect 31388 40292 31444 41132
rect 31612 41122 31668 41132
rect 31836 41122 31892 41132
rect 31948 40964 32004 41356
rect 32396 41300 32452 42588
rect 32508 42532 32564 42702
rect 32956 42662 33012 42700
rect 32508 42466 32564 42476
rect 32620 42642 32676 42654
rect 32620 42590 32622 42642
rect 32674 42590 32676 42642
rect 32620 41636 32676 42590
rect 33068 42532 33124 42924
rect 32620 41570 32676 41580
rect 32956 42476 33124 42532
rect 32396 41244 32900 41300
rect 32116 41076 32172 41086
rect 32116 41074 32788 41076
rect 32116 41022 32118 41074
rect 32170 41022 32788 41074
rect 32116 41020 32788 41022
rect 32116 41010 32172 41020
rect 31724 40908 32004 40964
rect 31612 40404 31668 40414
rect 31724 40404 31780 40908
rect 32060 40852 32116 40862
rect 31948 40404 32004 40414
rect 31612 40402 31780 40404
rect 31612 40350 31614 40402
rect 31666 40350 31780 40402
rect 31612 40348 31780 40350
rect 31836 40402 32004 40404
rect 31836 40350 31950 40402
rect 32002 40350 32004 40402
rect 31836 40348 32004 40350
rect 31612 40338 31668 40348
rect 31276 40290 31444 40292
rect 31276 40238 31278 40290
rect 31330 40238 31444 40290
rect 31276 40236 31444 40238
rect 31276 40226 31332 40236
rect 31612 40180 31668 40190
rect 30940 39900 31444 39956
rect 30828 39620 30884 39630
rect 30940 39620 30996 39900
rect 30828 39618 30996 39620
rect 30828 39566 30830 39618
rect 30882 39566 30996 39618
rect 30828 39564 30996 39566
rect 30828 39554 30884 39564
rect 29596 38210 29652 38220
rect 30100 38612 30436 38668
rect 30492 39340 30772 39396
rect 30100 38274 30156 38612
rect 30100 38222 30102 38274
rect 30154 38222 30156 38274
rect 30100 38210 30156 38222
rect 30268 38500 30324 38510
rect 29260 38164 29316 38174
rect 29260 38015 29316 38108
rect 29260 37963 29262 38015
rect 29314 37963 29316 38015
rect 29596 38052 29652 38062
rect 29260 37951 29316 37963
rect 29372 37994 29428 38006
rect 29372 37942 29374 37994
rect 29426 37942 29428 37994
rect 29596 37970 29598 37996
rect 29650 37970 29652 37996
rect 29596 37958 29652 37970
rect 29820 37994 29876 38006
rect 29372 37940 29428 37942
rect 29372 37874 29428 37884
rect 29820 37942 29822 37994
rect 29874 37942 29876 37994
rect 29820 37828 29876 37942
rect 29820 37762 29876 37772
rect 29260 37268 29316 37278
rect 29260 37174 29316 37212
rect 29820 37268 29876 37278
rect 29596 37042 29652 37054
rect 29596 36990 29598 37042
rect 29650 36990 29652 37042
rect 29596 36484 29652 36990
rect 29316 36372 29372 36382
rect 29316 36278 29372 36316
rect 29596 35754 29652 36428
rect 29260 35733 29316 35745
rect 29260 35681 29262 35733
rect 29314 35681 29316 35733
rect 29260 35588 29316 35681
rect 29260 35028 29316 35532
rect 29372 35726 29428 35738
rect 29372 35674 29374 35726
rect 29426 35674 29428 35726
rect 29372 35476 29428 35674
rect 29372 35410 29428 35420
rect 29596 35702 29598 35754
rect 29650 35702 29652 35754
rect 29260 34972 29540 35028
rect 29372 34804 29428 34814
rect 29148 34524 29316 34580
rect 29148 34356 29204 34366
rect 29148 34186 29204 34300
rect 29148 34134 29150 34186
rect 29202 34134 29204 34186
rect 29148 34122 29204 34134
rect 29036 33282 29092 33292
rect 29260 32676 29316 34524
rect 29372 34186 29428 34748
rect 29372 34134 29374 34186
rect 29426 34134 29428 34186
rect 29372 34122 29428 34134
rect 29260 32610 29316 32620
rect 29148 32564 29204 32574
rect 28700 32562 29204 32564
rect 28700 32510 28702 32562
rect 28754 32510 29150 32562
rect 29202 32510 29204 32562
rect 28700 32508 29204 32510
rect 28700 32498 28756 32508
rect 28812 31780 28868 32508
rect 29148 32498 29204 32508
rect 29036 31780 29092 31790
rect 28812 31778 29092 31780
rect 28812 31726 29038 31778
rect 29090 31726 29092 31778
rect 28812 31724 29092 31726
rect 28588 31106 28700 31118
rect 28588 31054 28646 31106
rect 28698 31054 28700 31106
rect 28588 31052 28700 31054
rect 28644 31042 28700 31052
rect 28588 30884 28644 30894
rect 28588 29652 28644 30828
rect 28700 30212 28756 30222
rect 28812 30212 28868 31724
rect 29036 31714 29092 31724
rect 29484 31332 29540 34972
rect 29596 34356 29652 35702
rect 29820 36594 29876 37212
rect 29820 36542 29822 36594
rect 29874 36542 29876 36594
rect 29820 35754 29876 36542
rect 30156 37266 30212 37278
rect 30156 37214 30158 37266
rect 30210 37214 30212 37266
rect 30156 35822 30212 37214
rect 29820 35702 29822 35754
rect 29874 35702 29876 35754
rect 30100 35810 30212 35822
rect 30100 35758 30102 35810
rect 30154 35758 30212 35810
rect 30100 35756 30212 35758
rect 30100 35746 30156 35756
rect 29820 35690 29876 35702
rect 30268 35252 30324 38444
rect 30380 38050 30436 38062
rect 30380 37998 30382 38050
rect 30434 37998 30436 38050
rect 30380 37828 30436 37998
rect 30380 37762 30436 37772
rect 30492 37268 30548 39340
rect 30660 38890 30716 38902
rect 30660 38838 30662 38890
rect 30714 38838 30716 38890
rect 30660 38836 30716 38838
rect 30660 38780 30772 38836
rect 30604 38052 30660 38062
rect 30716 38052 30772 38780
rect 30828 38834 30884 38846
rect 30828 38782 30830 38834
rect 30882 38782 30884 38834
rect 30828 38500 30884 38782
rect 30828 38434 30884 38444
rect 30940 38286 30996 39564
rect 31276 39786 31332 39798
rect 31276 39734 31278 39786
rect 31330 39734 31332 39786
rect 31276 39284 31332 39734
rect 31388 39618 31444 39900
rect 31388 39566 31390 39618
rect 31442 39566 31444 39618
rect 31388 39554 31444 39566
rect 31612 39618 31668 40124
rect 31612 39566 31614 39618
rect 31666 39566 31668 39618
rect 31612 39554 31668 39566
rect 31220 39228 31332 39284
rect 31220 38890 31276 39228
rect 31220 38838 31222 38890
rect 31274 38838 31276 38890
rect 31220 38826 31276 38838
rect 31612 39172 31668 39182
rect 31612 38890 31668 39116
rect 31612 38838 31614 38890
rect 31666 38838 31668 38890
rect 31612 38826 31668 38838
rect 31724 39060 31780 39070
rect 31724 38890 31780 39004
rect 31724 38838 31726 38890
rect 31778 38838 31780 38890
rect 31724 38826 31780 38838
rect 31052 38724 31108 38734
rect 31836 38724 31892 40348
rect 31948 40338 32004 40348
rect 32060 39508 32116 40796
rect 32172 39732 32228 39742
rect 32172 39730 32340 39732
rect 32172 39678 32174 39730
rect 32226 39678 32340 39730
rect 32172 39676 32340 39678
rect 32172 39666 32228 39676
rect 32060 39452 32228 39508
rect 31948 38948 32004 38958
rect 31948 38890 32004 38892
rect 31948 38838 31950 38890
rect 32002 38838 32004 38890
rect 31948 38826 32004 38838
rect 32172 38862 32228 39452
rect 32172 38836 32174 38862
rect 32226 38836 32228 38862
rect 32172 38770 32228 38780
rect 31052 38722 31892 38724
rect 31052 38670 31054 38722
rect 31106 38670 31892 38722
rect 31052 38668 31892 38670
rect 31052 38658 31108 38668
rect 31780 38500 31836 38510
rect 30884 38274 30996 38286
rect 30884 38222 30886 38274
rect 30938 38222 30996 38274
rect 30884 38220 30996 38222
rect 31612 38388 31668 38398
rect 30884 38210 30940 38220
rect 31052 38108 31556 38164
rect 31052 38052 31108 38108
rect 30716 37996 31108 38052
rect 30604 37492 30660 37996
rect 31500 37994 31556 38108
rect 31332 37940 31388 37950
rect 31332 37882 31388 37884
rect 31332 37830 31334 37882
rect 31386 37830 31388 37882
rect 31332 37818 31388 37830
rect 31500 37942 31502 37994
rect 31554 37942 31556 37994
rect 31612 38050 31668 38332
rect 31780 38274 31836 38444
rect 31780 38222 31782 38274
rect 31834 38222 31836 38274
rect 31780 38210 31836 38222
rect 32172 38276 32228 38286
rect 31612 37998 31614 38050
rect 31666 37998 31668 38050
rect 31612 37986 31668 37998
rect 30996 37492 31052 37502
rect 30604 37490 31052 37492
rect 30604 37438 30998 37490
rect 31050 37438 31052 37490
rect 30604 37436 31052 37438
rect 30996 37426 31052 37436
rect 30828 37268 30884 37278
rect 30492 37212 30660 37268
rect 30492 37042 30548 37054
rect 30492 36990 30494 37042
rect 30546 36990 30548 37042
rect 30380 36932 30436 36942
rect 30380 36036 30436 36876
rect 30492 36596 30548 36990
rect 30492 36530 30548 36540
rect 30604 36260 30660 37212
rect 30828 37174 30884 37212
rect 30604 36204 31444 36260
rect 30380 35970 30436 35980
rect 31220 36036 31276 36046
rect 31220 35922 31276 35980
rect 31220 35870 31222 35922
rect 31274 35870 31276 35922
rect 31220 35858 31276 35870
rect 30660 35588 30716 35598
rect 30660 35494 30716 35532
rect 30044 35196 30324 35252
rect 29596 34290 29652 34300
rect 29820 34914 29876 34926
rect 29820 34862 29822 34914
rect 29874 34862 29876 34914
rect 29820 34356 29876 34862
rect 30044 34692 30100 35196
rect 30044 34636 30436 34692
rect 29820 34290 29876 34300
rect 30044 34468 30100 34478
rect 29652 34132 29708 34142
rect 29932 34132 29988 34142
rect 29652 34130 29988 34132
rect 29652 34078 29654 34130
rect 29706 34078 29934 34130
rect 29986 34078 29988 34130
rect 29652 34076 29988 34078
rect 29652 34066 29708 34076
rect 29932 34066 29988 34076
rect 29708 33348 29764 33358
rect 29708 33254 29764 33292
rect 29820 32340 29876 32350
rect 29820 31890 29876 32284
rect 29820 31838 29822 31890
rect 29874 31838 29876 31890
rect 29820 31826 29876 31838
rect 29484 31266 29540 31276
rect 28756 30156 28868 30212
rect 28924 30994 28980 31006
rect 28924 30942 28926 30994
rect 28978 30942 28980 30994
rect 28700 30118 28756 30156
rect 28924 29876 28980 30942
rect 28924 29810 28980 29820
rect 29036 30996 29092 31006
rect 29036 29652 29092 30940
rect 30044 30884 30100 34412
rect 30268 34356 30324 34366
rect 30268 34262 30324 34300
rect 30380 32116 30436 34636
rect 31276 34130 31332 34142
rect 31276 34078 31278 34130
rect 31330 34078 31332 34130
rect 30940 33908 30996 33918
rect 30492 33906 30996 33908
rect 30492 33854 30942 33906
rect 30994 33854 30996 33906
rect 30492 33852 30996 33854
rect 30492 33458 30548 33852
rect 30940 33842 30996 33852
rect 31276 33684 31332 34078
rect 31388 33796 31444 36204
rect 31500 34804 31556 37942
rect 31892 37380 31948 37390
rect 31892 37286 31948 37324
rect 32060 37266 32116 37278
rect 32060 37214 32062 37266
rect 32114 37214 32116 37266
rect 32060 37044 32116 37214
rect 32060 36978 32116 36988
rect 31724 36596 31780 36606
rect 31724 36502 31780 36540
rect 31612 36148 31668 36158
rect 31612 35922 31668 36092
rect 31612 35870 31614 35922
rect 31666 35870 31668 35922
rect 31612 35858 31668 35870
rect 32060 36036 32116 36046
rect 31948 35698 32004 35710
rect 31948 35646 31950 35698
rect 32002 35646 32004 35698
rect 31948 35028 32004 35646
rect 32060 35698 32116 35980
rect 32060 35646 32062 35698
rect 32114 35646 32116 35698
rect 32060 35634 32116 35646
rect 31948 34962 32004 34972
rect 31500 34738 31556 34748
rect 31724 34804 31780 34814
rect 31724 34710 31780 34748
rect 31668 34468 31724 34478
rect 31668 34354 31724 34412
rect 31668 34302 31670 34354
rect 31722 34302 31724 34354
rect 31668 34290 31724 34302
rect 31388 33740 31780 33796
rect 31276 33628 31668 33684
rect 30492 33406 30494 33458
rect 30546 33406 30548 33458
rect 30492 33394 30548 33406
rect 31612 32788 31668 33628
rect 31612 32722 31668 32732
rect 31052 32676 31108 32686
rect 31052 32589 31108 32620
rect 31052 32537 31054 32589
rect 31106 32537 31108 32589
rect 31052 32525 31108 32537
rect 31612 32562 31668 32574
rect 30380 32050 30436 32060
rect 31612 32510 31614 32562
rect 31666 32510 31668 32562
rect 30380 31556 30436 31566
rect 30380 31220 30436 31500
rect 30380 31126 30436 31164
rect 31612 31118 31668 32510
rect 31724 31892 31780 33740
rect 31948 32340 32004 32350
rect 31948 32246 32004 32284
rect 32172 32340 32228 38220
rect 32172 32274 32228 32284
rect 32284 36708 32340 39676
rect 32732 39618 32788 41020
rect 32566 39562 32622 39574
rect 32566 39510 32568 39562
rect 32620 39510 32622 39562
rect 32732 39566 32734 39618
rect 32786 39566 32788 39618
rect 32732 39554 32788 39566
rect 32844 39618 32900 41244
rect 32844 39566 32846 39618
rect 32898 39566 32900 39618
rect 32844 39554 32900 39566
rect 32566 39284 32622 39510
rect 32622 39228 32676 39284
rect 32566 39218 32676 39228
rect 32452 38722 32508 38734
rect 32452 38670 32454 38722
rect 32506 38670 32508 38722
rect 32452 38668 32508 38670
rect 32452 38612 32564 38668
rect 32508 38052 32564 38612
rect 32508 37986 32564 37996
rect 32620 37828 32676 39218
rect 32956 38276 33012 42476
rect 33180 40964 33236 42924
rect 33796 42868 33852 43262
rect 33796 42802 33852 42812
rect 34076 42756 34132 42766
rect 34076 42662 34132 42700
rect 33740 41972 33796 41982
rect 34188 41972 34244 44716
rect 34392 44324 34448 44716
rect 34636 44548 34692 44558
rect 34860 44548 34916 45724
rect 35644 44994 35700 45006
rect 35644 44942 35646 44994
rect 35698 44942 35700 44994
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 34636 44546 34916 44548
rect 34636 44494 34638 44546
rect 34690 44494 34916 44546
rect 34636 44492 34916 44494
rect 34636 44482 34692 44492
rect 34392 44230 34448 44268
rect 35196 44324 35252 44334
rect 35196 44232 35198 44268
rect 35250 44232 35252 44268
rect 34748 44212 34804 44222
rect 35196 44220 35252 44232
rect 35532 44322 35588 44334
rect 35532 44270 35534 44322
rect 35586 44270 35588 44322
rect 34748 43594 34804 44156
rect 35532 44212 35588 44270
rect 35532 44146 35588 44156
rect 35644 43988 35700 44942
rect 35756 44434 35812 46396
rect 36092 45780 36148 47362
rect 36316 47406 36318 47458
rect 36370 47406 36372 47458
rect 36316 47236 36372 47406
rect 37324 47458 37380 47470
rect 37324 47406 37326 47458
rect 37378 47406 37380 47458
rect 36316 47170 36372 47180
rect 36932 47236 36988 47246
rect 36932 47142 36988 47180
rect 36316 46674 36372 46686
rect 36316 46622 36318 46674
rect 36370 46622 36372 46674
rect 36316 45892 36372 46622
rect 36652 46564 36708 46574
rect 36708 46508 36820 46564
rect 36652 46470 36708 46508
rect 36316 45826 36372 45836
rect 36092 45714 36148 45724
rect 36484 45666 36540 45678
rect 36484 45614 36486 45666
rect 36538 45614 36540 45666
rect 36484 45332 36540 45614
rect 36484 45266 36540 45276
rect 36316 45220 36372 45230
rect 36316 45162 36372 45164
rect 36204 45141 36260 45153
rect 36204 45089 36206 45141
rect 36258 45089 36260 45141
rect 36316 45110 36318 45162
rect 36370 45110 36372 45162
rect 36764 45162 36820 46508
rect 36876 45892 36932 45902
rect 36876 45798 36932 45836
rect 37324 45780 37380 47406
rect 38276 47460 38332 47470
rect 38276 47366 38332 47404
rect 39676 47458 39732 47470
rect 40460 47460 40516 47470
rect 39676 47406 39678 47458
rect 39730 47406 39732 47458
rect 37660 47236 37716 47246
rect 37436 47234 37716 47236
rect 37436 47182 37662 47234
rect 37714 47182 37716 47234
rect 37436 47180 37716 47182
rect 37436 46004 37492 47180
rect 37660 47170 37716 47180
rect 39340 46676 39396 46686
rect 39676 46676 39732 47406
rect 40236 47458 40516 47460
rect 40236 47406 40462 47458
rect 40514 47406 40516 47458
rect 40236 47404 40516 47406
rect 40236 46842 40292 47404
rect 40460 47394 40516 47404
rect 42812 47458 42868 47470
rect 42812 47406 42814 47458
rect 42866 47406 42868 47458
rect 41916 47348 41972 47358
rect 40236 46790 40238 46842
rect 40290 46790 40292 46842
rect 40236 46778 40292 46790
rect 40572 47124 40628 47134
rect 40236 46689 40292 46701
rect 39340 46674 39732 46676
rect 39340 46622 39342 46674
rect 39394 46622 39732 46674
rect 39340 46620 39732 46622
rect 39340 46610 39396 46620
rect 38556 46562 38612 46574
rect 38556 46510 38558 46562
rect 38610 46510 38612 46562
rect 38556 46228 38612 46510
rect 38556 46172 38836 46228
rect 37660 46004 37716 46014
rect 37436 46002 37716 46004
rect 37436 45950 37662 46002
rect 37714 45950 37716 46002
rect 37436 45948 37716 45950
rect 37660 45938 37716 45948
rect 37324 45724 37548 45780
rect 36316 45098 36372 45110
rect 36540 45134 36596 45146
rect 36204 44996 36260 45089
rect 36204 44930 36260 44940
rect 36540 45082 36542 45134
rect 36594 45082 36596 45134
rect 36764 45110 36766 45162
rect 36818 45110 36820 45162
rect 36764 45098 36820 45110
rect 36876 45332 36932 45342
rect 36540 44884 36596 45082
rect 36540 44548 36596 44828
rect 36540 44492 36708 44548
rect 35756 44382 35758 44434
rect 35810 44382 35812 44434
rect 35756 44370 35812 44382
rect 36092 44324 36148 44334
rect 35924 44322 36148 44324
rect 35924 44270 36094 44322
rect 36146 44270 36148 44322
rect 35924 44268 36148 44270
rect 35924 44266 35980 44268
rect 35924 44214 35926 44266
rect 35978 44214 35980 44266
rect 36092 44258 36148 44268
rect 35924 43988 35980 44214
rect 35532 43932 35980 43988
rect 36260 44098 36316 44110
rect 36260 44046 36262 44098
rect 36314 44046 36316 44098
rect 35532 43652 35588 43932
rect 34748 43542 34750 43594
rect 34802 43542 34804 43594
rect 35383 43596 35588 43652
rect 35383 43594 35439 43596
rect 34748 43530 34804 43542
rect 34972 43566 35028 43578
rect 34972 43514 34974 43566
rect 35026 43514 35028 43566
rect 35140 43573 35196 43585
rect 35140 43540 35142 43573
rect 34748 43428 34804 43438
rect 34468 43314 34524 43326
rect 34468 43262 34470 43314
rect 34522 43262 34524 43314
rect 34468 42868 34524 43262
rect 34468 42802 34524 42812
rect 34524 42698 34580 42710
rect 34524 42646 34526 42698
rect 34578 42646 34580 42698
rect 34524 42644 34580 42646
rect 34524 42578 34580 42588
rect 34748 42698 34804 43372
rect 34972 43316 35028 43514
rect 34972 43250 35028 43260
rect 35084 43521 35142 43540
rect 35194 43521 35196 43573
rect 35383 43542 35385 43594
rect 35437 43542 35439 43594
rect 35383 43530 35439 43542
rect 35644 43540 35700 43550
rect 35084 43484 35196 43521
rect 35084 42868 35140 43484
rect 35644 43370 35700 43484
rect 35532 43316 35588 43326
rect 35644 43318 35646 43370
rect 35698 43318 35700 43370
rect 35756 43538 35812 43550
rect 35756 43486 35758 43538
rect 35810 43486 35812 43538
rect 35756 43428 35812 43486
rect 35756 43362 35812 43372
rect 36092 43540 36148 43550
rect 36260 43540 36316 44046
rect 36092 43538 36316 43540
rect 36092 43486 36094 43538
rect 36146 43486 36316 43538
rect 36092 43484 36316 43486
rect 36428 43764 36484 43774
rect 35644 43306 35700 43318
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 34748 42646 34750 42698
rect 34802 42646 34804 42698
rect 34748 42420 34804 42646
rect 34748 42354 34804 42364
rect 34860 42812 35140 42868
rect 35308 42866 35364 42878
rect 35308 42814 35310 42866
rect 35362 42814 35364 42866
rect 34692 42196 34748 42206
rect 34860 42196 34916 42812
rect 35028 42698 35084 42710
rect 35028 42646 35030 42698
rect 35082 42646 35084 42698
rect 35028 42644 35084 42646
rect 35028 42578 35084 42588
rect 35308 42532 35364 42814
rect 35420 42868 35476 42878
rect 35420 42739 35476 42812
rect 35420 42687 35422 42739
rect 35474 42687 35476 42739
rect 35420 42675 35476 42687
rect 35532 42532 35588 43260
rect 35644 42868 35700 42878
rect 35644 42754 35700 42812
rect 35980 42756 36036 42766
rect 35644 42702 35646 42754
rect 35698 42702 35700 42754
rect 35644 42690 35700 42702
rect 35756 42754 36036 42756
rect 35756 42702 35982 42754
rect 36034 42702 36036 42754
rect 35756 42700 36036 42702
rect 35308 42466 35364 42476
rect 35420 42476 35588 42532
rect 34692 42194 34916 42196
rect 34692 42142 34694 42194
rect 34746 42142 34916 42194
rect 34692 42140 34916 42142
rect 34972 42420 35028 42430
rect 34692 42130 34748 42140
rect 33740 41970 33908 41972
rect 33740 41918 33742 41970
rect 33794 41918 33908 41970
rect 33740 41916 33908 41918
rect 33740 41906 33796 41916
rect 33292 41188 33348 41198
rect 33292 41094 33348 41132
rect 33628 41188 33684 41198
rect 33180 40908 33348 40964
rect 33068 40628 33124 40638
rect 33068 40458 33124 40572
rect 33068 40406 33070 40458
rect 33122 40406 33124 40458
rect 33068 40394 33124 40406
rect 33180 40430 33236 40442
rect 33180 40378 33182 40430
rect 33234 40378 33236 40430
rect 32956 38210 33012 38220
rect 33068 40292 33124 40302
rect 32956 38052 33012 38062
rect 32956 37958 33012 37996
rect 32788 37828 32844 37838
rect 32620 37826 32844 37828
rect 32620 37774 32790 37826
rect 32842 37774 32844 37826
rect 32620 37772 32844 37774
rect 32396 37380 32452 37390
rect 32396 37286 32452 37324
rect 32620 37044 32676 37772
rect 32788 37762 32844 37772
rect 32620 36978 32676 36988
rect 32284 32116 32340 36652
rect 33068 36596 33124 40236
rect 33180 39060 33236 40378
rect 33292 40292 33348 40908
rect 33628 40458 33684 41132
rect 33852 40526 33908 41916
rect 33964 41916 34244 41972
rect 34860 41972 34916 41982
rect 34972 41972 35028 42364
rect 34860 41970 35028 41972
rect 34860 41918 34862 41970
rect 34914 41918 35028 41970
rect 34860 41916 35028 41918
rect 33964 40740 34020 41916
rect 34860 41906 34916 41916
rect 34076 41746 34132 41758
rect 34076 41694 34078 41746
rect 34130 41694 34132 41746
rect 34076 41300 34132 41694
rect 34076 41234 34132 41244
rect 33964 40684 34132 40740
rect 33852 40514 33964 40526
rect 33852 40462 33910 40514
rect 33962 40462 33964 40514
rect 33852 40460 33964 40462
rect 33404 40430 33460 40442
rect 33404 40378 33406 40430
rect 33458 40404 33460 40430
rect 33628 40406 33630 40458
rect 33682 40406 33684 40458
rect 33908 40450 33964 40460
rect 33458 40378 33572 40404
rect 33628 40394 33684 40406
rect 33404 40348 33572 40378
rect 33292 40226 33348 40236
rect 33348 39394 33404 39406
rect 33348 39342 33350 39394
rect 33402 39342 33404 39394
rect 33348 39172 33404 39342
rect 33348 39106 33404 39116
rect 33180 38994 33236 39004
rect 33516 38948 33572 40348
rect 34076 40068 34132 40684
rect 34468 40628 34524 40638
rect 34468 40534 34524 40572
rect 34860 40404 34916 40414
rect 34860 40310 34916 40348
rect 34076 40002 34132 40012
rect 34972 39956 35028 41916
rect 35252 42308 35308 42318
rect 35252 41860 35308 42252
rect 35420 41860 35476 42476
rect 35756 42196 35812 42700
rect 35980 42690 36036 42700
rect 36092 42644 36148 43484
rect 36092 42578 36148 42588
rect 36316 42532 36372 42542
rect 36204 42530 36372 42532
rect 36204 42478 36318 42530
rect 36370 42478 36372 42530
rect 36204 42476 36372 42478
rect 35588 42140 35812 42196
rect 36092 42420 36148 42430
rect 35588 42082 35644 42140
rect 35588 42030 35590 42082
rect 35642 42030 35644 42082
rect 35588 42018 35644 42030
rect 35980 42084 36036 42094
rect 35868 41998 35924 42010
rect 35868 41946 35870 41998
rect 35922 41946 35924 41998
rect 35644 41860 35700 41870
rect 35420 41804 35588 41860
rect 35252 41766 35308 41804
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35196 41300 35252 41310
rect 35196 41206 35252 41244
rect 35196 40740 35252 40750
rect 35196 40404 35252 40684
rect 34860 39900 35028 39956
rect 35084 40402 35252 40404
rect 35084 40350 35198 40402
rect 35250 40350 35252 40402
rect 35084 40348 35252 40350
rect 34636 39620 34692 39630
rect 34356 39618 34692 39620
rect 34356 39566 34638 39618
rect 34690 39566 34692 39618
rect 34356 39564 34692 39566
rect 33796 39394 33852 39406
rect 33796 39342 33798 39394
rect 33850 39342 33852 39394
rect 33796 39284 33852 39342
rect 34356 39394 34412 39564
rect 34636 39554 34692 39564
rect 34356 39342 34358 39394
rect 34410 39342 34412 39394
rect 34356 39284 34412 39342
rect 34860 39396 34916 39900
rect 35084 39730 35140 40348
rect 35196 40338 35252 40348
rect 35308 40402 35364 40414
rect 35308 40350 35310 40402
rect 35362 40350 35364 40402
rect 35308 40292 35364 40350
rect 35308 40226 35364 40236
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35084 39678 35086 39730
rect 35138 39678 35140 39730
rect 35084 39666 35140 39678
rect 35420 39844 35476 39854
rect 34972 39620 35028 39630
rect 34972 39551 34974 39564
rect 35026 39551 35028 39564
rect 34972 39526 35028 39551
rect 35420 39620 35476 39788
rect 35420 39526 35476 39564
rect 34860 39340 35028 39396
rect 33796 39218 33852 39228
rect 33964 39228 34412 39284
rect 33516 38882 33572 38892
rect 33180 38836 33236 38846
rect 33180 38742 33236 38780
rect 33292 38724 33348 38734
rect 33292 38274 33348 38668
rect 33292 38222 33294 38274
rect 33346 38222 33348 38274
rect 33292 38210 33348 38222
rect 33740 38612 33796 38622
rect 33740 37604 33796 38556
rect 33964 38500 34020 39228
rect 33964 38434 34020 38444
rect 34860 38836 34916 38846
rect 34860 38286 34916 38780
rect 34804 38274 34916 38286
rect 34804 38222 34806 38274
rect 34858 38222 34916 38274
rect 34804 38220 34916 38222
rect 34972 38276 35028 39340
rect 35084 38724 35140 38762
rect 35084 38658 35140 38668
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 34972 38220 35252 38276
rect 34804 38210 34860 38220
rect 35084 38052 35140 38062
rect 34636 38050 35140 38052
rect 34636 37998 35086 38050
rect 35138 37998 35140 38050
rect 34636 37996 35140 37998
rect 33908 37828 33964 37838
rect 33908 37734 33964 37772
rect 34468 37826 34524 37838
rect 34468 37774 34470 37826
rect 34522 37774 34524 37826
rect 34468 37604 34524 37774
rect 33740 37548 34020 37604
rect 33292 37268 33348 37278
rect 33292 37174 33348 37212
rect 32620 36540 33124 36596
rect 33292 36932 33348 36942
rect 32508 36482 32564 36494
rect 32508 36430 32510 36482
rect 32562 36430 32564 36482
rect 32508 35924 32564 36430
rect 32508 35858 32564 35868
rect 32396 35474 32452 35486
rect 32396 35422 32398 35474
rect 32450 35422 32452 35474
rect 32396 35028 32452 35422
rect 32396 34962 32452 34972
rect 32452 34802 32508 34814
rect 32452 34750 32454 34802
rect 32506 34750 32508 34802
rect 32452 34244 32508 34750
rect 32452 34178 32508 34188
rect 32620 33572 32676 36540
rect 33180 36484 33236 36494
rect 33180 36390 33236 36428
rect 32844 36258 32900 36270
rect 32844 36206 32846 36258
rect 32898 36206 32900 36258
rect 32732 35700 32788 35710
rect 32844 35700 32900 36206
rect 32788 35644 32900 35700
rect 33180 35700 33236 35710
rect 32732 34914 32788 35644
rect 33180 35606 33236 35644
rect 33292 35530 33348 36876
rect 33852 36820 33908 36830
rect 33852 36370 33908 36764
rect 33852 36318 33854 36370
rect 33906 36318 33908 36370
rect 33628 36148 33684 36158
rect 33292 35478 33294 35530
rect 33346 35478 33348 35530
rect 33292 35466 33348 35478
rect 33404 35700 33460 35710
rect 32732 34862 32734 34914
rect 32786 34862 32788 34914
rect 32732 34850 32788 34862
rect 32956 35028 33012 35038
rect 32956 34914 33012 34972
rect 32956 34862 32958 34914
rect 33010 34862 33012 34914
rect 32956 34850 33012 34862
rect 33404 34914 33460 35644
rect 33516 35698 33572 35710
rect 33516 35646 33518 35698
rect 33570 35646 33572 35698
rect 33516 35028 33572 35646
rect 33516 34962 33572 34972
rect 33404 34862 33406 34914
rect 33458 34862 33460 34914
rect 33404 34850 33460 34862
rect 33516 34804 33572 34814
rect 33404 34692 33460 34702
rect 33404 34130 33460 34636
rect 33516 34580 33572 34748
rect 33628 34692 33684 36092
rect 33740 35028 33796 35038
rect 33740 34970 33796 34972
rect 33740 34918 33742 34970
rect 33794 34918 33796 34970
rect 33740 34906 33796 34918
rect 33852 34804 33908 36318
rect 33852 34738 33908 34748
rect 33628 34636 33796 34692
rect 33516 34524 33628 34580
rect 33404 34078 33406 34130
rect 33458 34078 33460 34130
rect 33572 34186 33628 34524
rect 33572 34134 33574 34186
rect 33626 34134 33628 34186
rect 33740 34242 33796 34636
rect 33852 34356 33908 34366
rect 33964 34356 34020 37548
rect 34468 37538 34524 37548
rect 34168 37380 34224 37390
rect 34168 37322 34224 37324
rect 34168 37270 34170 37322
rect 34222 37270 34224 37322
rect 34412 37380 34468 37390
rect 34636 37380 34692 37996
rect 35084 37986 35140 37996
rect 34412 37378 34692 37380
rect 34412 37326 34414 37378
rect 34466 37326 34692 37378
rect 34412 37324 34692 37326
rect 34412 37314 34468 37324
rect 34168 37258 34224 37270
rect 35196 37044 35252 38220
rect 35532 38164 35588 41804
rect 35644 41636 35700 41804
rect 35868 41860 35924 41946
rect 35868 41794 35924 41804
rect 35644 41570 35700 41580
rect 35980 41186 36036 42028
rect 36092 42026 36148 42364
rect 36092 41974 36094 42026
rect 36146 41974 36148 42026
rect 36092 41962 36148 41974
rect 36204 41972 36260 42476
rect 36316 42466 36372 42476
rect 36428 42308 36484 43708
rect 36316 42252 36484 42308
rect 36540 43538 36596 43550
rect 36540 43486 36542 43538
rect 36594 43486 36596 43538
rect 36316 42026 36372 42252
rect 36316 41974 36318 42026
rect 36370 41974 36372 42026
rect 36540 42084 36596 43486
rect 36652 42420 36708 44492
rect 36652 42354 36708 42364
rect 36316 41962 36372 41974
rect 36428 42005 36484 42017
rect 36204 41906 36260 41916
rect 36428 41953 36430 42005
rect 36482 41953 36484 42005
rect 35980 41134 35982 41186
rect 36034 41134 36036 41186
rect 35980 40292 36036 41134
rect 36428 41524 36484 41953
rect 36540 41972 36596 42028
rect 36652 41972 36708 41982
rect 36540 41970 36708 41972
rect 36540 41918 36654 41970
rect 36706 41918 36708 41970
rect 36540 41916 36708 41918
rect 36428 41188 36484 41468
rect 36652 41412 36708 41916
rect 36876 41748 36932 45276
rect 37492 45218 37548 45724
rect 38332 45332 38388 45342
rect 38780 45332 38836 46172
rect 39564 45778 39620 45790
rect 39564 45726 39566 45778
rect 39618 45726 39620 45778
rect 38892 45332 38948 45342
rect 38780 45330 38948 45332
rect 38780 45278 38894 45330
rect 38946 45278 38948 45330
rect 38780 45276 38948 45278
rect 37492 45166 37494 45218
rect 37546 45166 37548 45218
rect 37492 45154 37548 45166
rect 38220 45220 38276 45230
rect 38220 45162 38276 45164
rect 37772 45134 37828 45146
rect 37044 45108 37100 45118
rect 37044 45014 37100 45052
rect 37772 45082 37774 45134
rect 37826 45082 37828 45134
rect 37772 44772 37828 45082
rect 37996 45134 38052 45146
rect 37996 45082 37998 45134
rect 38050 45082 38052 45134
rect 37996 44884 38052 45082
rect 37996 44818 38052 44828
rect 38220 45110 38222 45162
rect 38274 45110 38276 45162
rect 37772 44706 37828 44716
rect 37996 44548 38052 44558
rect 37436 44546 38052 44548
rect 37436 44494 37998 44546
rect 38050 44494 38052 44546
rect 37436 44492 38052 44494
rect 36988 44434 37044 44446
rect 36988 44382 36990 44434
rect 37042 44382 37044 44434
rect 36988 42868 37044 44382
rect 37324 44322 37380 44334
rect 37100 44278 37156 44290
rect 37100 44226 37102 44278
rect 37154 44226 37156 44278
rect 37100 43988 37156 44226
rect 37324 44270 37326 44322
rect 37378 44270 37380 44322
rect 37324 44212 37380 44270
rect 37324 44146 37380 44156
rect 37100 43932 37268 43988
rect 36988 42802 37044 42812
rect 37100 43764 37156 43774
rect 37100 42726 37156 43708
rect 37212 43316 37268 43932
rect 37324 43540 37380 43550
rect 37436 43540 37492 44492
rect 37996 44482 38052 44492
rect 37660 44324 37716 44334
rect 37324 43538 37492 43540
rect 37324 43486 37326 43538
rect 37378 43486 37492 43538
rect 37324 43484 37492 43486
rect 37548 44322 37716 44324
rect 37548 44270 37662 44322
rect 37714 44270 37716 44322
rect 37548 44268 37716 44270
rect 37324 43474 37380 43484
rect 37212 43250 37268 43260
rect 37548 43204 37604 44268
rect 37660 44258 37716 44268
rect 38220 43764 38276 45110
rect 38332 45162 38388 45276
rect 38892 45266 38948 45276
rect 39564 45220 39620 45726
rect 38332 45110 38334 45162
rect 38386 45110 38388 45162
rect 39340 45164 39620 45220
rect 38332 45098 38388 45110
rect 38556 45108 38612 45118
rect 38556 45014 38612 45052
rect 38668 44884 38724 44894
rect 38556 44210 38612 44222
rect 38556 44158 38558 44210
rect 38610 44158 38612 44210
rect 38276 43708 38500 43764
rect 38220 43698 38276 43708
rect 37548 43148 37884 43204
rect 36876 41682 36932 41692
rect 36988 42698 37044 42710
rect 36988 42646 36990 42698
rect 37042 42646 37044 42698
rect 37100 42674 37102 42726
rect 37154 42674 37156 42726
rect 37548 42980 37604 42990
rect 37548 42726 37604 42924
rect 37828 42978 37884 43148
rect 37828 42926 37830 42978
rect 37882 42926 37884 42978
rect 37828 42914 37884 42926
rect 38444 42978 38500 43708
rect 38556 43540 38612 44158
rect 38556 43474 38612 43484
rect 38668 43316 38724 44828
rect 39340 44772 39396 45164
rect 39508 44994 39564 45006
rect 39508 44942 39510 44994
rect 39562 44942 39564 44994
rect 39508 44884 39564 44942
rect 39508 44818 39564 44828
rect 39340 43876 39396 44716
rect 39676 44660 39732 46620
rect 40012 46676 40068 46686
rect 40012 46582 40068 46620
rect 40236 46637 40238 46689
rect 40290 46637 40292 46689
rect 40236 46340 40292 46637
rect 40236 46284 40404 46340
rect 40348 46058 40404 46284
rect 40348 46006 40350 46058
rect 40402 46006 40404 46058
rect 40348 45994 40404 46006
rect 40460 45890 40516 45902
rect 40460 45838 40462 45890
rect 40514 45838 40516 45890
rect 40460 45780 40516 45838
rect 40460 45714 40516 45724
rect 40572 45444 40628 47068
rect 41356 46844 41804 46900
rect 40404 45388 40628 45444
rect 39956 45332 40012 45342
rect 39956 45238 40012 45276
rect 40404 45330 40460 45388
rect 40404 45278 40406 45330
rect 40458 45278 40460 45330
rect 40404 45266 40460 45278
rect 39676 44594 39732 44604
rect 40236 45108 40292 45118
rect 39340 43810 39396 43820
rect 40236 43708 40292 45052
rect 40460 44436 40516 44446
rect 40460 44342 40516 44380
rect 40124 43652 40292 43708
rect 40348 43652 40404 43662
rect 38444 42926 38446 42978
rect 38498 42926 38500 42978
rect 38444 42914 38500 42926
rect 38556 43260 38724 43316
rect 39228 43426 39284 43438
rect 39228 43374 39230 43426
rect 39282 43374 39284 43426
rect 37100 42662 37156 42674
rect 37324 42698 37380 42710
rect 36988 41636 37044 42646
rect 37324 42646 37326 42698
rect 37378 42646 37380 42698
rect 37548 42674 37550 42726
rect 37602 42674 37604 42726
rect 37548 42662 37604 42674
rect 38108 42756 38164 42766
rect 38108 42662 38164 42700
rect 37324 42420 37380 42646
rect 37324 42354 37380 42364
rect 37436 41972 37492 41982
rect 37436 41878 37492 41916
rect 36988 41570 37044 41580
rect 38220 41636 38276 41646
rect 36652 41356 37716 41412
rect 36428 41132 36540 41188
rect 36484 40962 36540 41132
rect 36484 40910 36486 40962
rect 36538 40910 36540 40962
rect 36484 40852 36540 40910
rect 37156 40962 37212 40974
rect 37156 40910 37158 40962
rect 37210 40910 37212 40962
rect 36484 40796 36708 40852
rect 36428 40628 36484 40638
rect 36428 40458 36484 40572
rect 36428 40406 36430 40458
rect 36482 40406 36484 40458
rect 36428 40394 36484 40406
rect 36540 40430 36596 40442
rect 35868 40236 35980 40292
rect 35756 39396 35812 39406
rect 35420 38108 35588 38164
rect 35644 39394 35812 39396
rect 35644 39342 35758 39394
rect 35810 39342 35812 39394
rect 35644 39340 35812 39342
rect 35644 38948 35700 39340
rect 35756 39330 35812 39340
rect 35308 38050 35364 38062
rect 35308 37998 35310 38050
rect 35362 37998 35364 38050
rect 35308 37156 35364 37998
rect 35308 37090 35364 37100
rect 35420 37044 35476 38108
rect 35644 38022 35700 38892
rect 35868 39060 35924 40236
rect 35980 40226 36036 40236
rect 36540 40378 36542 40430
rect 36594 40378 36596 40430
rect 36540 40180 36596 40378
rect 36540 40114 36596 40124
rect 36540 39620 36596 39630
rect 36540 39406 36596 39564
rect 36484 39394 36596 39406
rect 36484 39342 36486 39394
rect 36538 39342 36596 39394
rect 36484 39330 36596 39342
rect 35868 39004 36260 39060
rect 35868 38834 35924 39004
rect 35868 38782 35870 38834
rect 35922 38782 35924 38834
rect 35868 38770 35924 38782
rect 35980 38836 36036 38846
rect 35980 38742 36036 38780
rect 36092 38724 36148 38734
rect 35532 37994 35588 38006
rect 35532 37942 35534 37994
rect 35586 37942 35588 37994
rect 35644 37970 35646 38022
rect 35698 37970 35700 38022
rect 35644 37958 35700 37970
rect 35756 38612 35812 38622
rect 35532 37604 35588 37942
rect 35756 37828 35812 38556
rect 35980 38612 36148 38668
rect 35980 38052 36036 38612
rect 35924 38015 36036 38052
rect 35924 37963 35926 38015
rect 35978 37996 36036 38015
rect 35978 37963 35980 37996
rect 35924 37951 35980 37963
rect 36092 37994 36148 38006
rect 36092 37942 36094 37994
rect 36146 37942 36148 37994
rect 35756 37772 35924 37828
rect 35532 37538 35588 37548
rect 35756 37268 35812 37278
rect 35644 37266 35812 37268
rect 35644 37214 35758 37266
rect 35810 37214 35812 37266
rect 35644 37212 35812 37214
rect 35420 36988 35588 37044
rect 35196 36978 35252 36988
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35532 36148 35588 36988
rect 35532 36082 35588 36092
rect 35644 36484 35700 37212
rect 35756 37202 35812 37212
rect 35756 36596 35812 36606
rect 35868 36596 35924 37772
rect 36092 37380 36148 37942
rect 36204 37716 36260 39004
rect 36316 38612 36372 38622
rect 36316 38518 36372 38556
rect 36372 38052 36428 38062
rect 36372 37958 36428 37996
rect 36204 37660 36372 37716
rect 36092 37314 36148 37324
rect 36316 37268 36372 37660
rect 36428 37268 36484 37278
rect 36316 37266 36484 37268
rect 36316 37214 36430 37266
rect 36482 37214 36484 37266
rect 36316 37212 36484 37214
rect 36428 37202 36484 37212
rect 36148 37156 36204 37166
rect 36148 37062 36204 37100
rect 36540 36708 36596 39330
rect 35756 36594 35924 36596
rect 35756 36542 35758 36594
rect 35810 36542 35924 36594
rect 35756 36540 35924 36542
rect 36316 36652 36596 36708
rect 35756 36530 35812 36540
rect 35420 35924 35476 35934
rect 35644 35924 35700 36428
rect 35476 35868 35700 35924
rect 36204 36148 36260 36158
rect 35420 35830 35476 35868
rect 34412 35700 34468 35710
rect 34412 35698 35140 35700
rect 34412 35646 34414 35698
rect 34466 35646 35140 35698
rect 34412 35644 35140 35646
rect 34412 35634 34468 35644
rect 34076 35476 34132 35486
rect 34076 35474 34244 35476
rect 34076 35422 34078 35474
rect 34130 35422 34244 35474
rect 34076 35420 34244 35422
rect 34076 35410 34132 35420
rect 34076 35028 34132 35038
rect 34076 34934 34132 34972
rect 34076 34858 34132 34870
rect 34076 34806 34078 34858
rect 34130 34806 34132 34858
rect 34076 34804 34132 34806
rect 34076 34738 34132 34748
rect 33908 34300 34020 34356
rect 33852 34290 33908 34300
rect 34188 34244 34244 35420
rect 34412 35364 34468 35374
rect 34300 34914 34356 34926
rect 34300 34862 34302 34914
rect 34354 34862 34356 34914
rect 34300 34692 34356 34862
rect 34300 34626 34356 34636
rect 33740 34190 33742 34242
rect 33794 34190 33796 34242
rect 33740 34178 33796 34190
rect 33990 34188 34244 34244
rect 33572 34122 33628 34134
rect 33852 34130 33908 34142
rect 33404 34066 33460 34078
rect 33852 34078 33854 34130
rect 33906 34078 33908 34130
rect 33740 34020 33796 34030
rect 32396 33516 33348 33572
rect 32396 33458 32452 33516
rect 32396 33406 32398 33458
rect 32450 33406 32452 33458
rect 32396 33394 32452 33406
rect 33068 33348 33124 33358
rect 32956 33346 33124 33348
rect 32956 33294 33070 33346
rect 33122 33294 33124 33346
rect 32956 33292 33124 33294
rect 32564 32676 32620 32686
rect 32564 32582 32620 32620
rect 31948 32060 32340 32116
rect 32396 32340 32452 32350
rect 31724 31890 31892 31892
rect 31724 31838 31726 31890
rect 31778 31838 31892 31890
rect 31724 31836 31892 31838
rect 31724 31826 31780 31836
rect 31556 31106 31668 31118
rect 31556 31054 31558 31106
rect 31610 31054 31668 31106
rect 31556 31052 31668 31054
rect 31556 31042 31612 31052
rect 31836 31050 31892 31836
rect 30716 30996 30772 31006
rect 31108 30996 31164 31006
rect 30492 30994 31164 30996
rect 30492 30942 30718 30994
rect 30770 30942 31110 30994
rect 31162 30942 31164 30994
rect 31836 30998 31838 31050
rect 31890 30998 31892 31050
rect 31836 30986 31892 30998
rect 30492 30940 31164 30942
rect 30100 30828 30212 30884
rect 30044 30818 30100 30828
rect 28588 29586 28644 29596
rect 28812 29596 29092 29652
rect 28476 28980 28532 29148
rect 28812 29092 28868 29596
rect 28924 29316 28980 29326
rect 28924 29314 29092 29316
rect 28924 29262 28926 29314
rect 28978 29262 29092 29314
rect 28924 29260 29092 29262
rect 28924 29250 28980 29260
rect 28812 29036 28980 29092
rect 28476 28766 28532 28924
rect 28140 28756 28196 28766
rect 28028 28700 28140 28756
rect 28476 28754 28588 28766
rect 28476 28702 28534 28754
rect 28586 28702 28588 28754
rect 28476 28700 28588 28702
rect 27916 28590 27918 28642
rect 27970 28590 27972 28642
rect 27916 28578 27972 28590
rect 28140 28642 28196 28700
rect 28532 28690 28588 28700
rect 28140 28590 28142 28642
rect 28194 28590 28196 28642
rect 28140 28578 28196 28590
rect 28812 28644 28868 28654
rect 27916 28084 27972 28094
rect 27916 27858 27972 28028
rect 27916 27806 27918 27858
rect 27970 27806 27972 27858
rect 27916 27636 27972 27806
rect 28812 27858 28868 28588
rect 28812 27806 28814 27858
rect 28866 27806 28868 27858
rect 28812 27794 28868 27806
rect 28924 28420 28980 29036
rect 28924 27858 28980 28364
rect 29036 28196 29092 29260
rect 29372 28980 29428 28990
rect 29204 28532 29260 28542
rect 29036 28130 29092 28140
rect 29148 28530 29260 28532
rect 29148 28478 29206 28530
rect 29258 28478 29260 28530
rect 29148 28466 29260 28478
rect 28924 27806 28926 27858
rect 28978 27806 28980 27858
rect 28924 27794 28980 27806
rect 28532 27636 28588 27646
rect 27916 27570 27972 27580
rect 28476 27634 28588 27636
rect 28476 27582 28534 27634
rect 28586 27582 28588 27634
rect 28476 27570 28588 27582
rect 27804 27234 27860 27244
rect 26908 27022 26910 27074
rect 26962 27022 26964 27074
rect 26908 27010 26964 27022
rect 27020 27074 27076 27086
rect 27020 27022 27022 27074
rect 27074 27022 27076 27074
rect 27020 26964 27076 27022
rect 27356 27076 27412 27086
rect 27356 26982 27412 27020
rect 28084 27076 28140 27086
rect 28364 27076 28420 27086
rect 28084 26982 28140 27020
rect 28252 27074 28420 27076
rect 28252 27022 28366 27074
rect 28418 27022 28420 27074
rect 28252 27020 28420 27022
rect 27020 26898 27076 26908
rect 27188 26516 27244 26526
rect 27188 26514 28084 26516
rect 27188 26462 27190 26514
rect 27242 26462 28084 26514
rect 27188 26460 28084 26462
rect 27188 26450 27244 26460
rect 26908 26290 26964 26302
rect 26908 26238 26910 26290
rect 26962 26238 26964 26290
rect 26908 25396 26964 26238
rect 27020 26290 27076 26302
rect 27020 26238 27022 26290
rect 27074 26238 27076 26290
rect 27020 26180 27076 26238
rect 27020 26114 27076 26124
rect 27580 26290 27636 26302
rect 27580 26238 27582 26290
rect 27634 26238 27636 26290
rect 27580 25508 27636 26238
rect 27580 25442 27636 25452
rect 27804 26292 27860 26302
rect 27804 25478 27860 26236
rect 27804 25426 27806 25478
rect 27858 25426 27860 25478
rect 27804 25414 27860 25426
rect 27916 26180 27972 26190
rect 26908 25340 27076 25396
rect 26796 25106 26852 25116
rect 26684 24882 26740 24892
rect 25396 23378 25508 23390
rect 25396 23326 25398 23378
rect 25450 23326 25508 23378
rect 25396 23314 25508 23326
rect 25452 21924 25508 23314
rect 25452 21858 25508 21868
rect 25564 24444 26068 24500
rect 25228 20962 25284 20972
rect 25340 21362 25396 21374
rect 25340 21310 25342 21362
rect 25394 21310 25396 21362
rect 25340 20916 25396 21310
rect 25340 20850 25396 20860
rect 24220 20524 24612 20580
rect 24108 20300 24276 20356
rect 23492 20242 23604 20254
rect 23492 20190 23494 20242
rect 23546 20190 23604 20242
rect 23492 20188 23604 20190
rect 23492 19908 23548 20188
rect 24052 20132 24108 20142
rect 24052 20038 24108 20076
rect 23492 19842 23548 19852
rect 24220 19236 24276 20300
rect 24444 19796 24500 19806
rect 24444 19702 24500 19740
rect 24556 19460 24612 20524
rect 24780 20018 24836 20748
rect 24780 19966 24782 20018
rect 24834 19966 24836 20018
rect 24780 19954 24836 19966
rect 24892 20802 25172 20804
rect 24892 20750 25118 20802
rect 25170 20750 25172 20802
rect 24892 20748 25172 20750
rect 24892 20132 24948 20748
rect 25116 20738 25172 20748
rect 24052 19234 24276 19236
rect 24052 19182 24222 19234
rect 24274 19182 24276 19234
rect 24052 19180 24276 19182
rect 23884 19124 23940 19134
rect 23884 19030 23940 19068
rect 24052 18674 24108 19180
rect 24220 19170 24276 19180
rect 24444 19458 24612 19460
rect 24444 19406 24558 19458
rect 24610 19406 24612 19458
rect 24444 19404 24612 19406
rect 24052 18622 24054 18674
rect 24106 18622 24108 18674
rect 23436 18452 23492 18462
rect 23324 18396 23436 18452
rect 23324 18282 23380 18294
rect 23324 18230 23326 18282
rect 23378 18230 23380 18282
rect 23324 18004 23380 18230
rect 23100 17948 23380 18004
rect 23100 17668 23156 17948
rect 23436 17892 23492 18396
rect 23100 17574 23156 17612
rect 23324 17836 23492 17892
rect 24052 17892 24108 18622
rect 24220 18452 24276 18462
rect 24220 18358 24276 18396
rect 23324 17666 23380 17836
rect 24052 17826 24108 17836
rect 23324 17614 23326 17666
rect 23378 17614 23380 17666
rect 23772 17668 23828 17678
rect 23324 17602 23380 17614
rect 23492 17610 23548 17622
rect 23492 17558 23494 17610
rect 23546 17558 23548 17610
rect 23772 17574 23828 17612
rect 24332 17668 24388 17678
rect 22764 17444 22820 17454
rect 22764 17442 23268 17444
rect 22764 17390 22766 17442
rect 22818 17390 23268 17442
rect 22764 17388 23268 17390
rect 22764 17378 22820 17388
rect 23100 17108 23156 17118
rect 22764 16882 22820 16894
rect 22764 16830 22766 16882
rect 22818 16830 22820 16882
rect 22764 16772 22820 16830
rect 23100 16882 23156 17052
rect 23100 16830 23102 16882
rect 23154 16830 23156 16882
rect 23100 16818 23156 16830
rect 22764 15428 22820 16716
rect 22988 16100 23044 16110
rect 23212 16100 23268 17388
rect 23492 17332 23548 17558
rect 23660 17556 23716 17566
rect 23660 17462 23716 17500
rect 24052 17556 24108 17566
rect 24052 17554 24276 17556
rect 24052 17502 24054 17554
rect 24106 17502 24276 17554
rect 24052 17500 24276 17502
rect 24052 17490 24108 17500
rect 23324 17276 23548 17332
rect 23660 17332 23716 17342
rect 23324 16772 23380 17276
rect 23548 17108 23604 17118
rect 23436 16996 23492 17006
rect 23436 16902 23492 16940
rect 23324 16706 23380 16716
rect 22988 15540 23044 16044
rect 22988 15474 23044 15484
rect 23100 16098 23268 16100
rect 23100 16046 23214 16098
rect 23266 16046 23268 16098
rect 23100 16044 23268 16046
rect 22764 15362 22820 15372
rect 23100 15148 23156 16044
rect 23212 16034 23268 16044
rect 23324 16266 23380 16278
rect 23324 16214 23326 16266
rect 23378 16214 23380 16266
rect 23324 16100 23380 16214
rect 23324 16034 23380 16044
rect 23548 16098 23604 17052
rect 23548 16046 23550 16098
rect 23602 16046 23604 16098
rect 23548 16034 23604 16046
rect 23660 15876 23716 17276
rect 24108 17108 24164 17118
rect 24108 16938 24164 17052
rect 24108 16886 24110 16938
rect 24162 16886 24164 16938
rect 24108 16874 24164 16886
rect 24220 16324 24276 17500
rect 24332 16882 24388 17612
rect 24444 17108 24500 19404
rect 24556 19394 24612 19404
rect 24892 19236 24948 20076
rect 25228 20045 25284 20058
rect 25228 20020 25230 20045
rect 25282 20020 25284 20045
rect 25564 20020 25620 24444
rect 27020 24388 27076 25340
rect 27244 25172 27300 25182
rect 26852 24332 27076 24388
rect 27132 24612 27188 24622
rect 25900 24276 25956 24286
rect 25732 24052 25788 24062
rect 25900 24052 25956 24220
rect 25788 23996 25956 24052
rect 25732 23958 25788 23996
rect 25900 23940 25956 23996
rect 26684 24164 26740 24174
rect 26572 23940 26628 23950
rect 25900 23922 26012 23940
rect 25900 23884 25958 23922
rect 25956 23870 25958 23884
rect 26010 23870 26012 23922
rect 25956 23858 26012 23870
rect 26124 23882 26180 23894
rect 26124 23830 26126 23882
rect 26178 23830 26180 23882
rect 26012 23182 26068 23194
rect 25732 23156 25788 23166
rect 25732 23062 25788 23100
rect 26012 23156 26014 23182
rect 26066 23156 26068 23182
rect 25900 22484 25956 22494
rect 26012 22484 26068 23100
rect 26124 23044 26180 23830
rect 26348 23882 26404 23894
rect 26348 23830 26350 23882
rect 26402 23830 26404 23882
rect 26572 23858 26574 23884
rect 26626 23858 26628 23884
rect 26572 23846 26628 23858
rect 26348 23548 26404 23830
rect 26236 23492 26404 23548
rect 26236 23210 26292 23492
rect 26348 23426 26404 23436
rect 26236 23158 26238 23210
rect 26290 23158 26292 23210
rect 26460 23268 26516 23278
rect 26684 23268 26740 24108
rect 26852 24162 26908 24332
rect 26852 24110 26854 24162
rect 26906 24110 26908 24162
rect 26852 24098 26908 24110
rect 27132 23938 27188 24556
rect 27244 24164 27300 25116
rect 27804 24612 27860 24622
rect 27244 24098 27300 24108
rect 27356 24610 27860 24612
rect 27356 24558 27806 24610
rect 27858 24558 27860 24610
rect 27356 24556 27860 24558
rect 27132 23886 27134 23938
rect 27186 23886 27188 23938
rect 27132 23874 27188 23886
rect 27356 23940 27412 24556
rect 27804 24546 27860 24556
rect 27356 23846 27412 23884
rect 27636 23828 27692 23838
rect 26460 23201 26516 23212
rect 26404 23189 26516 23201
rect 26404 23184 26406 23189
rect 26236 23146 26292 23158
rect 26348 23137 26406 23184
rect 26458 23137 26516 23189
rect 26647 23210 26740 23268
rect 26647 23158 26649 23210
rect 26701 23158 26740 23210
rect 27468 23826 27692 23828
rect 27468 23774 27638 23826
rect 27690 23774 27692 23826
rect 27468 23772 27692 23774
rect 26647 23146 26740 23158
rect 26348 23128 26516 23137
rect 26348 23125 26460 23128
rect 26348 23044 26404 23125
rect 26124 22988 26404 23044
rect 26684 22820 26740 23146
rect 26796 23154 26852 23166
rect 26796 23102 26798 23154
rect 26850 23102 26852 23154
rect 26796 23044 26852 23102
rect 27020 23156 27076 23166
rect 27468 23156 27524 23772
rect 27636 23762 27692 23772
rect 27020 23062 27076 23100
rect 27132 23100 27524 23156
rect 27804 23154 27860 23166
rect 27804 23102 27806 23154
rect 27858 23102 27860 23154
rect 26796 22978 26852 22988
rect 26684 22764 26908 22820
rect 25900 22482 26068 22484
rect 25900 22430 25902 22482
rect 25954 22430 26068 22482
rect 25900 22428 26068 22430
rect 26852 22482 26908 22764
rect 26852 22430 26854 22482
rect 26906 22430 26908 22482
rect 25900 22418 25956 22428
rect 26852 22418 26908 22430
rect 26572 22260 26628 22270
rect 25676 21588 25732 21598
rect 25676 21494 25732 21532
rect 26572 21586 26628 22204
rect 26572 21534 26574 21586
rect 26626 21534 26628 21586
rect 26572 21522 26628 21534
rect 26964 21588 27020 21598
rect 26964 21494 27020 21532
rect 26236 21364 26292 21374
rect 25900 21362 26292 21364
rect 25900 21310 26238 21362
rect 26290 21310 26292 21362
rect 25900 21308 26292 21310
rect 25900 20914 25956 21308
rect 26236 21298 26292 21308
rect 25900 20862 25902 20914
rect 25954 20862 25956 20914
rect 25900 20850 25956 20862
rect 25228 19954 25284 19964
rect 25340 19964 25620 20020
rect 24892 19142 24948 19180
rect 24556 18340 24612 18350
rect 24556 18246 24612 18284
rect 24892 18340 24948 18350
rect 24780 17666 24836 17678
rect 24780 17614 24782 17666
rect 24834 17614 24836 17666
rect 24780 17556 24836 17614
rect 24780 17490 24836 17500
rect 24612 17442 24668 17454
rect 24612 17390 24614 17442
rect 24666 17390 24668 17442
rect 24612 17332 24668 17390
rect 24612 17266 24668 17276
rect 24444 17052 24780 17108
rect 24332 16830 24334 16882
rect 24386 16830 24388 16882
rect 24724 16938 24780 17052
rect 24724 16886 24726 16938
rect 24778 16886 24780 16938
rect 24724 16874 24780 16886
rect 24332 16818 24388 16830
rect 24220 16258 24276 16268
rect 24556 16770 24612 16782
rect 24556 16718 24558 16770
rect 24610 16718 24612 16770
rect 24220 16100 24276 16110
rect 23548 15820 23716 15876
rect 23884 15874 23940 15886
rect 23884 15822 23886 15874
rect 23938 15822 23940 15874
rect 23212 15316 23268 15326
rect 23212 15222 23268 15260
rect 22988 15092 23156 15148
rect 22652 13122 22708 13132
rect 22876 13779 22932 13791
rect 22876 13727 22878 13779
rect 22930 13727 22932 13779
rect 22428 12910 22430 12962
rect 22482 12910 22484 12962
rect 22428 12898 22484 12910
rect 22764 12962 22820 12974
rect 22764 12910 22766 12962
rect 22818 12910 22820 12962
rect 22092 12740 22148 12750
rect 22764 12740 22820 12910
rect 22092 12738 22820 12740
rect 22092 12686 22094 12738
rect 22146 12686 22820 12738
rect 22092 12684 22820 12686
rect 22092 12674 22148 12684
rect 21924 12404 21980 12414
rect 21924 12290 21980 12348
rect 21924 12238 21926 12290
rect 21978 12238 21980 12290
rect 21924 12226 21980 12238
rect 19740 11676 20244 11732
rect 20412 12122 20468 12134
rect 20412 12070 20414 12122
rect 20466 12070 20468 12122
rect 21308 12126 21310 12178
rect 21362 12126 21364 12178
rect 21308 12114 21364 12126
rect 21420 12178 21476 12190
rect 21420 12126 21422 12178
rect 21474 12126 21476 12178
rect 20412 11732 20468 12070
rect 19740 11620 19796 11676
rect 20412 11666 20468 11676
rect 20972 11954 21028 11966
rect 20972 11902 20974 11954
rect 21026 11902 21028 11954
rect 19740 11526 19796 11564
rect 20748 11620 20804 11630
rect 20076 11396 20132 11406
rect 19628 11394 20132 11396
rect 19628 11342 20078 11394
rect 20130 11342 20132 11394
rect 19628 11340 20132 11342
rect 20076 11330 20132 11340
rect 20412 11396 20468 11406
rect 20412 11302 20468 11340
rect 20748 11394 20804 11564
rect 20748 11342 20750 11394
rect 20802 11342 20804 11394
rect 20748 11330 20804 11342
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 20338 10836 20394 10846
rect 20338 10648 20394 10780
rect 20338 10596 20340 10648
rect 20392 10596 20394 10648
rect 20338 10584 20394 10596
rect 20524 10724 20580 10734
rect 20524 10610 20580 10668
rect 20972 10724 21028 11902
rect 21420 11844 21476 12126
rect 21420 11778 21476 11788
rect 21644 12178 21700 12190
rect 21644 12126 21646 12178
rect 21698 12126 21700 12178
rect 21644 11630 21700 12126
rect 22764 12180 22820 12684
rect 22876 12404 22932 13727
rect 22988 13524 23044 15092
rect 23212 14420 23268 14430
rect 22988 13458 23044 13468
rect 23100 14084 23156 14094
rect 23100 13186 23156 14028
rect 23212 13802 23268 14364
rect 23212 13750 23214 13802
rect 23266 13750 23268 13802
rect 23212 13738 23268 13750
rect 23436 14308 23492 14318
rect 23100 13134 23102 13186
rect 23154 13134 23156 13186
rect 23100 13122 23156 13134
rect 23212 13412 23268 13422
rect 22876 12338 22932 12348
rect 22932 12234 22988 12246
rect 22932 12182 22934 12234
rect 22986 12182 22988 12234
rect 22932 12180 22988 12182
rect 23100 12180 23156 12190
rect 23212 12180 23268 13356
rect 23436 12962 23492 14252
rect 23548 13636 23604 15820
rect 23884 15652 23940 15822
rect 23884 15586 23940 15596
rect 23772 15482 23828 15494
rect 23772 15430 23774 15482
rect 23826 15430 23828 15482
rect 23660 15353 23716 15365
rect 23660 15301 23662 15353
rect 23714 15301 23716 15353
rect 23660 15204 23716 15301
rect 23660 15138 23716 15148
rect 23772 13802 23828 15430
rect 23884 15316 23940 15326
rect 23884 15222 23940 15260
rect 24220 14308 24276 16044
rect 24444 16100 24500 16110
rect 24556 16100 24612 16718
rect 24444 16098 24612 16100
rect 24444 16046 24446 16098
rect 24498 16046 24612 16098
rect 24444 16044 24612 16046
rect 24444 16034 24500 16044
rect 24724 15988 24780 15998
rect 24724 15894 24780 15932
rect 24892 15764 24948 18284
rect 25228 17780 25284 17790
rect 25228 17638 25284 17724
rect 25228 17586 25230 17638
rect 25282 17586 25284 17638
rect 25228 17574 25284 17586
rect 25340 17444 25396 19964
rect 25564 19796 25620 19806
rect 25340 17378 25396 17388
rect 25452 17668 25508 17678
rect 25452 16334 25508 17612
rect 25564 17220 25620 19740
rect 25676 19236 25732 19246
rect 25676 19234 25956 19236
rect 25676 19182 25678 19234
rect 25730 19182 25956 19234
rect 25676 19180 25956 19182
rect 25676 19170 25732 19180
rect 25900 18676 25956 19180
rect 26012 18676 26068 18686
rect 25900 18674 26068 18676
rect 25900 18622 26014 18674
rect 26066 18622 26068 18674
rect 25900 18620 26068 18622
rect 26012 18610 26068 18620
rect 26348 18564 26404 18574
rect 26348 18450 26404 18508
rect 26348 18398 26350 18450
rect 26402 18398 26404 18450
rect 26348 18386 26404 18398
rect 27132 18452 27188 23100
rect 27300 22932 27356 22942
rect 27804 22932 27860 23102
rect 27300 22930 27524 22932
rect 27300 22878 27302 22930
rect 27354 22878 27524 22930
rect 27300 22876 27524 22878
rect 27300 22866 27356 22876
rect 27468 21812 27524 22876
rect 27804 22484 27860 22876
rect 27916 22596 27972 26124
rect 28028 25506 28084 26460
rect 28252 25618 28308 27020
rect 28364 27010 28420 27020
rect 28364 26852 28420 26862
rect 28364 26290 28420 26796
rect 28364 26238 28366 26290
rect 28418 26238 28420 26290
rect 28364 26226 28420 26238
rect 28252 25566 28254 25618
rect 28306 25566 28308 25618
rect 28252 25554 28308 25566
rect 28476 25620 28532 27570
rect 28588 27188 28644 27198
rect 28588 27074 28644 27132
rect 28588 27022 28590 27074
rect 28642 27022 28644 27074
rect 28588 27010 28644 27022
rect 29036 27076 29092 27086
rect 29036 26982 29092 27020
rect 29148 26908 29204 28466
rect 29372 28420 29428 28924
rect 29708 28868 29764 28878
rect 29484 28644 29540 28654
rect 29484 28550 29540 28588
rect 29708 28642 29764 28812
rect 29708 28590 29710 28642
rect 29762 28590 29764 28642
rect 29708 28578 29764 28590
rect 29372 28364 29540 28420
rect 29372 28196 29428 28206
rect 29372 28082 29428 28140
rect 29372 28030 29374 28082
rect 29426 28030 29428 28082
rect 29372 28018 29428 28030
rect 28588 26852 29204 26908
rect 29372 26964 29428 27002
rect 29372 26898 29428 26908
rect 28588 25844 28644 26852
rect 28588 25788 28868 25844
rect 28476 25564 28644 25620
rect 28028 25454 28030 25506
rect 28082 25454 28084 25506
rect 28028 25442 28084 25454
rect 28420 25450 28476 25462
rect 28420 25398 28422 25450
rect 28474 25398 28476 25450
rect 28420 24836 28476 25398
rect 28140 24780 28476 24836
rect 28140 24052 28196 24780
rect 28588 24724 28644 25564
rect 28140 23938 28196 23996
rect 28364 24668 28644 24724
rect 28140 23886 28142 23938
rect 28194 23886 28196 23938
rect 28140 23874 28196 23886
rect 28252 23940 28308 23950
rect 28252 23846 28308 23884
rect 28140 23492 28196 23502
rect 28140 23198 28196 23436
rect 28140 23146 28142 23198
rect 28194 23146 28196 23198
rect 28140 23134 28196 23146
rect 28252 23044 28308 23054
rect 27916 22530 27972 22540
rect 28140 23042 28308 23044
rect 28140 22990 28254 23042
rect 28306 22990 28308 23042
rect 28140 22988 28308 22990
rect 27804 22418 27860 22428
rect 27916 22372 27972 22382
rect 27916 22290 27918 22316
rect 27970 22290 27972 22316
rect 27636 22260 27692 22270
rect 27636 22166 27692 22204
rect 27468 21746 27524 21756
rect 27804 21588 27860 21598
rect 27468 21586 27860 21588
rect 27468 21534 27806 21586
rect 27858 21534 27860 21586
rect 27468 21532 27860 21534
rect 27468 20132 27524 21532
rect 27804 21522 27860 21532
rect 27804 20916 27860 20926
rect 27916 20916 27972 22290
rect 28140 22314 28196 22988
rect 28252 22978 28308 22988
rect 28364 22484 28420 24668
rect 28532 24500 28588 24510
rect 28532 24162 28588 24444
rect 28532 24110 28534 24162
rect 28586 24110 28588 24162
rect 28532 24098 28588 24110
rect 28812 23604 28868 25788
rect 29036 25508 29092 25518
rect 28588 23548 28868 23604
rect 28924 25396 28980 25406
rect 28588 23492 28644 23548
rect 28140 22262 28142 22314
rect 28194 22262 28196 22314
rect 28140 21812 28196 22262
rect 28140 21746 28196 21756
rect 28252 22428 28420 22484
rect 28476 22596 28532 22606
rect 27804 20914 27972 20916
rect 27804 20862 27806 20914
rect 27858 20862 27972 20914
rect 27804 20860 27972 20862
rect 27804 20850 27860 20860
rect 27468 20018 27524 20076
rect 27468 19966 27470 20018
rect 27522 19966 27524 20018
rect 27468 19954 27524 19966
rect 28252 20132 28308 22428
rect 28476 22335 28532 22540
rect 28364 22314 28420 22326
rect 28364 22262 28366 22314
rect 28418 22262 28420 22314
rect 28476 22283 28478 22335
rect 28530 22283 28532 22335
rect 28476 22271 28532 22283
rect 28364 22148 28420 22262
rect 28588 22148 28644 23436
rect 28700 23156 28756 23166
rect 28700 23062 28756 23100
rect 28364 22092 28588 22148
rect 28588 22054 28644 22092
rect 28924 21812 28980 25340
rect 29036 24946 29092 25452
rect 29484 25172 29540 28364
rect 30044 28196 30100 28206
rect 30044 28082 30100 28140
rect 30044 28030 30046 28082
rect 30098 28030 30100 28082
rect 30044 28018 30100 28030
rect 29708 27858 29764 27870
rect 29708 27806 29710 27858
rect 29762 27806 29764 27858
rect 29708 27300 29764 27806
rect 29708 27234 29764 27244
rect 29484 25106 29540 25116
rect 29708 27074 29764 27086
rect 29708 27022 29710 27074
rect 29762 27022 29764 27074
rect 29036 24894 29038 24946
rect 29090 24894 29092 24946
rect 29036 23938 29092 24894
rect 29708 24500 29764 27022
rect 30044 26852 30100 26862
rect 29820 26850 30100 26852
rect 29820 26798 30046 26850
rect 30098 26798 30100 26850
rect 29820 26796 30100 26798
rect 29820 25618 29876 26796
rect 30044 26786 30100 26796
rect 30156 25844 30212 30828
rect 30324 29092 30380 29102
rect 30324 28866 30380 29036
rect 30324 28814 30326 28866
rect 30378 28814 30380 28866
rect 30324 28802 30380 28814
rect 30380 27972 30436 27982
rect 30380 27858 30436 27916
rect 30380 27806 30382 27858
rect 30434 27806 30436 27858
rect 30268 26404 30324 26414
rect 30380 26404 30436 27806
rect 30492 26908 30548 30940
rect 30716 30930 30772 30940
rect 31108 30930 31164 30940
rect 31724 30210 31780 30222
rect 31724 30158 31726 30210
rect 31778 30158 31780 30210
rect 31724 29988 31780 30158
rect 30604 29876 30660 29886
rect 30604 28642 30660 29820
rect 31724 29652 31780 29932
rect 31836 30210 31892 30222
rect 31836 30158 31838 30210
rect 31890 30158 31892 30210
rect 31836 29876 31892 30158
rect 31836 29810 31892 29820
rect 31948 29764 32004 32060
rect 32172 31892 32228 31902
rect 32060 31836 32172 31892
rect 32060 31050 32116 31836
rect 32172 31798 32228 31836
rect 32284 31734 32340 31746
rect 32284 31682 32286 31734
rect 32338 31682 32340 31734
rect 32284 31220 32340 31682
rect 32396 31444 32452 32284
rect 32956 32004 33012 33292
rect 33068 33282 33124 33292
rect 33124 32788 33180 32798
rect 33124 32674 33180 32732
rect 33124 32622 33126 32674
rect 33178 32622 33180 32674
rect 33124 32610 33180 32622
rect 33292 32676 33348 33516
rect 33628 32788 33684 32798
rect 33516 32732 33628 32788
rect 33292 32620 33404 32676
rect 33348 32618 33404 32620
rect 33348 32566 33350 32618
rect 33402 32566 33404 32618
rect 33348 32554 33404 32566
rect 33068 32004 33124 32014
rect 32956 31948 33068 32004
rect 32396 31378 32452 31388
rect 32620 31778 32676 31790
rect 32620 31726 32622 31778
rect 32674 31726 32676 31778
rect 32060 30998 32062 31050
rect 32114 30998 32116 31050
rect 32060 30986 32116 30998
rect 32172 31164 32340 31220
rect 32396 31220 32452 31230
rect 32172 30446 32228 31164
rect 32396 31050 32452 31164
rect 32284 31022 32340 31034
rect 32284 30996 32286 31022
rect 32338 30996 32340 31022
rect 32396 30998 32398 31050
rect 32450 30998 32452 31050
rect 32396 30986 32452 30998
rect 32508 30996 32564 31006
rect 32284 30930 32340 30940
rect 32116 30436 32228 30446
rect 32508 30436 32564 30940
rect 32620 30884 32676 31726
rect 33068 31778 33124 31948
rect 33068 31726 33070 31778
rect 33122 31726 33124 31778
rect 33068 31714 33124 31726
rect 33404 31444 33460 31454
rect 33236 30884 33292 30894
rect 32620 30882 33292 30884
rect 32620 30830 33238 30882
rect 33290 30830 33292 30882
rect 32620 30828 33292 30830
rect 33180 30818 33292 30828
rect 32732 30436 32788 30446
rect 32116 30434 32452 30436
rect 32116 30382 32118 30434
rect 32170 30382 32452 30434
rect 32116 30380 32452 30382
rect 32508 30434 32788 30436
rect 32508 30382 32734 30434
rect 32786 30382 32788 30434
rect 32508 30380 32788 30382
rect 32116 30370 32172 30380
rect 32396 30210 32452 30380
rect 32732 30370 32788 30380
rect 33068 30212 33124 30222
rect 32396 30158 32398 30210
rect 32450 30158 32452 30210
rect 32396 30146 32452 30158
rect 32620 30210 33124 30212
rect 32620 30158 33070 30210
rect 33122 30158 33124 30210
rect 32620 30156 33124 30158
rect 31948 29698 32004 29708
rect 31724 29596 31892 29652
rect 31276 29426 31332 29438
rect 31276 29374 31278 29426
rect 31330 29374 31332 29426
rect 30828 29316 30884 29326
rect 31276 29316 31332 29374
rect 30828 29314 31332 29316
rect 30828 29262 30830 29314
rect 30882 29262 31332 29314
rect 30828 29260 31332 29262
rect 30828 29250 30884 29260
rect 30940 28756 30996 28766
rect 30604 28590 30606 28642
rect 30658 28590 30660 28642
rect 30604 28578 30660 28590
rect 30828 28642 30884 28654
rect 30828 28590 30830 28642
rect 30882 28590 30884 28642
rect 30828 27748 30884 28590
rect 30940 28420 30996 28700
rect 31052 28644 31108 28654
rect 31052 28642 31220 28644
rect 31052 28590 31054 28642
rect 31106 28590 31220 28642
rect 31052 28588 31220 28590
rect 31052 28578 31108 28588
rect 30940 28364 31108 28420
rect 31052 28026 31108 28364
rect 31052 27974 31054 28026
rect 31106 27974 31108 28026
rect 31052 27962 31108 27974
rect 31164 28196 31220 28588
rect 31164 27858 31220 28140
rect 31164 27806 31166 27858
rect 31218 27806 31220 27858
rect 31164 27794 31220 27806
rect 31276 27860 31332 29260
rect 31388 29426 31444 29438
rect 31388 29374 31390 29426
rect 31442 29374 31444 29426
rect 31388 27972 31444 29374
rect 31668 29204 31724 29214
rect 31388 27906 31444 27916
rect 31612 29202 31724 29204
rect 31612 29150 31670 29202
rect 31722 29150 31724 29202
rect 31612 29138 31724 29150
rect 31276 27794 31332 27804
rect 30828 27682 30884 27692
rect 31612 27748 31668 29138
rect 31836 28868 31892 29596
rect 31836 28810 31892 28812
rect 31836 28758 31838 28810
rect 31890 28758 31892 28810
rect 31836 28746 31892 28758
rect 32620 28754 32676 30156
rect 33068 30146 33124 30156
rect 32620 28702 32622 28754
rect 32674 28702 32676 28754
rect 31724 28644 31780 28654
rect 32172 28644 32228 28654
rect 31724 28642 32452 28644
rect 31724 28590 31726 28642
rect 31778 28590 32174 28642
rect 32226 28590 32452 28642
rect 31724 28588 32452 28590
rect 31724 28578 31780 28588
rect 31836 27860 31892 28588
rect 32172 28578 32228 28588
rect 32396 28082 32452 28588
rect 32396 28030 32398 28082
rect 32450 28030 32452 28082
rect 32396 28018 32452 28030
rect 32508 28598 32564 28610
rect 32508 28546 32510 28598
rect 32562 28546 32564 28598
rect 32508 28196 32564 28546
rect 32620 28420 32676 28702
rect 32732 29764 32788 29774
rect 33180 29764 33236 30818
rect 33404 30324 33460 31388
rect 33516 30996 33572 32732
rect 33628 32722 33684 32732
rect 33628 32590 33684 32602
rect 33628 32564 33630 32590
rect 33682 32564 33684 32590
rect 33628 32498 33684 32508
rect 33740 31220 33796 33964
rect 33852 33908 33908 34078
rect 33990 34020 34046 34188
rect 33852 33842 33908 33852
rect 33964 33964 34046 34020
rect 34412 34020 34468 35308
rect 34916 35364 34972 35374
rect 34916 34914 34972 35308
rect 34916 34862 34918 34914
rect 34970 34862 34972 34914
rect 34916 34850 34972 34862
rect 34972 34356 35028 34366
rect 33852 33460 33908 33470
rect 33964 33460 34020 33964
rect 34412 33954 34468 33964
rect 34524 34354 35028 34356
rect 34524 34302 34974 34354
rect 35026 34302 35028 34354
rect 34524 34300 35028 34302
rect 34132 33908 34188 33918
rect 34132 33814 34188 33852
rect 34524 33684 34580 34300
rect 34972 34290 35028 34300
rect 33852 33458 34020 33460
rect 33852 33406 33854 33458
rect 33906 33406 34020 33458
rect 33852 33404 34020 33406
rect 34076 33628 34580 33684
rect 34636 34130 34692 34142
rect 34636 34078 34638 34130
rect 34690 34078 34692 34130
rect 34636 33684 34692 34078
rect 34636 33628 35028 33684
rect 33852 33394 33908 33404
rect 33964 33124 34020 33134
rect 33852 32788 33908 32798
rect 33852 32618 33908 32732
rect 33852 32566 33854 32618
rect 33906 32566 33908 32618
rect 33852 32554 33908 32566
rect 33964 32618 34020 33068
rect 33964 32566 33966 32618
rect 34018 32566 34020 32618
rect 33964 32554 34020 32566
rect 34076 32452 34132 33628
rect 34860 32900 34916 32910
rect 34412 32788 34468 32798
rect 34412 32618 34468 32732
rect 34300 32597 34356 32609
rect 33852 32396 34132 32452
rect 34188 32564 34244 32574
rect 33852 31890 33908 32396
rect 34188 32116 34244 32508
rect 33852 31838 33854 31890
rect 33906 31838 33908 31890
rect 33852 31826 33908 31838
rect 34076 32060 34244 32116
rect 34300 32545 34302 32597
rect 34354 32545 34356 32597
rect 34412 32566 34414 32618
rect 34466 32566 34468 32618
rect 34860 32618 34916 32844
rect 34412 32554 34468 32566
rect 34636 32590 34692 32602
rect 34636 32564 34638 32590
rect 34690 32564 34692 32590
rect 34300 32340 34356 32545
rect 34860 32566 34862 32618
rect 34914 32566 34916 32618
rect 34860 32554 34916 32566
rect 34636 32498 34692 32508
rect 34300 32116 34356 32284
rect 34076 31892 34132 32060
rect 34300 32050 34356 32060
rect 33740 31164 33908 31220
rect 33628 31108 33684 31118
rect 33628 31050 33684 31052
rect 33628 30998 33630 31050
rect 33682 30998 33684 31050
rect 33628 30986 33684 30998
rect 33740 31022 33796 31034
rect 33516 30884 33572 30940
rect 33740 30970 33742 31022
rect 33794 30970 33796 31022
rect 33740 30884 33796 30970
rect 33516 30828 33796 30884
rect 33852 30548 33908 31164
rect 34076 31062 34132 31836
rect 34972 31556 35028 33628
rect 35084 32686 35140 35644
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35644 35196 36148 35252
rect 35644 35082 35700 35196
rect 35532 35028 35588 35038
rect 35644 35030 35646 35082
rect 35698 35030 35700 35082
rect 35644 35018 35700 35030
rect 35980 35026 36036 35038
rect 35196 34914 35252 34926
rect 35196 34862 35198 34914
rect 35250 34862 35252 34914
rect 35196 33908 35252 34862
rect 35532 34914 35588 34972
rect 35532 34862 35534 34914
rect 35586 34862 35588 34914
rect 35532 34850 35588 34862
rect 35980 34974 35982 35026
rect 36034 34974 36036 35026
rect 35308 34130 35364 34142
rect 35308 34078 35310 34130
rect 35362 34078 35364 34130
rect 35308 33908 35364 34078
rect 35980 34132 36036 34974
rect 36092 34899 36148 35196
rect 36092 34847 36094 34899
rect 36146 34847 36148 34899
rect 36092 34835 36148 34847
rect 36092 34132 36148 34142
rect 35980 34130 36148 34132
rect 35980 34078 36094 34130
rect 36146 34078 36148 34130
rect 35980 34076 36148 34078
rect 36092 34066 36148 34076
rect 35644 34020 35700 34030
rect 35308 33852 35588 33908
rect 35196 33842 35252 33852
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35532 32788 35588 33852
rect 35644 33236 35700 33964
rect 35644 33170 35700 33180
rect 35756 33572 35812 33582
rect 35756 33458 35812 33516
rect 35756 33406 35758 33458
rect 35810 33406 35812 33458
rect 35756 32900 35812 33406
rect 35756 32834 35812 32844
rect 35084 32674 35196 32686
rect 35084 32622 35142 32674
rect 35194 32622 35196 32674
rect 35084 32620 35196 32622
rect 35140 32610 35196 32620
rect 35532 32562 35588 32732
rect 35532 32510 35534 32562
rect 35586 32510 35588 32562
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 34468 31500 35028 31556
rect 35532 32004 35588 32510
rect 34020 31050 34132 31062
rect 34020 30998 34022 31050
rect 34074 30998 34132 31050
rect 34020 30996 34132 30998
rect 34188 31444 34244 31454
rect 34188 31050 34244 31388
rect 34188 30998 34190 31050
rect 34242 30998 34244 31050
rect 34468 31106 34524 31500
rect 34468 31054 34470 31106
rect 34522 31054 34524 31106
rect 34468 31042 34524 31054
rect 34748 31108 34804 31118
rect 34020 30986 34076 30996
rect 34188 30986 34244 30998
rect 33404 30258 33460 30268
rect 33628 30492 33908 30548
rect 33628 30222 33684 30492
rect 33292 30212 33348 30222
rect 33292 30118 33348 30156
rect 33572 30210 33684 30222
rect 33572 30158 33574 30210
rect 33626 30158 33684 30210
rect 33572 30156 33684 30158
rect 33964 30210 34020 30222
rect 33964 30158 33966 30210
rect 34018 30158 34020 30210
rect 34636 30210 34692 30222
rect 33572 30146 33628 30156
rect 32732 28420 32788 29708
rect 32956 29708 33236 29764
rect 32844 28756 32900 28766
rect 32844 28642 32900 28700
rect 32844 28590 32846 28642
rect 32898 28590 32900 28642
rect 32844 28578 32900 28590
rect 32732 28364 32900 28420
rect 32620 28354 32676 28364
rect 32508 27972 32564 28140
rect 32508 27916 32788 27972
rect 32060 27860 32116 27870
rect 31836 27858 32004 27860
rect 31836 27806 31838 27858
rect 31890 27806 32004 27858
rect 31836 27804 32004 27806
rect 31836 27794 31892 27804
rect 31612 27682 31668 27692
rect 30772 27300 30828 27310
rect 30772 27206 30828 27244
rect 31052 27074 31108 27086
rect 31052 27022 31054 27074
rect 31106 27022 31108 27074
rect 30492 26852 30660 26908
rect 30268 26402 30436 26404
rect 30268 26350 30270 26402
rect 30322 26350 30436 26402
rect 30268 26348 30436 26350
rect 30268 26338 30324 26348
rect 29820 25566 29822 25618
rect 29874 25566 29876 25618
rect 29820 25554 29876 25566
rect 30044 25788 30212 25844
rect 30604 25844 30660 26852
rect 31052 26404 31108 27022
rect 31276 27076 31332 27086
rect 31556 27076 31612 27086
rect 31276 27074 31612 27076
rect 31276 27022 31278 27074
rect 31330 27022 31558 27074
rect 31610 27022 31612 27074
rect 31276 27020 31612 27022
rect 31276 27010 31332 27020
rect 31556 27010 31612 27020
rect 31836 27076 31892 27086
rect 31836 26982 31892 27020
rect 31948 27074 32004 27804
rect 32060 27766 32116 27804
rect 32340 27188 32396 27198
rect 32340 27094 32396 27132
rect 31948 27022 31950 27074
rect 32002 27022 32004 27074
rect 31948 27010 32004 27022
rect 32620 27076 32676 27086
rect 32620 26982 32676 27020
rect 32732 27074 32788 27916
rect 32732 27022 32734 27074
rect 32786 27022 32788 27074
rect 32732 27010 32788 27022
rect 31052 26338 31108 26348
rect 31388 26628 31444 26638
rect 31388 26290 31444 26572
rect 32284 26404 32340 26414
rect 31388 26238 31390 26290
rect 31442 26238 31444 26290
rect 31724 26328 31780 26340
rect 31724 26292 31726 26328
rect 31778 26292 31780 26328
rect 32284 26310 32340 26348
rect 31388 26226 31444 26238
rect 31612 26234 31668 26246
rect 30884 26180 30940 26190
rect 31612 26182 31614 26234
rect 31666 26182 31668 26234
rect 31724 26226 31780 26236
rect 32452 26234 32508 26246
rect 30884 26178 30996 26180
rect 30884 26126 30886 26178
rect 30938 26126 30996 26178
rect 30884 26114 30996 26126
rect 30044 25396 30100 25788
rect 30604 25778 30660 25788
rect 30044 25330 30100 25340
rect 30940 25396 30996 26114
rect 31220 26068 31276 26078
rect 31612 26068 31668 26182
rect 31220 26066 31668 26068
rect 31220 26014 31222 26066
rect 31274 26014 31668 26066
rect 31220 26012 31668 26014
rect 32452 26182 32454 26234
rect 32506 26182 32508 26234
rect 31220 26002 31276 26012
rect 30940 25330 30996 25340
rect 31164 25844 31220 25854
rect 30716 25284 30772 25294
rect 30044 25172 30100 25182
rect 29708 24434 29764 24444
rect 29932 24948 29988 24958
rect 29820 23940 29876 23950
rect 29036 23886 29038 23938
rect 29090 23886 29092 23938
rect 29036 23874 29092 23886
rect 29708 23938 29876 23940
rect 29708 23886 29822 23938
rect 29874 23886 29876 23938
rect 29708 23884 29876 23886
rect 29596 23492 29652 23502
rect 29596 23210 29652 23436
rect 29036 23156 29092 23166
rect 29316 23156 29372 23166
rect 29036 23154 29372 23156
rect 29036 23102 29038 23154
rect 29090 23102 29318 23154
rect 29370 23102 29372 23154
rect 29596 23158 29598 23210
rect 29650 23158 29652 23210
rect 29596 23146 29652 23158
rect 29708 23156 29764 23884
rect 29820 23874 29876 23884
rect 29036 23100 29372 23102
rect 29036 23090 29092 23100
rect 29316 23090 29372 23100
rect 29820 23380 29876 23390
rect 29820 23210 29876 23324
rect 29820 23158 29822 23210
rect 29874 23158 29876 23210
rect 29820 23146 29876 23158
rect 29708 23090 29764 23100
rect 29316 22484 29372 22494
rect 29316 22390 29372 22428
rect 29932 22484 29988 24892
rect 30044 23716 30100 25116
rect 30716 24749 30772 25228
rect 31052 25284 31108 25294
rect 30716 24697 30718 24749
rect 30770 24697 30772 24749
rect 30716 24685 30772 24697
rect 30940 24836 30996 24846
rect 30940 23716 30996 24780
rect 30044 23660 30212 23716
rect 30044 23268 30100 23278
rect 30044 23210 30100 23212
rect 30044 23158 30046 23210
rect 30098 23158 30100 23210
rect 30044 23146 30100 23158
rect 30156 23212 30212 23660
rect 30716 23660 30996 23716
rect 30380 23492 30436 23502
rect 30156 23210 30324 23212
rect 30156 23158 30158 23210
rect 30210 23158 30324 23210
rect 30156 23156 30324 23158
rect 30156 23146 30212 23156
rect 29932 22418 29988 22428
rect 29484 22372 29540 22382
rect 29484 22278 29540 22316
rect 29708 22372 29764 22382
rect 29708 22370 29876 22372
rect 29708 22318 29710 22370
rect 29762 22318 29876 22370
rect 29708 22316 29876 22318
rect 29708 22306 29764 22316
rect 28812 21756 28980 21812
rect 29708 21812 29764 21822
rect 28588 21476 28644 21486
rect 28364 21474 28644 21476
rect 28364 21422 28590 21474
rect 28642 21422 28644 21474
rect 28364 21420 28644 21422
rect 28364 21026 28420 21420
rect 28588 21410 28644 21420
rect 28364 20974 28366 21026
rect 28418 20974 28420 21026
rect 28364 20962 28420 20974
rect 28812 20916 28868 21756
rect 29484 21252 29540 21262
rect 28812 20860 28980 20916
rect 28700 20804 28756 20814
rect 28700 20710 28756 20748
rect 28084 19796 28140 19806
rect 27916 19794 28140 19796
rect 27916 19742 28086 19794
rect 28138 19742 28140 19794
rect 27916 19740 28140 19742
rect 27580 19572 27636 19582
rect 27356 19460 27412 19470
rect 27356 18696 27412 19404
rect 27580 19346 27636 19516
rect 27580 19294 27582 19346
rect 27634 19294 27636 19346
rect 27580 19282 27636 19294
rect 27300 18674 27412 18696
rect 27300 18622 27302 18674
rect 27354 18622 27412 18674
rect 27300 18610 27412 18622
rect 27132 18386 27188 18396
rect 27356 18340 27412 18610
rect 27916 18564 27972 19740
rect 28084 19730 28140 19740
rect 28140 19460 28196 19470
rect 28140 19234 28196 19404
rect 28140 19182 28142 19234
rect 28194 19182 28196 19234
rect 28140 19170 28196 19182
rect 28252 19236 28308 20076
rect 28812 20132 28868 20142
rect 28812 20074 28868 20076
rect 28364 20046 28420 20058
rect 28364 19994 28366 20046
rect 28418 19994 28420 20046
rect 28364 19572 28420 19994
rect 28364 19506 28420 19516
rect 28588 20046 28644 20058
rect 28588 19994 28590 20046
rect 28642 19994 28644 20046
rect 28812 20022 28814 20074
rect 28866 20022 28868 20074
rect 28812 20010 28868 20022
rect 28924 20074 28980 20860
rect 29204 20804 29260 20814
rect 29204 20710 29260 20748
rect 29484 20774 29540 21196
rect 29484 20722 29486 20774
rect 29538 20722 29540 20774
rect 29484 20710 29540 20722
rect 29708 20774 29764 21756
rect 29820 21364 29876 22316
rect 29988 22258 30044 22270
rect 29988 22206 29990 22258
rect 30042 22206 30044 22258
rect 29988 21812 30044 22206
rect 29988 21746 30044 21756
rect 30156 22148 30212 22158
rect 30156 21588 30212 22092
rect 30268 21924 30324 23156
rect 30268 21858 30324 21868
rect 29820 21298 29876 21308
rect 29932 21532 30212 21588
rect 29708 20722 29710 20774
rect 29762 20722 29764 20774
rect 29708 20710 29764 20722
rect 29932 20774 29988 21532
rect 29932 20722 29934 20774
rect 29986 20722 29988 20774
rect 29932 20710 29988 20722
rect 30044 20746 30100 20758
rect 30044 20694 30046 20746
rect 30098 20694 30100 20746
rect 29596 20580 29652 20590
rect 28924 20022 28926 20074
rect 28978 20022 28980 20074
rect 28476 19348 28532 19358
rect 28588 19348 28644 19994
rect 28924 19684 28980 20022
rect 29148 20356 29204 20366
rect 29148 20018 29204 20300
rect 29484 20132 29540 20142
rect 29148 19966 29150 20018
rect 29202 19966 29204 20018
rect 29148 19954 29204 19966
rect 29260 20076 29484 20132
rect 29260 19908 29316 20076
rect 29484 20038 29540 20076
rect 29260 19684 29316 19852
rect 28924 19618 28980 19628
rect 29148 19628 29316 19684
rect 28476 19346 28588 19348
rect 28476 19294 28478 19346
rect 28530 19294 28588 19346
rect 28476 19292 28588 19294
rect 28476 19282 28532 19292
rect 28588 19254 28644 19292
rect 28308 19204 28364 19236
rect 28308 19180 28310 19204
rect 28252 19152 28310 19180
rect 28362 19152 28364 19204
rect 28252 19142 28364 19152
rect 28308 19140 28364 19142
rect 29148 19199 29204 19628
rect 29596 19460 29652 20524
rect 30044 20356 30100 20694
rect 30044 20290 30100 20300
rect 30268 20244 30324 20254
rect 30380 20244 30436 23436
rect 30548 22596 30604 22606
rect 30548 22148 30604 22540
rect 30548 22054 30604 22092
rect 30604 21924 30660 21934
rect 30492 21474 30548 21486
rect 30492 21422 30494 21474
rect 30546 21422 30548 21474
rect 30492 21364 30548 21422
rect 30492 21298 30548 21308
rect 30604 20926 30660 21868
rect 30548 20914 30660 20926
rect 30548 20862 30550 20914
rect 30602 20862 30660 20914
rect 30548 20860 30660 20862
rect 30716 21588 30772 23660
rect 30884 22932 30940 22942
rect 30884 22838 30940 22876
rect 30716 20916 30772 21532
rect 30940 21812 30996 21822
rect 30940 21586 30996 21756
rect 31052 21700 31108 25228
rect 31164 24836 31220 25788
rect 32452 25732 32508 26182
rect 32452 25676 32564 25732
rect 31724 25396 31780 25406
rect 31612 25394 31780 25396
rect 31612 25342 31726 25394
rect 31778 25342 31780 25394
rect 31612 25340 31780 25342
rect 31164 24770 31220 24780
rect 31407 24836 31463 24846
rect 31407 24778 31463 24780
rect 31276 24724 31332 24734
rect 31407 24726 31409 24778
rect 31461 24726 31463 24778
rect 31407 24714 31463 24726
rect 31612 24724 31668 25340
rect 31724 25330 31780 25340
rect 32508 25396 32564 25676
rect 32844 25630 32900 28364
rect 32508 25330 32564 25340
rect 32788 25618 32900 25630
rect 32788 25566 32790 25618
rect 32842 25566 32900 25618
rect 32788 25564 32900 25566
rect 32340 25284 32396 25294
rect 32340 25190 32396 25228
rect 32788 24836 32844 25564
rect 32956 24948 33012 29708
rect 33572 29652 33628 29662
rect 33572 29558 33628 29596
rect 33404 29428 33460 29438
rect 33516 29428 33572 29438
rect 33964 29428 34020 30158
rect 34300 30154 34356 30166
rect 34300 30102 34302 30154
rect 34354 30102 34356 30154
rect 34300 30100 34356 30102
rect 34188 30042 34244 30054
rect 34188 29990 34190 30042
rect 34242 29990 34244 30042
rect 34076 29876 34132 29886
rect 34076 29594 34132 29820
rect 34076 29542 34078 29594
rect 34130 29542 34132 29594
rect 34076 29530 34132 29542
rect 33404 29426 33516 29428
rect 33404 29374 33406 29426
rect 33458 29374 33516 29426
rect 33404 29372 33516 29374
rect 33404 29362 33460 29372
rect 33348 28868 33404 28878
rect 33348 28774 33404 28812
rect 33068 28644 33124 28654
rect 33068 28550 33124 28588
rect 33516 28644 33572 29372
rect 33852 29426 34020 29428
rect 33852 29374 33966 29426
rect 34018 29374 34020 29426
rect 33852 29372 34020 29374
rect 33516 28308 33572 28588
rect 33292 28252 33572 28308
rect 33628 29316 33684 29326
rect 33124 27636 33180 27646
rect 32956 24882 33012 24892
rect 33068 27634 33180 27636
rect 33068 27582 33126 27634
rect 33178 27582 33180 27634
rect 33068 27570 33180 27582
rect 32788 24770 32844 24780
rect 31164 24498 31220 24510
rect 31164 24446 31166 24498
rect 31218 24446 31220 24498
rect 31164 23940 31220 24446
rect 31164 23874 31220 23884
rect 31164 23154 31220 23166
rect 31164 23102 31166 23154
rect 31218 23102 31220 23154
rect 31164 23044 31220 23102
rect 31276 23154 31332 24668
rect 31612 24658 31668 24668
rect 32284 24724 32340 24762
rect 32284 24658 32340 24668
rect 32620 24052 32676 24062
rect 32620 23938 32676 23996
rect 32620 23886 32622 23938
rect 32674 23886 32676 23938
rect 32620 23874 32676 23886
rect 33068 23940 33124 27570
rect 33292 27412 33348 28252
rect 33404 27860 33460 27870
rect 33404 27766 33460 27804
rect 33628 27858 33684 29260
rect 33852 28420 33908 29372
rect 33964 29362 34020 29372
rect 34188 29316 34244 29990
rect 34300 29652 34356 30044
rect 34300 29586 34356 29596
rect 34636 30158 34638 30210
rect 34690 30158 34692 30210
rect 34300 29453 34356 29466
rect 34300 29428 34302 29453
rect 34354 29428 34356 29453
rect 34636 29428 34692 30158
rect 34300 29362 34356 29372
rect 34412 29372 34636 29428
rect 34188 29250 34244 29260
rect 33852 28354 33908 28364
rect 33964 28756 34020 28766
rect 33964 28532 34020 28700
rect 34300 28644 34356 28654
rect 34412 28644 34468 29372
rect 34636 29334 34692 29372
rect 34300 28642 34468 28644
rect 34300 28590 34302 28642
rect 34354 28590 34468 28642
rect 34300 28588 34468 28590
rect 34524 28644 34580 28654
rect 34300 28578 34356 28588
rect 34524 28551 34526 28588
rect 34578 28551 34580 28588
rect 34524 28539 34580 28551
rect 33964 28476 34244 28532
rect 33628 27806 33630 27858
rect 33682 27806 33684 27858
rect 33628 27794 33684 27806
rect 33740 27860 33796 27870
rect 33740 27766 33796 27804
rect 33964 27858 34020 28476
rect 34188 28474 34244 28476
rect 34188 28422 34190 28474
rect 34242 28422 34244 28474
rect 34188 28410 34244 28422
rect 34244 28308 34300 28318
rect 34244 27970 34300 28252
rect 34244 27918 34246 27970
rect 34298 27918 34300 27970
rect 34244 27906 34300 27918
rect 34748 27860 34804 31052
rect 34972 30994 35028 31006
rect 35196 30996 35252 31006
rect 34972 30942 34974 30994
rect 35026 30942 35028 30994
rect 34972 29988 35028 30942
rect 35084 30994 35252 30996
rect 35084 30942 35198 30994
rect 35250 30942 35252 30994
rect 35084 30940 35252 30942
rect 35532 30996 35588 31948
rect 36204 31958 36260 36092
rect 36316 33348 36372 36652
rect 36540 36484 36596 36494
rect 36540 36390 36596 36428
rect 36428 35252 36484 35262
rect 36428 34914 36484 35196
rect 36428 34862 36430 34914
rect 36482 34862 36484 34914
rect 36428 34850 36484 34862
rect 36652 34356 36708 40796
rect 37156 40628 37212 40910
rect 36764 40430 36820 40442
rect 36764 40404 36766 40430
rect 36818 40404 36820 40430
rect 36764 40338 36820 40348
rect 36988 40430 37044 40442
rect 36988 40404 36990 40430
rect 37042 40404 37044 40430
rect 36988 40338 37044 40348
rect 37156 40292 37212 40572
rect 37436 40852 37492 40862
rect 37268 40516 37324 40526
rect 37268 40422 37324 40460
rect 37324 40292 37380 40302
rect 37156 40236 37268 40292
rect 36764 40180 36820 40190
rect 36764 39396 36820 40124
rect 36988 39620 37044 39630
rect 36988 39531 36990 39564
rect 37042 39531 37044 39564
rect 36988 39519 37044 39531
rect 37100 39562 37156 39574
rect 37100 39510 37102 39562
rect 37154 39510 37156 39562
rect 37100 39396 37156 39510
rect 36764 39340 37156 39396
rect 36764 39060 36820 39340
rect 36876 39172 36932 39182
rect 36932 39116 37044 39172
rect 36876 39106 36932 39116
rect 36764 38994 36820 39004
rect 36876 38948 36932 38958
rect 36876 38890 36932 38892
rect 36764 38869 36820 38881
rect 36764 38817 36766 38869
rect 36818 38817 36820 38869
rect 36876 38838 36878 38890
rect 36930 38838 36932 38890
rect 36876 38826 36932 38838
rect 36764 38724 36820 38817
rect 36764 34468 36820 38668
rect 36876 38052 36932 38062
rect 36876 37958 36932 37996
rect 36988 36708 37044 39116
rect 37100 39060 37156 39070
rect 37100 38890 37156 39004
rect 37100 38838 37102 38890
rect 37154 38838 37156 38890
rect 37100 38836 37156 38838
rect 37100 38760 37156 38780
rect 37212 38668 37268 40236
rect 37324 39590 37380 40236
rect 37324 39538 37326 39590
rect 37378 39538 37380 39590
rect 37324 39060 37380 39538
rect 37436 39508 37492 40796
rect 37548 40402 37604 41356
rect 37660 41186 37716 41356
rect 37660 41134 37662 41186
rect 37714 41134 37716 41186
rect 37660 41122 37716 41134
rect 37548 40350 37550 40402
rect 37602 40350 37604 40402
rect 37548 39732 37604 40350
rect 37884 40628 37940 40638
rect 37884 39854 37940 40572
rect 37828 39842 37940 39854
rect 37828 39790 37830 39842
rect 37882 39790 37940 39842
rect 37828 39788 37940 39790
rect 37828 39778 37884 39788
rect 37548 39666 37604 39676
rect 38108 39732 38164 39742
rect 37772 39620 37828 39630
rect 37548 39562 37604 39574
rect 37548 39510 37550 39562
rect 37602 39510 37604 39562
rect 37548 39508 37604 39510
rect 37436 39452 37604 39508
rect 37324 38994 37380 39004
rect 37362 38850 37418 38862
rect 37362 38798 37364 38850
rect 37416 38836 37418 38850
rect 37604 38836 37660 38874
rect 37416 38798 37492 38836
rect 37362 38780 37492 38798
rect 37212 38612 37380 38668
rect 37212 37826 37268 37838
rect 37212 37774 37214 37826
rect 37266 37774 37268 37826
rect 37212 37266 37268 37774
rect 37212 37214 37214 37266
rect 37266 37214 37268 37266
rect 37212 37202 37268 37214
rect 37100 36708 37156 36718
rect 36988 36706 37156 36708
rect 36988 36654 37102 36706
rect 37154 36654 37156 36706
rect 36988 36652 37156 36654
rect 37100 36642 37156 36652
rect 37100 36036 37156 36046
rect 37100 35725 37156 35980
rect 37324 35924 37380 38612
rect 37436 38612 37492 38780
rect 37604 38770 37660 38780
rect 37436 38546 37492 38556
rect 37772 38050 37828 39564
rect 38108 39618 38164 39676
rect 38108 39566 38110 39618
rect 38162 39566 38164 39618
rect 38108 39554 38164 39566
rect 37996 38836 38052 38846
rect 37996 38742 38052 38780
rect 37772 37998 37774 38050
rect 37826 37998 37828 38050
rect 37772 37986 37828 37998
rect 38220 37492 38276 41580
rect 38332 41412 38388 41422
rect 38332 40402 38388 41356
rect 38556 40740 38612 43260
rect 39228 43204 39284 43374
rect 39228 43138 39284 43148
rect 40124 43314 40180 43652
rect 40124 43262 40126 43314
rect 40178 43262 40180 43314
rect 38332 40350 38334 40402
rect 38386 40350 38388 40402
rect 38332 40338 38388 40350
rect 38444 40684 38612 40740
rect 38668 42756 38724 42766
rect 38444 39172 38500 40684
rect 38668 40628 38724 42700
rect 38556 40572 38724 40628
rect 38780 42754 38836 42766
rect 38780 42702 38782 42754
rect 38834 42702 38836 42754
rect 38780 40628 38836 42702
rect 39788 42756 39844 42766
rect 40124 42756 40180 43262
rect 40348 43092 40404 43596
rect 40460 43540 40516 43550
rect 40460 43446 40516 43484
rect 40348 43036 40516 43092
rect 39788 42754 40180 42756
rect 39788 42702 39790 42754
rect 39842 42702 40180 42754
rect 39788 42700 40180 42702
rect 40348 42754 40404 42766
rect 40348 42702 40350 42754
rect 40402 42702 40404 42754
rect 39788 42690 39844 42700
rect 39116 42530 39172 42542
rect 39116 42478 39118 42530
rect 39170 42478 39172 42530
rect 39116 41412 39172 42478
rect 40348 42084 40404 42702
rect 40460 42586 40516 43036
rect 40460 42534 40462 42586
rect 40514 42534 40516 42586
rect 40460 42522 40516 42534
rect 39676 41970 39732 41982
rect 39676 41918 39678 41970
rect 39730 41918 39732 41970
rect 39116 41346 39172 41356
rect 39340 41860 39396 41870
rect 38556 40068 38612 40572
rect 38780 40562 38836 40572
rect 39340 40628 39396 41804
rect 39340 40562 39396 40572
rect 39676 40516 39732 41918
rect 40236 41972 40292 41982
rect 40012 41746 40068 41758
rect 40012 41694 40014 41746
rect 40066 41694 40068 41746
rect 39900 41158 39956 41170
rect 39900 41106 39902 41158
rect 39954 41106 39956 41158
rect 39900 40964 39956 41106
rect 39900 40898 39956 40908
rect 39676 40450 39732 40460
rect 38556 40012 38724 40068
rect 38668 39844 38724 40012
rect 40012 39956 40068 41694
rect 40124 41186 40180 41198
rect 40124 41134 40126 41186
rect 40178 41134 40180 41186
rect 40124 40740 40180 41134
rect 40124 40674 40180 40684
rect 40236 40852 40292 41916
rect 40236 40514 40292 40796
rect 40236 40462 40238 40514
rect 40290 40462 40292 40514
rect 40236 40450 40292 40462
rect 38668 39778 38724 39788
rect 38892 39900 40068 39956
rect 38892 39730 38948 39900
rect 38892 39678 38894 39730
rect 38946 39678 38948 39730
rect 38892 39666 38948 39678
rect 38444 39106 38500 39116
rect 38948 38724 39004 38734
rect 38948 38630 39004 38668
rect 38332 38610 38388 38622
rect 38332 38558 38334 38610
rect 38386 38558 38388 38610
rect 38332 38164 38388 38558
rect 38556 38164 38612 38174
rect 38332 38162 38612 38164
rect 38332 38110 38558 38162
rect 38610 38110 38612 38162
rect 38332 38108 38612 38110
rect 38556 38098 38612 38108
rect 39116 37828 39172 37838
rect 38220 37436 38500 37492
rect 37436 36484 37492 36494
rect 38276 36484 38332 36494
rect 37436 36482 38332 36484
rect 37436 36430 37438 36482
rect 37490 36430 38278 36482
rect 38330 36430 38332 36482
rect 37436 36428 38332 36430
rect 37436 36418 37492 36428
rect 37828 36258 37884 36270
rect 37828 36206 37830 36258
rect 37882 36206 37884 36258
rect 37828 36036 37884 36206
rect 37828 35970 37884 35980
rect 37324 35868 37492 35924
rect 37100 35673 37102 35725
rect 37154 35673 37156 35725
rect 37100 35364 37156 35673
rect 37324 35700 37380 35738
rect 37324 35634 37380 35644
rect 37324 35476 37380 35486
rect 37100 35308 37268 35364
rect 36932 34867 36988 34879
rect 36932 34815 36934 34867
rect 36986 34815 36988 34867
rect 36932 34804 36988 34815
rect 36932 34738 36988 34748
rect 36764 34402 36820 34412
rect 36652 34290 36708 34300
rect 37100 33796 37156 33806
rect 36316 33292 36708 33348
rect 36372 33124 36428 33134
rect 36372 33030 36428 33068
rect 36540 33124 36596 33134
rect 36316 32788 36372 32798
rect 36316 32562 36372 32732
rect 36316 32510 36318 32562
rect 36370 32510 36372 32562
rect 36316 32498 36372 32510
rect 36204 31946 36316 31958
rect 36204 31894 36262 31946
rect 36314 31894 36316 31946
rect 36204 31892 36316 31894
rect 36260 31882 36316 31892
rect 36092 31778 36148 31790
rect 36092 31726 36094 31778
rect 36146 31726 36148 31778
rect 35756 31668 35812 31678
rect 36092 31668 36148 31726
rect 35756 31666 36148 31668
rect 35756 31614 35758 31666
rect 35810 31614 36148 31666
rect 35756 31612 36148 31614
rect 35756 31444 35812 31612
rect 35756 31378 35812 31388
rect 35756 30996 35812 31006
rect 35532 30994 35812 30996
rect 35532 30942 35758 30994
rect 35810 30942 35812 30994
rect 35532 30940 35812 30942
rect 35084 30436 35140 30940
rect 35196 30930 35252 30940
rect 35756 30930 35812 30940
rect 36540 30994 36596 33068
rect 36540 30942 36542 30994
rect 36594 30942 36596 30994
rect 36540 30930 36596 30942
rect 35476 30772 35532 30810
rect 36652 30772 36708 33292
rect 35476 30706 35532 30716
rect 35756 30716 36708 30772
rect 36764 33012 36820 33022
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35084 30380 35364 30436
rect 35196 30212 35252 30222
rect 34972 29922 35028 29932
rect 35084 30210 35252 30212
rect 35084 30158 35198 30210
rect 35250 30158 35252 30210
rect 35084 30156 35252 30158
rect 35084 28868 35140 30156
rect 35196 30146 35252 30156
rect 35308 30212 35364 30380
rect 35308 30042 35364 30156
rect 35308 29990 35310 30042
rect 35362 29990 35364 30042
rect 35532 30154 35588 30166
rect 35532 30102 35534 30154
rect 35586 30102 35588 30154
rect 35532 30100 35588 30102
rect 35532 30034 35588 30044
rect 35308 29978 35364 29990
rect 35364 29652 35420 29662
rect 35364 29558 35420 29596
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35364 28868 35420 28878
rect 34972 28866 35420 28868
rect 34972 28814 35366 28866
rect 35418 28814 35420 28866
rect 34972 28812 35420 28814
rect 34972 28642 35028 28812
rect 35364 28802 35420 28812
rect 35644 28868 35700 28878
rect 34972 28590 34974 28642
rect 35026 28590 35028 28642
rect 34972 28578 35028 28590
rect 35196 28642 35252 28654
rect 35196 28590 35198 28642
rect 35250 28590 35252 28642
rect 33964 27806 33966 27858
rect 34018 27806 34020 27858
rect 33964 27794 34020 27806
rect 34636 27804 34804 27860
rect 34972 28420 35028 28430
rect 35196 28420 35252 28590
rect 35028 28364 35252 28420
rect 33180 27356 33348 27412
rect 33852 27748 33908 27758
rect 33180 26290 33236 27356
rect 33180 26238 33182 26290
rect 33234 26238 33236 26290
rect 33180 25284 33236 26238
rect 33292 27076 33348 27086
rect 33292 26290 33348 27020
rect 33516 27076 33572 27086
rect 33516 26982 33572 27020
rect 33852 27074 33908 27692
rect 33852 27022 33854 27074
rect 33906 27022 33908 27074
rect 33852 27010 33908 27022
rect 34076 27074 34132 27086
rect 34076 27022 34078 27074
rect 34130 27022 34132 27074
rect 34076 26964 34132 27022
rect 34188 27076 34244 27086
rect 34188 26982 34244 27020
rect 34468 27076 34524 27114
rect 34468 27010 34524 27020
rect 34636 26908 34692 27804
rect 34748 27636 34804 27646
rect 34748 27634 34916 27636
rect 34748 27582 34750 27634
rect 34802 27582 34916 27634
rect 34748 27580 34916 27582
rect 34748 27570 34804 27580
rect 34748 27076 34804 27086
rect 34748 26982 34804 27020
rect 34076 26898 34132 26908
rect 33292 26238 33294 26290
rect 33346 26238 33348 26290
rect 33292 26226 33348 26238
rect 33852 26852 33908 26862
rect 33572 26068 33628 26078
rect 33572 25974 33628 26012
rect 33852 25506 33908 26796
rect 34524 26852 34692 26908
rect 34188 26740 34244 26750
rect 34076 26328 34132 26340
rect 34076 26292 34078 26328
rect 34130 26292 34132 26328
rect 34188 26292 34244 26684
rect 33852 25454 33854 25506
rect 33906 25454 33908 25506
rect 33852 25442 33908 25454
rect 33964 26234 34020 26246
rect 33964 26182 33966 26234
rect 34018 26182 34020 26234
rect 34132 26236 34244 26292
rect 34076 26226 34132 26236
rect 33516 25396 33572 25406
rect 33180 25218 33236 25228
rect 33348 25284 33404 25294
rect 33516 25284 33572 25340
rect 33348 25282 33572 25284
rect 33348 25230 33350 25282
rect 33402 25230 33572 25282
rect 33348 25228 33572 25230
rect 33348 25218 33404 25228
rect 33516 25060 33572 25228
rect 33684 25284 33740 25294
rect 33964 25284 34020 26182
rect 34188 25468 34244 26236
rect 34524 25732 34580 26852
rect 34860 26740 34916 27580
rect 34972 27524 35028 28364
rect 35084 27858 35140 27870
rect 35084 27806 35086 27858
rect 35138 27806 35140 27858
rect 35084 27748 35140 27806
rect 35084 27682 35140 27692
rect 34972 27468 35140 27524
rect 34860 26674 34916 26684
rect 34972 27074 35028 27086
rect 34972 27022 34974 27074
rect 35026 27022 35028 27074
rect 34972 26516 35028 27022
rect 35084 26964 35140 27468
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35252 27076 35308 27086
rect 35532 27076 35588 27086
rect 35252 27074 35588 27076
rect 35252 27022 35254 27074
rect 35306 27022 35534 27074
rect 35586 27022 35588 27074
rect 35252 27020 35588 27022
rect 35252 27010 35308 27020
rect 35532 27010 35588 27020
rect 35644 26908 35700 28812
rect 35084 26852 35364 26908
rect 34636 26460 35028 26516
rect 34636 26402 34692 26460
rect 34636 26350 34638 26402
rect 34690 26350 34692 26402
rect 34636 26338 34692 26350
rect 35308 26402 35364 26852
rect 35308 26350 35310 26402
rect 35362 26350 35364 26402
rect 35308 26338 35364 26350
rect 35532 26852 35700 26908
rect 34804 26234 34860 26246
rect 34804 26182 34806 26234
rect 34858 26182 34860 26234
rect 34804 26068 34860 26182
rect 35084 26068 35140 26078
rect 34804 26012 34972 26068
rect 34524 25676 34692 25732
rect 34524 25508 34580 25518
rect 34188 25416 34190 25468
rect 34242 25416 34244 25468
rect 34188 25404 34244 25416
rect 34300 25506 34580 25508
rect 34300 25454 34526 25506
rect 34578 25454 34580 25506
rect 34300 25452 34580 25454
rect 33684 25282 34020 25284
rect 33684 25230 33686 25282
rect 33738 25230 34020 25282
rect 33684 25228 34020 25230
rect 33684 25218 33740 25228
rect 33516 25004 33684 25060
rect 33180 24948 33236 24958
rect 33180 24854 33236 24892
rect 33516 24722 33572 24734
rect 33516 24670 33518 24722
rect 33570 24670 33572 24722
rect 33516 24500 33572 24670
rect 33628 24612 33684 25004
rect 34300 24958 34356 25452
rect 34524 25442 34580 25452
rect 34244 24946 34356 24958
rect 34244 24894 34246 24946
rect 34298 24894 34356 24946
rect 34244 24892 34356 24894
rect 34244 24882 34300 24892
rect 34076 24724 34132 24734
rect 34076 24630 34132 24668
rect 34636 24724 34692 25676
rect 34748 25508 34804 25518
rect 34748 25414 34804 25452
rect 34916 25450 34972 26012
rect 34916 25398 34918 25450
rect 34970 25398 34972 25450
rect 35084 25506 35140 26012
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35532 25732 35588 26852
rect 35420 25676 35588 25732
rect 35084 25454 35086 25506
rect 35138 25454 35140 25506
rect 35084 25442 35140 25454
rect 35308 25508 35364 25518
rect 35308 25414 35364 25452
rect 34916 25396 34972 25398
rect 34916 25330 34972 25340
rect 35308 25284 35364 25294
rect 35308 24834 35364 25228
rect 35308 24782 35310 24834
rect 35362 24782 35364 24834
rect 35308 24770 35364 24782
rect 34916 24724 34972 24734
rect 34692 24668 34804 24724
rect 34636 24658 34692 24668
rect 33908 24612 33964 24622
rect 33628 24610 33964 24612
rect 33628 24558 33910 24610
rect 33962 24558 33964 24610
rect 33628 24556 33964 24558
rect 33292 23940 33348 23950
rect 33068 23938 33348 23940
rect 33068 23886 33294 23938
rect 33346 23886 33348 23938
rect 33068 23884 33348 23886
rect 33516 23940 33572 24444
rect 33908 24388 33964 24556
rect 34580 24388 34636 24398
rect 33908 24332 34356 24388
rect 34076 24052 34132 24062
rect 33628 23940 33684 23950
rect 33516 23938 33684 23940
rect 33516 23886 33630 23938
rect 33682 23886 33684 23938
rect 33908 23912 33964 23920
rect 33516 23884 33684 23886
rect 31724 23826 31780 23838
rect 31724 23774 31726 23826
rect 31778 23774 31780 23826
rect 31724 23492 31780 23774
rect 32284 23716 32340 23726
rect 31724 23426 31780 23436
rect 32172 23714 32340 23716
rect 32172 23662 32286 23714
rect 32338 23662 32340 23714
rect 32172 23660 32340 23662
rect 32172 23380 32228 23660
rect 32284 23650 32340 23660
rect 32956 23714 33012 23726
rect 32956 23662 32958 23714
rect 33010 23662 33012 23714
rect 32172 23210 32228 23324
rect 32956 23380 33012 23662
rect 33292 23716 33348 23884
rect 33628 23874 33684 23884
rect 33852 23908 33964 23912
rect 33852 23856 33910 23908
rect 33962 23856 33964 23908
rect 33852 23844 33964 23856
rect 33852 23716 33908 23844
rect 33292 23660 33908 23716
rect 32956 23314 33012 23324
rect 31948 23182 32004 23194
rect 31276 23102 31278 23154
rect 31330 23102 31332 23154
rect 31276 23090 31332 23102
rect 31668 23156 31724 23166
rect 31668 23062 31724 23100
rect 31948 23130 31950 23182
rect 32002 23130 32004 23182
rect 32172 23158 32174 23210
rect 32226 23158 32228 23210
rect 32172 23146 32228 23158
rect 32396 23268 32452 23278
rect 32620 23268 32676 23278
rect 32396 23210 32452 23212
rect 32396 23158 32398 23210
rect 32450 23158 32452 23210
rect 32396 23146 32452 23158
rect 32583 23212 32620 23222
rect 32583 23210 32676 23212
rect 32583 23158 32585 23210
rect 32637 23158 32676 23210
rect 32583 23156 32676 23158
rect 32956 23156 33012 23166
rect 32583 23146 32639 23156
rect 31164 22482 31220 22988
rect 31948 23044 32004 23130
rect 32956 23062 33012 23100
rect 33516 23156 33572 23166
rect 31948 22978 32004 22988
rect 31164 22430 31166 22482
rect 31218 22430 31220 22482
rect 31164 22418 31220 22430
rect 31500 22932 31556 22942
rect 33292 22932 33348 22942
rect 31276 21700 31332 21710
rect 31052 21644 31220 21700
rect 30940 21534 30942 21586
rect 30994 21534 30996 21586
rect 30940 21522 30996 21534
rect 30548 20850 30604 20860
rect 30716 20850 30772 20860
rect 30380 20188 30548 20244
rect 30268 20132 30324 20188
rect 30156 20076 30324 20132
rect 30156 20074 30212 20076
rect 30156 20022 30158 20074
rect 30210 20022 30212 20074
rect 30156 20010 30212 20022
rect 30380 20018 30436 20030
rect 30380 19966 30382 20018
rect 30434 19966 30436 20018
rect 29596 19394 29652 19404
rect 29708 19796 29764 19806
rect 29484 19348 29540 19358
rect 29148 19147 29150 19199
rect 29202 19147 29204 19199
rect 29148 19135 29204 19147
rect 29260 19236 29316 19246
rect 29260 19154 29262 19180
rect 29314 19154 29316 19180
rect 29260 19142 29316 19154
rect 29484 19206 29540 19292
rect 29484 19154 29486 19206
rect 29538 19154 29540 19206
rect 29484 19142 29540 19154
rect 29708 19206 29764 19740
rect 30380 19796 30436 19966
rect 30380 19730 30436 19740
rect 30156 19684 30212 19694
rect 30492 19684 30548 20188
rect 31052 20020 31108 20030
rect 30772 19962 30828 19974
rect 30156 19460 30212 19628
rect 30156 19394 30212 19404
rect 30488 19628 30548 19684
rect 30604 19906 30660 19918
rect 30604 19854 30606 19906
rect 30658 19854 30660 19906
rect 29708 19154 29710 19206
rect 29762 19154 29764 19206
rect 29708 19142 29764 19154
rect 30488 19196 30544 19628
rect 30488 19144 30490 19196
rect 30542 19144 30544 19196
rect 28588 19124 28644 19134
rect 27916 18498 27972 18508
rect 28028 18788 28084 18798
rect 28028 18450 28084 18732
rect 28028 18398 28030 18450
rect 28082 18398 28084 18450
rect 28028 18386 28084 18398
rect 28140 18452 28196 18462
rect 28140 18450 28308 18452
rect 28140 18398 28142 18450
rect 28194 18398 28308 18450
rect 28140 18396 28308 18398
rect 28140 18386 28196 18396
rect 27356 18274 27412 18284
rect 27692 18340 27748 18350
rect 27692 18246 27748 18284
rect 26236 17780 26292 17790
rect 25844 17778 26292 17780
rect 25844 17726 26238 17778
rect 26290 17726 26292 17778
rect 25844 17724 26292 17726
rect 25844 17666 25900 17724
rect 26236 17714 26292 17724
rect 26348 17780 26404 17790
rect 25844 17614 25846 17666
rect 25898 17614 25900 17666
rect 25844 17602 25900 17614
rect 25564 17154 25620 17164
rect 25676 17554 25732 17566
rect 25676 17502 25678 17554
rect 25730 17502 25732 17554
rect 25452 16322 25564 16334
rect 25452 16270 25510 16322
rect 25562 16270 25564 16322
rect 25452 16268 25564 16270
rect 25508 16258 25564 16268
rect 25676 16212 25732 17502
rect 25676 16146 25732 16156
rect 25788 17444 25844 17454
rect 25340 16098 25396 16110
rect 25340 16046 25342 16098
rect 25394 16046 25396 16098
rect 24780 15708 24948 15764
rect 25116 15988 25172 15998
rect 24668 15652 24724 15662
rect 24500 15540 24556 15550
rect 24500 15446 24556 15484
rect 24332 15428 24388 15438
rect 24332 15314 24388 15372
rect 24332 15262 24334 15314
rect 24386 15262 24388 15314
rect 24332 15250 24388 15262
rect 23772 13750 23774 13802
rect 23826 13750 23828 13802
rect 23772 13738 23828 13750
rect 23970 14252 24276 14308
rect 23970 13786 24026 14252
rect 23970 13734 23972 13786
rect 24024 13734 24026 13786
rect 23970 13722 24026 13734
rect 24668 13748 24724 15596
rect 24668 13682 24724 13692
rect 23548 13580 23828 13636
rect 23436 12910 23438 12962
rect 23490 12910 23492 12962
rect 23436 12898 23492 12910
rect 22764 12124 23044 12180
rect 22988 11956 23044 12124
rect 23100 12178 23268 12180
rect 23100 12126 23102 12178
rect 23154 12126 23268 12178
rect 23772 12234 23828 13580
rect 23772 12182 23774 12234
rect 23826 12182 23828 12234
rect 23772 12170 23828 12182
rect 23996 13634 24052 13646
rect 23996 13582 23998 13634
rect 24050 13582 24052 13634
rect 23996 12234 24052 13582
rect 24108 13524 24164 13534
rect 24108 12404 24164 13468
rect 24780 13300 24836 15708
rect 25116 15314 25172 15932
rect 25116 15262 25118 15314
rect 25170 15262 25172 15314
rect 25116 15250 25172 15262
rect 24892 15204 24948 15214
rect 25340 15148 25396 16046
rect 24892 15092 25396 15148
rect 25564 16100 25620 16110
rect 25452 15092 25508 15102
rect 24892 14642 24948 15092
rect 25452 14998 25508 15036
rect 24892 14590 24894 14642
rect 24946 14590 24948 14642
rect 24892 14578 24948 14590
rect 25564 14308 25620 16044
rect 25788 15148 25844 17388
rect 26348 16938 26404 17724
rect 26796 17668 26852 17678
rect 26630 17610 26686 17622
rect 26630 17558 26632 17610
rect 26684 17558 26686 17610
rect 26796 17574 26852 17612
rect 26908 17666 26964 17678
rect 26908 17614 26910 17666
rect 26962 17614 26964 17666
rect 26630 17332 26686 17558
rect 26630 17266 26686 17276
rect 26908 17108 26964 17614
rect 26348 16886 26350 16938
rect 26402 16886 26404 16938
rect 26348 16874 26404 16886
rect 26572 17052 26964 17108
rect 27020 17668 27076 17678
rect 27020 17108 27076 17612
rect 27692 17668 27748 17678
rect 28084 17668 28140 17678
rect 27692 17666 28140 17668
rect 27692 17614 27694 17666
rect 27746 17614 28086 17666
rect 28138 17614 28140 17666
rect 27692 17612 28140 17614
rect 27244 17444 27300 17454
rect 26572 16882 26628 17052
rect 27020 17042 27076 17052
rect 27132 17220 27188 17230
rect 26572 16830 26574 16882
rect 26626 16830 26628 16882
rect 26012 15986 26068 15998
rect 26012 15934 26014 15986
rect 26066 15934 26068 15986
rect 26012 15316 26068 15934
rect 26404 15540 26460 15550
rect 26572 15540 26628 16830
rect 26796 16884 26852 16894
rect 26796 16790 26852 16828
rect 26964 16884 27020 16894
rect 26964 16790 27020 16828
rect 27132 16660 27188 17164
rect 27244 16882 27300 17388
rect 27356 17442 27412 17454
rect 27356 17390 27358 17442
rect 27410 17390 27412 17442
rect 27356 17332 27412 17390
rect 27542 17332 27598 17342
rect 27356 17276 27542 17332
rect 27244 16830 27246 16882
rect 27298 16830 27300 16882
rect 27244 16818 27300 16830
rect 27356 17108 27412 17118
rect 27356 16882 27412 17052
rect 27356 16830 27358 16882
rect 27410 16830 27412 16882
rect 27542 16920 27598 17276
rect 27692 17220 27748 17612
rect 28084 17602 28140 17612
rect 27692 17154 27748 17164
rect 27542 16868 27544 16920
rect 27596 16868 27598 16920
rect 27542 16856 27598 16868
rect 27916 16884 27972 16894
rect 27356 16818 27412 16830
rect 27916 16770 27972 16828
rect 27916 16718 27918 16770
rect 27970 16718 27972 16770
rect 27916 16706 27972 16718
rect 26404 15538 26628 15540
rect 26404 15486 26406 15538
rect 26458 15486 26628 15538
rect 26404 15484 26628 15486
rect 26684 16604 27188 16660
rect 26404 15474 26460 15484
rect 26012 15250 26068 15260
rect 26236 15316 26292 15326
rect 26236 15222 26292 15260
rect 25526 14252 25620 14308
rect 25676 15092 25844 15148
rect 25526 13784 25582 14252
rect 25228 13746 25284 13758
rect 25228 13694 25230 13746
rect 25282 13694 25284 13746
rect 25228 13412 25284 13694
rect 25340 13748 25396 13758
rect 25526 13732 25528 13784
rect 25580 13732 25582 13784
rect 25526 13720 25582 13732
rect 25340 13654 25396 13692
rect 25228 13346 25284 13356
rect 24780 13234 24836 13244
rect 25452 13076 25508 13086
rect 24220 12964 24276 12974
rect 24220 12962 24500 12964
rect 24220 12910 24222 12962
rect 24274 12910 24500 12962
rect 24220 12908 24500 12910
rect 24220 12898 24276 12908
rect 24108 12348 24388 12404
rect 23996 12182 23998 12234
rect 24050 12182 24052 12234
rect 23996 12170 24052 12182
rect 23100 12124 23268 12126
rect 23100 12114 23156 12124
rect 23492 12122 23548 12134
rect 23324 12066 23380 12078
rect 23324 12014 23326 12066
rect 23378 12014 23380 12066
rect 22988 11900 23156 11956
rect 21084 11620 21140 11630
rect 21644 11618 21756 11630
rect 21644 11566 21702 11618
rect 21754 11566 21756 11618
rect 21644 11564 21756 11566
rect 21084 10846 21140 11564
rect 21700 11554 21756 11564
rect 21980 11396 22036 11406
rect 21980 11302 22036 11340
rect 22092 11394 22148 11406
rect 22092 11342 22094 11394
rect 22146 11342 22148 11394
rect 22092 11284 22148 11342
rect 22092 11218 22148 11228
rect 22764 11394 22820 11406
rect 22764 11342 22766 11394
rect 22818 11342 22820 11394
rect 21084 10834 21196 10846
rect 21084 10782 21142 10834
rect 21194 10782 21196 10834
rect 21084 10780 21196 10782
rect 21140 10770 21196 10780
rect 21678 10836 21734 10846
rect 20972 10658 21028 10668
rect 21532 10724 21588 10734
rect 20524 10558 20526 10610
rect 20578 10558 20580 10610
rect 20524 10546 20580 10558
rect 20636 10612 20692 10622
rect 20636 10518 20692 10556
rect 21420 10610 21476 10622
rect 21420 10558 21422 10610
rect 21474 10558 21476 10610
rect 19292 10434 19348 10444
rect 21420 10500 21476 10558
rect 21532 10610 21588 10668
rect 21532 10558 21534 10610
rect 21586 10558 21588 10610
rect 21532 10546 21588 10558
rect 21678 10648 21734 10780
rect 21678 10596 21680 10648
rect 21732 10596 21734 10648
rect 21420 10434 21476 10444
rect 19404 10386 19460 10398
rect 19964 10388 20020 10398
rect 19404 10334 19406 10386
rect 19458 10334 19460 10386
rect 19292 9828 19348 9838
rect 19292 9734 19348 9772
rect 19404 9492 19460 10334
rect 19684 10386 20020 10388
rect 19684 10334 19966 10386
rect 20018 10334 20020 10386
rect 19684 10332 20020 10334
rect 19684 9882 19740 10332
rect 19964 10322 20020 10332
rect 20412 10388 20468 10398
rect 21678 10388 21734 10596
rect 21980 10724 22036 10734
rect 21678 10332 21868 10388
rect 19684 9830 19686 9882
rect 19738 9830 19740 9882
rect 19684 9818 19740 9830
rect 20188 10276 20244 10286
rect 20188 9798 20244 10220
rect 20188 9746 20190 9798
rect 20242 9746 20244 9798
rect 20412 9826 20468 10332
rect 21420 9940 21476 9950
rect 20412 9774 20414 9826
rect 20466 9774 20468 9826
rect 20412 9762 20468 9774
rect 20804 9938 21476 9940
rect 20804 9886 21422 9938
rect 21474 9886 21476 9938
rect 20804 9884 21476 9886
rect 20804 9826 20860 9884
rect 21420 9874 21476 9884
rect 20804 9774 20806 9826
rect 20858 9774 20860 9826
rect 20804 9762 20860 9774
rect 21812 9826 21868 10332
rect 21812 9774 21814 9826
rect 21866 9774 21868 9826
rect 21812 9762 21868 9774
rect 21980 9826 22036 10668
rect 22484 10610 22540 10622
rect 22484 10558 22486 10610
rect 22538 10558 22540 10610
rect 22092 10500 22148 10510
rect 22484 10500 22540 10558
rect 22092 10498 22540 10500
rect 22092 10446 22094 10498
rect 22146 10446 22540 10498
rect 22092 10444 22540 10446
rect 22652 10498 22708 10510
rect 22652 10446 22654 10498
rect 22706 10446 22708 10498
rect 22092 10434 22148 10444
rect 22652 9940 22708 10446
rect 22652 9874 22708 9884
rect 21980 9774 21982 9826
rect 22034 9774 22036 9826
rect 21980 9762 22036 9774
rect 22092 9828 22148 9838
rect 20188 9734 20244 9746
rect 19516 9716 19572 9726
rect 19516 9622 19572 9660
rect 20636 9716 20692 9754
rect 22092 9734 22148 9772
rect 22316 9826 22372 9838
rect 22316 9774 22318 9826
rect 22370 9774 22372 9826
rect 20636 9650 20692 9660
rect 21308 9716 21364 9726
rect 20636 9492 20692 9502
rect 19404 9436 19628 9492
rect 19404 9268 19460 9278
rect 19404 9154 19460 9212
rect 19404 9102 19406 9154
rect 19458 9102 19460 9154
rect 19404 9090 19460 9102
rect 19572 9098 19628 9436
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19068 9042 19236 9044
rect 18116 8754 18172 8764
rect 17612 8530 17668 8540
rect 17612 8034 17668 8046
rect 17612 7982 17614 8034
rect 17666 7982 17668 8034
rect 17612 7476 17668 7982
rect 17276 6470 17278 6522
rect 17330 6470 17332 6522
rect 17276 6458 17332 6470
rect 17500 7474 17668 7476
rect 17500 7422 17614 7474
rect 17666 7422 17668 7474
rect 17500 7420 17668 7422
rect 16940 6300 17444 6356
rect 15708 6076 16212 6132
rect 15372 5906 15428 5918
rect 15372 5854 15374 5906
rect 15426 5854 15428 5906
rect 15036 5684 15092 5694
rect 14812 5682 15092 5684
rect 14812 5630 15038 5682
rect 15090 5630 15092 5682
rect 14812 5628 15092 5630
rect 14812 5234 14868 5628
rect 15036 5618 15092 5628
rect 15372 5460 15428 5854
rect 15708 5906 15764 6076
rect 15708 5854 15710 5906
rect 15762 5854 15764 5906
rect 15708 5842 15764 5854
rect 15932 5921 15988 5946
rect 15932 5908 15934 5921
rect 15986 5908 15988 5921
rect 16156 5908 16212 6076
rect 16380 5908 16436 5918
rect 16156 5906 16436 5908
rect 16156 5854 16382 5906
rect 16434 5854 16436 5906
rect 16156 5852 16436 5854
rect 15932 5842 15988 5852
rect 16044 5796 16100 5806
rect 16044 5794 16212 5796
rect 16044 5742 16046 5794
rect 16098 5742 16212 5794
rect 16044 5740 16212 5742
rect 16044 5730 16100 5740
rect 15372 5404 15988 5460
rect 14812 5182 14814 5234
rect 14866 5182 14868 5234
rect 14812 5170 14868 5182
rect 15932 5236 15988 5404
rect 15932 5180 16100 5236
rect 14028 5030 14084 5068
rect 15372 4900 15428 4910
rect 8876 4398 8878 4450
rect 8930 4398 8932 4450
rect 8876 4386 8932 4398
rect 14364 4564 14420 4574
rect 8316 4274 8372 4284
rect 14364 4338 14420 4508
rect 15372 4562 15428 4844
rect 15372 4510 15374 4562
rect 15426 4510 15428 4562
rect 15372 4498 15428 4510
rect 16044 4506 16100 5180
rect 15708 4452 15764 4462
rect 16044 4454 16046 4506
rect 16098 4454 16100 4506
rect 16044 4442 16100 4454
rect 16156 4452 16212 5740
rect 16268 5460 16324 5470
rect 16268 4564 16324 5404
rect 16380 5348 16436 5852
rect 16380 5282 16436 5292
rect 16492 5908 16548 5918
rect 16268 4508 16436 4564
rect 16156 4396 16268 4452
rect 14364 4286 14366 4338
rect 14418 4286 14420 4338
rect 14364 4274 14420 4286
rect 15036 4340 15092 4350
rect 15036 4246 15092 4284
rect 15708 4338 15764 4396
rect 16212 4394 16268 4396
rect 15708 4286 15710 4338
rect 15762 4286 15764 4338
rect 15708 4274 15764 4286
rect 16044 4338 16100 4350
rect 16044 4286 16046 4338
rect 16098 4286 16100 4338
rect 16212 4342 16214 4394
rect 16266 4342 16268 4394
rect 16212 4330 16268 4342
rect 16044 4228 16100 4286
rect 16380 4228 16436 4508
rect 16044 4172 16436 4228
rect 16492 4228 16548 5852
rect 16604 5460 16660 6300
rect 16940 6132 16996 6142
rect 16772 5684 16884 5694
rect 16772 5682 16828 5684
rect 16772 5630 16774 5682
rect 16826 5630 16828 5682
rect 16772 5628 16828 5630
rect 16772 5618 16884 5628
rect 16604 5394 16660 5404
rect 16716 5348 16772 5358
rect 16716 5234 16772 5292
rect 16716 5182 16718 5234
rect 16770 5182 16772 5234
rect 16716 5170 16772 5182
rect 16828 5012 16884 5618
rect 16716 4956 16884 5012
rect 16940 5124 16996 6076
rect 17388 5794 17444 6300
rect 17500 6132 17556 7420
rect 17612 7410 17668 7420
rect 17500 6066 17556 6076
rect 17612 6692 17668 6702
rect 17388 5742 17390 5794
rect 17442 5742 17444 5794
rect 17388 5730 17444 5742
rect 17500 5921 17556 5933
rect 17500 5869 17502 5921
rect 17554 5869 17556 5921
rect 17500 5684 17556 5869
rect 17612 5908 17668 6636
rect 17836 6690 17892 6702
rect 17836 6638 17838 6690
rect 17890 6638 17892 6690
rect 17724 5908 17780 5918
rect 17612 5906 17780 5908
rect 17612 5854 17726 5906
rect 17778 5854 17780 5906
rect 17612 5852 17780 5854
rect 17724 5842 17780 5852
rect 17500 5618 17556 5628
rect 17836 5684 17892 6638
rect 18284 6692 18340 8876
rect 19068 8990 19182 9042
rect 19234 8990 19236 9042
rect 19572 9046 19574 9098
rect 19626 9046 19628 9098
rect 19908 9210 19964 9222
rect 19908 9158 19910 9210
rect 19962 9158 19964 9210
rect 19908 9156 19964 9158
rect 19908 9090 19964 9100
rect 19572 9034 19628 9046
rect 19740 9044 19796 9054
rect 19068 8988 19236 8990
rect 18620 8260 18676 8270
rect 18620 8178 18622 8204
rect 18674 8178 18676 8204
rect 18620 8166 18676 8178
rect 18396 8036 18452 8046
rect 18396 7474 18452 7980
rect 19068 7700 19124 8988
rect 19180 8978 19236 8988
rect 19740 8950 19796 8988
rect 20524 9044 20580 9054
rect 20636 9044 20692 9436
rect 20524 9042 20692 9044
rect 20524 8990 20526 9042
rect 20578 8990 20692 9042
rect 20524 8988 20692 8990
rect 20524 8978 20580 8988
rect 18396 7422 18398 7474
rect 18450 7422 18452 7474
rect 18396 7410 18452 7422
rect 18620 7644 19124 7700
rect 19404 8372 19460 8382
rect 19404 7700 19460 8316
rect 20188 8372 20244 8382
rect 19852 8258 19908 8270
rect 19852 8206 19854 8258
rect 19906 8206 19908 8258
rect 19572 8148 19628 8158
rect 19852 8148 19908 8206
rect 19572 8146 19684 8148
rect 19572 8094 19574 8146
rect 19626 8094 19684 8146
rect 19572 8082 19684 8094
rect 19852 8082 19908 8092
rect 20076 8258 20132 8270
rect 20076 8206 20078 8258
rect 20130 8206 20132 8258
rect 19628 7700 19684 8082
rect 20076 8036 20132 8206
rect 20188 8258 20244 8316
rect 20188 8206 20190 8258
rect 20242 8206 20244 8258
rect 20188 8194 20244 8206
rect 20412 8148 20468 8158
rect 20076 7980 20356 8036
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19404 7644 19572 7700
rect 19628 7644 19908 7700
rect 18396 6692 18452 6702
rect 18620 6692 18676 7644
rect 19404 6804 19460 6814
rect 18284 6690 18452 6692
rect 18284 6638 18398 6690
rect 18450 6638 18452 6690
rect 18284 6636 18452 6638
rect 18396 6626 18452 6636
rect 18564 6636 18676 6692
rect 19068 6690 19124 6702
rect 19068 6638 19070 6690
rect 19122 6638 19124 6690
rect 18116 6580 18172 6590
rect 18116 6486 18172 6524
rect 18564 6522 18620 6636
rect 18564 6470 18566 6522
rect 18618 6470 18620 6522
rect 18564 6458 18620 6470
rect 19068 6356 19124 6638
rect 19404 6651 19460 6748
rect 19404 6599 19406 6651
rect 19458 6599 19460 6651
rect 19404 6587 19460 6599
rect 19516 6522 19572 7644
rect 19740 7476 19796 7486
rect 19628 6692 19684 6702
rect 19628 6598 19684 6636
rect 19516 6470 19518 6522
rect 19570 6470 19572 6522
rect 19516 6458 19572 6470
rect 19740 6468 19796 7420
rect 19852 6692 19908 7644
rect 20300 7588 20356 7980
rect 20300 7494 20356 7532
rect 19852 6626 19908 6636
rect 20076 6690 20132 6702
rect 20076 6638 20078 6690
rect 20130 6638 20132 6690
rect 19068 6244 19124 6300
rect 19628 6412 19796 6468
rect 20076 6468 20132 6638
rect 20300 6692 20356 6702
rect 20300 6598 20356 6636
rect 20412 6580 20468 8092
rect 20524 8036 20580 8046
rect 20524 7942 20580 7980
rect 20636 7476 20692 8988
rect 21308 9042 21364 9660
rect 22316 9492 22372 9774
rect 22764 9828 22820 11342
rect 23100 10638 23156 11900
rect 23324 11508 23380 12014
rect 23492 12070 23494 12122
rect 23546 12070 23548 12122
rect 23492 11732 23548 12070
rect 24332 12068 24388 12348
rect 24444 12290 24500 12908
rect 24444 12238 24446 12290
rect 24498 12238 24500 12290
rect 24444 12226 24500 12238
rect 24780 12740 24836 12750
rect 24612 12122 24668 12134
rect 24612 12070 24614 12122
rect 24666 12070 24668 12122
rect 24612 12068 24668 12070
rect 24332 12012 24668 12068
rect 24668 11732 24724 11742
rect 23492 11676 23828 11732
rect 23548 11508 23604 11518
rect 23324 11506 23604 11508
rect 23324 11454 23550 11506
rect 23602 11454 23604 11506
rect 23324 11452 23604 11454
rect 23548 11442 23604 11452
rect 22876 10612 22932 10622
rect 22876 10518 22932 10556
rect 23100 10586 23102 10638
rect 23154 10586 23156 10638
rect 23100 10276 23156 10586
rect 23772 10498 23828 11676
rect 24668 11060 24724 11676
rect 24444 11004 24724 11060
rect 24174 10836 24230 10846
rect 24174 10660 24230 10780
rect 24174 10608 24176 10660
rect 24228 10608 24230 10660
rect 24174 10596 24230 10608
rect 24332 10724 24388 10734
rect 24332 10610 24388 10668
rect 24332 10558 24334 10610
rect 24386 10558 24388 10610
rect 24332 10546 24388 10558
rect 24444 10612 24500 11004
rect 24444 10518 24500 10556
rect 24780 10836 24836 12684
rect 25452 12180 25508 13020
rect 25340 12178 25508 12180
rect 25340 12126 25454 12178
rect 25506 12126 25508 12178
rect 25340 12124 25508 12126
rect 25340 11620 25396 12124
rect 25452 12114 25508 12124
rect 25676 11732 25732 15092
rect 25900 13524 25956 13534
rect 25900 13430 25956 13468
rect 26572 13412 26628 13422
rect 25900 13300 25956 13310
rect 25788 12180 25844 12190
rect 25788 12086 25844 12124
rect 25340 11554 25396 11564
rect 25564 11676 25732 11732
rect 25452 11508 25508 11518
rect 25452 11414 25508 11452
rect 23772 10446 23774 10498
rect 23826 10446 23828 10498
rect 23772 10434 23828 10446
rect 23100 10210 23156 10220
rect 23660 9940 23716 9950
rect 23660 9846 23716 9884
rect 22876 9828 22932 9838
rect 22764 9826 22932 9828
rect 22764 9774 22878 9826
rect 22930 9774 22932 9826
rect 22764 9772 22932 9774
rect 22316 9426 22372 9436
rect 22876 9492 22932 9772
rect 22876 9426 22932 9436
rect 23324 9492 23380 9502
rect 21308 8990 21310 9042
rect 21362 8990 21364 9042
rect 21308 8978 21364 8990
rect 23212 8932 23268 8942
rect 22428 8930 23268 8932
rect 22428 8878 23214 8930
rect 23266 8878 23268 8930
rect 22428 8876 23268 8878
rect 22428 8596 22484 8876
rect 23212 8866 23268 8876
rect 22092 8540 22484 8596
rect 21924 8484 21980 8494
rect 21924 8390 21980 8428
rect 21588 8260 21644 8270
rect 21588 8166 21644 8204
rect 22092 8258 22148 8540
rect 23324 8484 23380 9436
rect 24780 9278 24836 10780
rect 25340 11396 25396 11406
rect 25340 10778 25396 11340
rect 25340 10726 25342 10778
rect 25394 10726 25396 10778
rect 25340 10714 25396 10726
rect 25452 10612 25508 10622
rect 25452 9940 25508 10556
rect 25564 10164 25620 11676
rect 25676 11508 25732 11518
rect 25676 10666 25732 11452
rect 25676 10614 25678 10666
rect 25730 10614 25732 10666
rect 25676 10602 25732 10614
rect 25788 11396 25844 11406
rect 25900 11396 25956 13244
rect 26124 12852 26180 12862
rect 26124 12850 26292 12852
rect 26124 12798 26126 12850
rect 26178 12798 26292 12850
rect 26124 12796 26292 12798
rect 26124 12786 26180 12796
rect 26124 12178 26180 12190
rect 26124 12126 26126 12178
rect 26178 12126 26180 12178
rect 26124 11508 26180 12126
rect 26236 12180 26292 12796
rect 26572 12516 26628 13356
rect 26684 13086 26740 16604
rect 27916 16212 27972 16222
rect 27916 16118 27972 16156
rect 27804 16100 27860 16110
rect 27804 15314 27860 16044
rect 28252 16100 28308 18396
rect 28588 17556 28644 19068
rect 29988 19122 30044 19134
rect 30488 19132 30544 19144
rect 29988 19070 29990 19122
rect 30042 19070 30044 19122
rect 29988 18788 30044 19070
rect 29988 18722 30044 18732
rect 28924 18340 28980 18350
rect 28924 18246 28980 18284
rect 30604 18004 30660 19854
rect 30772 19910 30774 19962
rect 30826 19910 30828 19962
rect 30772 19908 30828 19910
rect 30772 19842 30828 19852
rect 30828 19684 30884 19694
rect 30828 18450 30884 19628
rect 31052 19402 31108 19964
rect 31164 19460 31220 21644
rect 31276 21642 31332 21644
rect 31276 21590 31278 21642
rect 31330 21590 31332 21642
rect 31276 21578 31332 21590
rect 31276 21476 31332 21486
rect 31276 21382 31332 21420
rect 31388 21364 31444 21374
rect 31388 20746 31444 21308
rect 31388 20694 31390 20746
rect 31442 20694 31444 20746
rect 31388 20682 31444 20694
rect 31500 20074 31556 22876
rect 33068 22930 33348 22932
rect 33068 22878 33294 22930
rect 33346 22878 33348 22930
rect 33068 22876 33348 22878
rect 33068 22482 33124 22876
rect 33292 22866 33348 22876
rect 33068 22430 33070 22482
rect 33122 22430 33124 22482
rect 33068 22418 33124 22430
rect 33404 21812 33460 21822
rect 33404 21698 33460 21756
rect 33404 21646 33406 21698
rect 33458 21646 33460 21698
rect 33404 21634 33460 21646
rect 31612 21588 31668 21598
rect 31612 21494 31668 21532
rect 32956 21588 33012 21598
rect 32396 21476 32452 21486
rect 31276 20020 31332 20030
rect 31500 20022 31502 20074
rect 31554 20022 31556 20074
rect 32060 20804 32116 20814
rect 32060 20746 32116 20748
rect 32060 20694 32062 20746
rect 32114 20694 32116 20746
rect 32060 20244 32116 20694
rect 32396 20746 32452 21420
rect 32564 21474 32620 21486
rect 32564 21422 32566 21474
rect 32618 21422 32620 21474
rect 32564 21140 32620 21422
rect 32564 21074 32620 21084
rect 32956 20970 33012 21532
rect 32956 20918 32958 20970
rect 33010 20918 33012 20970
rect 32956 20906 33012 20918
rect 33068 20804 33124 20814
rect 32396 20694 32398 20746
rect 32450 20694 32452 20746
rect 32396 20682 32452 20694
rect 32956 20802 33124 20804
rect 32956 20750 33070 20802
rect 33122 20750 33124 20802
rect 32956 20748 33124 20750
rect 31500 20010 31556 20022
rect 31948 20020 32004 20030
rect 31276 19926 31332 19964
rect 31948 19926 32004 19964
rect 31612 19908 31668 19918
rect 31612 19814 31668 19852
rect 32060 19796 32116 20188
rect 32620 20634 32676 20646
rect 32620 20582 32622 20634
rect 32674 20582 32676 20634
rect 32452 19906 32508 19918
rect 32452 19854 32454 19906
rect 32506 19854 32508 19906
rect 32060 19740 32228 19796
rect 31388 19684 31444 19694
rect 31164 19404 31332 19460
rect 31052 19350 31054 19402
rect 31106 19350 31108 19402
rect 31052 19338 31108 19350
rect 31164 19236 31220 19246
rect 31164 19142 31220 19180
rect 30828 18398 30830 18450
rect 30882 18398 30884 18450
rect 30828 18386 30884 18398
rect 30604 17948 30996 18004
rect 28588 17106 28644 17500
rect 28588 17054 28590 17106
rect 28642 17054 28644 17106
rect 28588 17042 28644 17054
rect 29260 17554 29316 17566
rect 29260 17502 29262 17554
rect 29314 17502 29316 17554
rect 28924 16884 28980 16894
rect 28924 16790 28980 16828
rect 29260 16884 29316 17502
rect 30940 17444 30996 17948
rect 30604 17388 30996 17444
rect 31052 17668 31108 17678
rect 30156 17108 30212 17118
rect 29260 16818 29316 16828
rect 29596 16884 29652 16894
rect 30044 16884 30100 16894
rect 29596 16882 29876 16884
rect 29596 16830 29598 16882
rect 29650 16830 29876 16882
rect 29596 16828 29876 16830
rect 29596 16818 29652 16828
rect 29260 16660 29316 16670
rect 28812 16658 29316 16660
rect 28812 16606 29262 16658
rect 29314 16606 29316 16658
rect 28812 16604 29316 16606
rect 28252 16034 28308 16044
rect 28700 16100 28756 16110
rect 28700 16006 28756 16044
rect 28812 15372 28868 16604
rect 29260 16594 29316 16604
rect 29596 16212 29652 16222
rect 29596 16210 29764 16212
rect 29596 16158 29598 16210
rect 29650 16158 29764 16210
rect 29596 16156 29764 16158
rect 29596 16146 29652 16156
rect 29260 16098 29316 16110
rect 29260 16046 29262 16098
rect 29314 16046 29316 16098
rect 29260 15540 29316 16046
rect 29484 16054 29540 16066
rect 29484 16002 29486 16054
rect 29538 16002 29540 16054
rect 29484 15652 29540 16002
rect 29484 15586 29540 15596
rect 29260 15474 29316 15484
rect 27804 15262 27806 15314
rect 27858 15262 27860 15314
rect 27804 15250 27860 15262
rect 28588 15316 28868 15372
rect 28588 15314 28644 15316
rect 28588 15262 28590 15314
rect 28642 15262 28644 15314
rect 28588 15250 28644 15262
rect 26796 15092 26852 15102
rect 26796 14642 26852 15036
rect 26796 14590 26798 14642
rect 26850 14590 26852 14642
rect 26796 14578 26852 14590
rect 27580 14532 27636 14542
rect 27468 14530 27636 14532
rect 27468 14478 27582 14530
rect 27634 14478 27636 14530
rect 27468 14476 27636 14478
rect 26796 13746 26852 13758
rect 26796 13694 26798 13746
rect 26850 13694 26852 13746
rect 26796 13300 26852 13694
rect 26796 13234 26852 13244
rect 27468 13300 27524 14476
rect 27580 14466 27636 14476
rect 29372 14532 29428 14542
rect 29372 14438 29428 14476
rect 29708 14491 29764 16156
rect 29708 14439 29710 14491
rect 29762 14439 29764 14491
rect 29708 14427 29764 14439
rect 29820 14362 29876 16828
rect 30044 16098 30100 16828
rect 30156 16266 30212 17052
rect 30380 16996 30436 17006
rect 30380 16909 30436 16940
rect 30380 16857 30382 16909
rect 30434 16857 30436 16909
rect 30380 16845 30436 16857
rect 30156 16214 30158 16266
rect 30210 16214 30212 16266
rect 30156 16202 30212 16214
rect 30044 16046 30046 16098
rect 30098 16046 30100 16098
rect 30044 16034 30100 16046
rect 30604 15876 30660 17388
rect 31052 16660 31108 17612
rect 31164 17666 31220 17678
rect 31164 17614 31166 17666
rect 31218 17614 31220 17666
rect 31164 17220 31220 17614
rect 31164 17154 31220 17164
rect 31276 16996 31332 19404
rect 31388 19236 31444 19628
rect 31388 19170 31444 19180
rect 31724 19178 31780 19190
rect 31724 19126 31726 19178
rect 31778 19126 31780 19178
rect 31612 18450 31668 18462
rect 31612 18398 31614 18450
rect 31666 18398 31668 18450
rect 31612 17108 31668 18398
rect 31724 18338 31780 19126
rect 32172 19178 32228 19740
rect 32452 19460 32508 19854
rect 32452 19394 32508 19404
rect 32620 19348 32676 20582
rect 32956 19684 33012 20748
rect 33068 20738 33124 20748
rect 32956 19618 33012 19628
rect 33068 20356 33124 20366
rect 32620 19292 33012 19348
rect 32172 19126 32174 19178
rect 32226 19126 32228 19178
rect 32172 19114 32228 19126
rect 32844 19178 32900 19190
rect 32844 19126 32846 19178
rect 32898 19126 32900 19178
rect 32732 19066 32788 19078
rect 32732 19014 32734 19066
rect 32786 19014 32788 19066
rect 31948 18477 32004 18490
rect 31948 18452 31950 18477
rect 32002 18452 32004 18477
rect 31948 18386 32004 18396
rect 32284 18450 32340 18462
rect 32284 18398 32286 18450
rect 32338 18398 32340 18450
rect 31724 18286 31726 18338
rect 31778 18286 31780 18338
rect 31724 18274 31780 18286
rect 32284 17892 32340 18398
rect 32284 17826 32340 17836
rect 31948 17668 32004 17678
rect 32004 17638 32228 17668
rect 32004 17612 32174 17638
rect 31948 17574 32004 17612
rect 32172 17586 32174 17612
rect 32226 17586 32228 17638
rect 32172 17574 32228 17586
rect 32732 17108 32788 19014
rect 32844 18452 32900 19126
rect 32844 18386 32900 18396
rect 32956 17220 33012 19292
rect 33068 18506 33124 20300
rect 33236 20132 33292 20142
rect 33236 20038 33292 20076
rect 33516 20074 33572 23100
rect 33740 22372 33796 23660
rect 33908 23156 33964 23166
rect 33908 23062 33964 23100
rect 34076 22484 34132 23996
rect 34076 22418 34132 22428
rect 33740 22306 33796 22316
rect 33852 22370 33908 22382
rect 33852 22318 33854 22370
rect 33906 22318 33908 22370
rect 33740 21812 33796 21822
rect 33740 21252 33796 21756
rect 33852 21588 33908 22318
rect 34132 22260 34188 22270
rect 33852 21522 33908 21532
rect 33964 22258 34188 22260
rect 33964 22206 34134 22258
rect 34186 22206 34188 22258
rect 33964 22204 34188 22206
rect 33740 21196 33800 21252
rect 33516 20022 33518 20074
rect 33570 20022 33572 20074
rect 33516 20010 33572 20022
rect 33628 21028 33684 21038
rect 33628 20074 33684 20972
rect 33744 20764 33800 21196
rect 33744 20712 33746 20764
rect 33798 20712 33800 20764
rect 33964 20802 34020 22204
rect 34132 22194 34188 22204
rect 34300 22260 34356 24332
rect 34580 24050 34636 24332
rect 34580 23998 34582 24050
rect 34634 23998 34636 24050
rect 34580 23940 34636 23998
rect 34580 23874 34636 23884
rect 34748 23828 34804 24668
rect 34916 24612 34972 24668
rect 34748 23762 34804 23772
rect 34860 24610 34972 24612
rect 34860 24558 34918 24610
rect 34970 24558 34972 24610
rect 34860 24546 34972 24558
rect 34860 23716 34916 24546
rect 35420 24500 35476 25676
rect 35588 25508 35644 25518
rect 35588 25414 35644 25452
rect 35756 25172 35812 30716
rect 36764 30660 36820 32956
rect 37100 32562 37156 33740
rect 37212 32676 37268 35308
rect 37324 33796 37380 35420
rect 37324 33730 37380 33740
rect 37436 32788 37492 35868
rect 37660 35588 37716 35598
rect 37660 35494 37716 35532
rect 37884 35364 37940 35374
rect 37772 35082 37828 35094
rect 37772 35030 37774 35082
rect 37826 35030 37828 35082
rect 37660 34916 37716 34926
rect 37660 34822 37716 34860
rect 37772 34804 37828 35030
rect 37772 34738 37828 34748
rect 37884 34580 37940 35308
rect 38108 35028 38164 36428
rect 38276 36418 38332 36428
rect 38444 36148 38500 37436
rect 39116 37380 39172 37772
rect 40348 37828 40404 42028
rect 40460 42420 40516 42430
rect 40460 41410 40516 42364
rect 40460 41358 40462 41410
rect 40514 41358 40516 41410
rect 40460 41346 40516 41358
rect 40572 40964 40628 45388
rect 40684 46676 40740 46686
rect 40684 44548 40740 46620
rect 41188 46452 41244 46462
rect 40796 46450 41244 46452
rect 40796 46398 41190 46450
rect 41242 46398 41244 46450
rect 40796 46396 41244 46398
rect 40796 45890 40852 46396
rect 41188 46386 41244 46396
rect 41356 46228 41412 46844
rect 41748 46730 41804 46844
rect 41468 46676 41524 46686
rect 41468 46582 41524 46620
rect 41580 46674 41636 46686
rect 41580 46622 41582 46674
rect 41634 46622 41636 46674
rect 41748 46678 41750 46730
rect 41802 46678 41804 46730
rect 41748 46666 41804 46678
rect 41916 46674 41972 47292
rect 42364 47348 42420 47358
rect 42364 47254 42420 47292
rect 42812 46788 42868 47406
rect 42980 47348 43036 47358
rect 42980 47290 43036 47292
rect 42980 47238 42982 47290
rect 43034 47238 43036 47290
rect 42980 47226 43036 47238
rect 42364 46732 42868 46788
rect 40796 45838 40798 45890
rect 40850 45838 40852 45890
rect 40796 45826 40852 45838
rect 40908 46172 41524 46228
rect 40908 45108 40964 46172
rect 41356 46002 41412 46014
rect 41356 45950 41358 46002
rect 41410 45950 41412 46002
rect 41244 45890 41300 45902
rect 41244 45838 41246 45890
rect 41298 45838 41300 45890
rect 41244 45556 41300 45838
rect 41356 45780 41412 45950
rect 41468 45863 41524 46172
rect 41580 46004 41636 46622
rect 41916 46622 41918 46674
rect 41970 46622 41972 46674
rect 41580 45948 41860 46004
rect 41468 45811 41470 45863
rect 41522 45811 41524 45863
rect 41468 45799 41524 45811
rect 41804 45892 41860 45948
rect 41804 45798 41860 45836
rect 41356 45714 41412 45724
rect 41916 45556 41972 46622
rect 41244 45500 41972 45556
rect 42140 46676 42196 46686
rect 42140 45890 42196 46620
rect 42140 45838 42142 45890
rect 42194 45838 42196 45890
rect 42140 45668 42196 45838
rect 40908 45042 40964 45052
rect 40684 44482 40740 44492
rect 41244 44660 41300 44670
rect 41580 44660 41636 45500
rect 41784 45108 41840 45118
rect 41784 45014 41840 45052
rect 42028 44884 42084 44894
rect 41244 44324 41300 44604
rect 41244 44230 41300 44268
rect 41356 44604 41636 44660
rect 41692 44882 42084 44884
rect 41692 44830 42030 44882
rect 42082 44830 42084 44882
rect 41692 44828 42084 44830
rect 41356 43708 41412 44604
rect 41468 44436 41524 44446
rect 41468 44342 41524 44380
rect 41692 44278 41748 44828
rect 42028 44818 42084 44828
rect 41636 44266 41748 44278
rect 41636 44214 41638 44266
rect 41690 44214 41748 44266
rect 41804 44548 41860 44558
rect 41804 44322 41860 44492
rect 42140 44436 42196 45612
rect 42364 46564 42420 46732
rect 42588 46564 42644 46574
rect 42364 45444 42420 46508
rect 42364 45378 42420 45388
rect 42476 46562 42644 46564
rect 42476 46510 42590 46562
rect 42642 46510 42644 46562
rect 42476 46508 42644 46510
rect 42476 45220 42532 46508
rect 42588 46498 42644 46508
rect 42700 45892 42756 45902
rect 42700 45444 42756 45836
rect 43372 45556 43428 47966
rect 43820 48018 43876 48030
rect 43820 47966 43822 48018
rect 43874 47966 43876 48018
rect 43820 47458 43876 47966
rect 43820 47406 43822 47458
rect 43874 47406 43876 47458
rect 43820 46900 43876 47406
rect 44492 47572 44548 47582
rect 43820 46834 43876 46844
rect 44268 47236 44324 47246
rect 44268 46340 44324 47180
rect 44492 46674 44548 47516
rect 46396 47572 46452 47582
rect 46396 47478 46452 47516
rect 46732 47458 46788 47470
rect 45836 47430 45892 47442
rect 45836 47378 45838 47430
rect 45890 47378 45892 47430
rect 45724 47348 45780 47358
rect 44492 46622 44494 46674
rect 44546 46622 44548 46674
rect 44492 46610 44548 46622
rect 45276 46900 45332 46910
rect 45276 46676 45332 46844
rect 45388 46676 45444 46686
rect 45276 46674 45444 46676
rect 45276 46622 45278 46674
rect 45330 46622 45390 46674
rect 45442 46622 45444 46674
rect 45276 46620 45444 46622
rect 45276 46610 45332 46620
rect 45388 46610 45444 46620
rect 43820 46284 44324 46340
rect 43820 46114 43876 46284
rect 43820 46062 43822 46114
rect 43874 46062 43876 46114
rect 43820 46050 43876 46062
rect 45052 45890 45108 45902
rect 43576 45834 43632 45846
rect 43576 45782 43578 45834
rect 43630 45782 43632 45834
rect 43576 45668 43632 45782
rect 45052 45838 45054 45890
rect 45106 45838 45108 45890
rect 44884 45668 44940 45678
rect 43576 45602 43632 45612
rect 44604 45666 44940 45668
rect 44604 45614 44886 45666
rect 44938 45614 44940 45666
rect 44604 45612 44940 45614
rect 43260 45500 43428 45556
rect 44044 45556 44100 45566
rect 42700 45388 42980 45444
rect 42476 45154 42532 45164
rect 42364 45108 42420 45118
rect 42364 44660 42420 45052
rect 42700 45108 42756 45118
rect 42700 45014 42756 45052
rect 42532 44884 42588 44894
rect 42532 44882 42756 44884
rect 42532 44830 42534 44882
rect 42586 44830 42756 44882
rect 42532 44828 42756 44830
rect 42532 44818 42588 44828
rect 42364 44604 42588 44660
rect 42532 44546 42588 44604
rect 42532 44494 42534 44546
rect 42586 44494 42588 44546
rect 42532 44482 42588 44494
rect 42140 44370 42196 44380
rect 41804 44270 41806 44322
rect 41858 44270 41860 44322
rect 41804 44258 41860 44270
rect 41636 44212 41748 44214
rect 41636 44202 41692 44212
rect 40684 43652 41636 43708
rect 40684 42756 40740 43652
rect 41468 43568 41524 43580
rect 40796 43538 40852 43550
rect 40796 43486 40798 43538
rect 40850 43486 40852 43538
rect 40796 43204 40852 43486
rect 40964 43516 41470 43568
rect 41522 43516 41524 43568
rect 40964 43512 41524 43516
rect 40964 43370 41020 43512
rect 41468 43504 41524 43512
rect 41580 43428 41636 43652
rect 41692 43652 41748 43662
rect 41692 43594 41748 43596
rect 41692 43542 41694 43594
rect 41746 43542 41748 43594
rect 42700 43652 42756 44828
rect 42924 44548 42980 45388
rect 42812 44436 42868 44446
rect 42812 44322 42868 44380
rect 42812 44270 42814 44322
rect 42866 44270 42868 44322
rect 42812 44258 42868 44270
rect 42924 44322 42980 44492
rect 43148 45220 43204 45230
rect 43148 44324 43204 45164
rect 42924 44270 42926 44322
rect 42978 44270 42980 44322
rect 42924 44258 42980 44270
rect 43036 44322 43204 44324
rect 43036 44270 43150 44322
rect 43202 44270 43204 44322
rect 43036 44268 43204 44270
rect 43036 44100 43092 44268
rect 43148 44258 43204 44268
rect 43260 45133 43316 45500
rect 43260 45081 43262 45133
rect 43314 45081 43316 45133
rect 43260 44324 43316 45081
rect 43596 44996 43652 45006
rect 43484 44548 43540 44558
rect 43484 44454 43540 44492
rect 43260 44258 43316 44268
rect 42700 43586 42756 43596
rect 42812 44044 43092 44100
rect 41692 43530 41748 43542
rect 41972 43482 42028 43494
rect 41972 43430 41974 43482
rect 42026 43430 42028 43482
rect 41972 43428 42028 43430
rect 41580 43372 42028 43428
rect 40964 43318 40966 43370
rect 41018 43318 41020 43370
rect 40964 43306 41020 43318
rect 42252 43316 42308 43326
rect 42252 43222 42308 43260
rect 40796 43148 41636 43204
rect 40908 42756 40964 42766
rect 40684 42754 40964 42756
rect 40684 42702 40910 42754
rect 40962 42702 40964 42754
rect 40684 42700 40964 42702
rect 40908 42690 40964 42700
rect 41580 42756 41636 43148
rect 42028 42980 42084 42990
rect 42812 42980 42868 44044
rect 42924 43876 42980 43886
rect 42924 43538 42980 43820
rect 43092 43708 43148 43718
rect 43596 43708 43652 44940
rect 44044 44546 44100 45500
rect 44044 44494 44046 44546
rect 44098 44494 44100 44546
rect 44044 44482 44100 44494
rect 44492 45332 44548 45342
rect 44380 44324 44436 44334
rect 44380 44230 44436 44268
rect 43092 43706 43652 43708
rect 43092 43654 43094 43706
rect 43146 43654 43652 43706
rect 43092 43652 43652 43654
rect 43932 44100 43988 44110
rect 43092 43642 43148 43652
rect 42924 43486 42926 43538
rect 42978 43486 42980 43538
rect 42924 43474 42980 43486
rect 43708 43566 43764 43578
rect 43708 43514 43710 43566
rect 43762 43514 43764 43566
rect 43372 43316 43428 43326
rect 42028 42978 42644 42980
rect 42028 42926 42030 42978
rect 42082 42926 42644 42978
rect 42028 42924 42644 42926
rect 42028 42914 42084 42924
rect 41784 42756 41840 42766
rect 42364 42756 42420 42766
rect 41580 42754 41840 42756
rect 41580 42702 41786 42754
rect 41838 42702 41840 42754
rect 41580 42700 41840 42702
rect 40908 42532 40964 42542
rect 40908 41970 40964 42476
rect 40908 41918 40910 41970
rect 40962 41918 40964 41970
rect 40908 41906 40964 41918
rect 41580 41972 41636 42700
rect 41784 42690 41840 42700
rect 42028 42754 42420 42756
rect 42028 42702 42366 42754
rect 42418 42702 42420 42754
rect 42028 42700 42420 42702
rect 41784 42084 41840 42094
rect 41784 42026 41840 42028
rect 41784 41974 41786 42026
rect 41838 41974 41840 42026
rect 42028 42082 42084 42700
rect 42364 42690 42420 42700
rect 42588 42754 42644 42924
rect 42588 42702 42590 42754
rect 42642 42702 42644 42754
rect 42588 42690 42644 42702
rect 42700 42924 42868 42980
rect 43036 43092 43092 43102
rect 42700 42308 42756 42924
rect 42028 42030 42030 42082
rect 42082 42030 42084 42082
rect 42028 42018 42084 42030
rect 42476 42252 42756 42308
rect 42868 42756 42924 42766
rect 42868 42642 42924 42700
rect 42868 42590 42870 42642
rect 42922 42590 42924 42642
rect 41784 41962 41840 41974
rect 42476 41972 42532 42252
rect 42868 42196 42924 42590
rect 42868 42130 42924 42140
rect 42252 41970 42532 41972
rect 41580 41906 41636 41916
rect 42252 41918 42478 41970
rect 42530 41918 42532 41970
rect 42252 41916 42532 41918
rect 42252 41151 42308 41916
rect 42476 41906 42532 41916
rect 42588 41970 42644 41982
rect 42588 41918 42590 41970
rect 42642 41918 42644 41970
rect 42588 41300 42644 41918
rect 42868 41972 42924 41982
rect 42868 41878 42924 41916
rect 43036 41748 43092 43036
rect 43372 42754 43428 43260
rect 43708 42980 43764 43514
rect 43708 42914 43764 42924
rect 43932 43538 43988 44044
rect 44380 43876 44436 43886
rect 44380 43708 44436 43820
rect 44324 43652 44436 43708
rect 44324 43594 44380 43652
rect 43932 43486 43934 43538
rect 43986 43486 43988 43538
rect 43372 42702 43374 42754
rect 43426 42702 43428 42754
rect 43372 42690 43428 42702
rect 43540 42868 43596 42878
rect 43540 42698 43596 42812
rect 43540 42646 43542 42698
rect 43594 42646 43596 42698
rect 43820 42756 43876 42766
rect 43820 42662 43876 42700
rect 43540 42420 43596 42646
rect 42252 41099 42254 41151
rect 42306 41099 42308 41151
rect 42252 41087 42308 41099
rect 42364 41244 42644 41300
rect 42924 41692 43092 41748
rect 43372 42364 43596 42420
rect 43708 42642 43764 42654
rect 43708 42590 43710 42642
rect 43762 42590 43764 42642
rect 42364 41130 42420 41244
rect 42924 41188 42980 41692
rect 43092 41412 43148 41422
rect 43372 41412 43428 42364
rect 43484 42196 43540 42206
rect 43484 41970 43540 42140
rect 43484 41918 43486 41970
rect 43538 41918 43540 41970
rect 43484 41906 43540 41918
rect 43708 41972 43764 42590
rect 43932 42420 43988 43486
rect 44156 43540 44212 43550
rect 44324 43542 44326 43594
rect 44378 43542 44380 43594
rect 44324 43530 44380 43542
rect 44156 43446 44212 43484
rect 44100 42980 44156 42990
rect 44100 42886 44156 42924
rect 43932 42364 44100 42420
rect 44044 42026 44100 42364
rect 44492 42196 44548 45276
rect 44604 43594 44660 45612
rect 44884 45602 44940 45612
rect 44716 45444 44772 45454
rect 44716 43708 44772 45388
rect 44828 44490 44884 44502
rect 44828 44438 44830 44490
rect 44882 44438 44884 44490
rect 44828 44100 44884 44438
rect 44828 44034 44884 44044
rect 44940 44322 44996 44334
rect 44940 44270 44942 44322
rect 44994 44270 44996 44322
rect 44940 43988 44996 44270
rect 45052 44100 45108 45838
rect 45276 45890 45332 45902
rect 45276 45838 45278 45890
rect 45330 45838 45332 45890
rect 45276 45332 45332 45838
rect 45276 45266 45332 45276
rect 45500 45892 45556 45902
rect 45500 44548 45556 45836
rect 45612 45834 45668 45846
rect 45612 45782 45614 45834
rect 45666 45782 45668 45834
rect 45612 44558 45668 45782
rect 45724 45556 45780 47292
rect 45836 47012 45892 47378
rect 46508 47414 46564 47426
rect 46508 47362 46510 47414
rect 46562 47362 46564 47414
rect 46508 47236 46564 47362
rect 46508 47170 46564 47180
rect 46732 47406 46734 47458
rect 46786 47406 46788 47458
rect 45836 45668 45892 46956
rect 46732 46900 46788 47406
rect 47292 47458 47348 48076
rect 49308 47684 49364 48860
rect 47292 47406 47294 47458
rect 47346 47406 47348 47458
rect 47292 47394 47348 47406
rect 47964 47458 48020 47470
rect 47964 47406 47966 47458
rect 48018 47406 48020 47458
rect 47628 47236 47684 47246
rect 47628 47142 47684 47180
rect 46396 46844 46788 46900
rect 46060 46676 46116 46686
rect 45948 45892 46004 45902
rect 45948 45798 46004 45836
rect 46060 45722 46116 46620
rect 46172 46564 46228 46574
rect 46172 46470 46228 46508
rect 46284 46452 46340 46462
rect 46060 45670 46062 45722
rect 46114 45670 46116 45722
rect 45836 45612 46004 45668
rect 46060 45658 46116 45670
rect 46172 45780 46228 45790
rect 45724 45500 45892 45556
rect 45836 45162 45892 45500
rect 45724 45141 45780 45153
rect 45724 45108 45726 45141
rect 45778 45108 45780 45141
rect 45836 45110 45838 45162
rect 45890 45110 45892 45162
rect 45836 45098 45892 45110
rect 45724 45042 45780 45052
rect 45948 44996 46004 45612
rect 45836 44940 46004 44996
rect 46060 45134 46116 45146
rect 46060 45082 46062 45134
rect 46114 45082 46116 45134
rect 46060 44996 46116 45082
rect 45612 44546 45724 44558
rect 45612 44494 45670 44546
rect 45722 44494 45724 44546
rect 45612 44492 45724 44494
rect 45500 44482 45556 44492
rect 45668 44482 45724 44492
rect 45276 44324 45332 44334
rect 45276 44322 45444 44324
rect 45276 44270 45278 44322
rect 45330 44270 45444 44322
rect 45276 44268 45444 44270
rect 45276 44258 45332 44268
rect 45388 44212 45444 44268
rect 45388 44146 45444 44156
rect 45052 44044 45332 44100
rect 44940 43922 44996 43932
rect 45052 43876 45108 43886
rect 44716 43652 44996 43708
rect 44604 43542 44606 43594
rect 44658 43542 44660 43594
rect 44940 43594 44996 43652
rect 44604 43530 44660 43542
rect 44716 43566 44772 43578
rect 44716 43514 44718 43566
rect 44770 43514 44772 43566
rect 44940 43542 44942 43594
rect 44994 43542 44996 43594
rect 44940 43530 44996 43542
rect 44716 43092 44772 43514
rect 44492 42140 44660 42196
rect 43820 41972 43876 41982
rect 43708 41916 43820 41972
rect 44044 41974 44046 42026
rect 44098 41974 44100 42026
rect 44044 41962 44100 41974
rect 44268 41972 44324 41982
rect 43820 41878 43876 41916
rect 44268 41858 44324 41916
rect 44268 41806 44270 41858
rect 44322 41806 44324 41858
rect 44268 41794 44324 41806
rect 44492 41970 44548 41982
rect 44492 41918 44494 41970
rect 44546 41918 44548 41970
rect 43092 41410 43428 41412
rect 43092 41358 43094 41410
rect 43146 41358 43428 41410
rect 43092 41356 43428 41358
rect 43092 41346 43148 41356
rect 44492 41300 44548 41918
rect 44492 41234 44548 41244
rect 42364 41078 42366 41130
rect 42418 41078 42420 41130
rect 40572 40898 40628 40908
rect 41076 40964 41132 40974
rect 41524 40964 41580 40974
rect 41076 40870 41132 40908
rect 41244 40962 41580 40964
rect 41244 40910 41526 40962
rect 41578 40910 41580 40962
rect 41244 40908 41580 40910
rect 40460 40516 40516 40526
rect 40460 38612 40516 40460
rect 40796 40404 40852 40414
rect 40796 39730 40852 40348
rect 40796 39678 40798 39730
rect 40850 39678 40852 39730
rect 40796 39666 40852 39678
rect 40460 38162 40516 38556
rect 40460 38110 40462 38162
rect 40514 38110 40516 38162
rect 40460 38098 40516 38110
rect 40684 39396 40740 39406
rect 40348 37762 40404 37772
rect 40572 38052 40628 38062
rect 40404 37380 40460 37390
rect 39116 37286 39172 37324
rect 40348 37324 40404 37380
rect 40348 37286 40460 37324
rect 39732 37154 39788 37166
rect 39732 37102 39734 37154
rect 39786 37102 39788 37154
rect 38220 36092 38500 36148
rect 38556 36932 38612 36942
rect 38220 35474 38276 36092
rect 38556 35700 38612 36876
rect 39732 36932 39788 37102
rect 39732 36866 39788 36876
rect 40236 37044 40292 37054
rect 39340 36482 39396 36494
rect 39340 36430 39342 36482
rect 39394 36430 39396 36482
rect 39004 36260 39060 36270
rect 38220 35422 38222 35474
rect 38274 35422 38276 35474
rect 38220 35364 38276 35422
rect 38220 35298 38276 35308
rect 38332 35698 38612 35700
rect 38332 35646 38558 35698
rect 38610 35646 38612 35698
rect 38332 35644 38612 35646
rect 38108 34972 38276 35028
rect 37996 34916 38052 34926
rect 37996 34914 38164 34916
rect 37996 34862 37998 34914
rect 38050 34862 38164 34914
rect 37996 34860 38164 34862
rect 37996 34850 38052 34860
rect 37884 34514 37940 34524
rect 37996 34692 38052 34702
rect 37996 34244 38052 34636
rect 37996 34150 38052 34188
rect 37212 32610 37268 32620
rect 37324 32732 37492 32788
rect 38108 33570 38164 34860
rect 38108 33518 38110 33570
rect 38162 33518 38164 33570
rect 38108 32788 38164 33518
rect 37100 32510 37102 32562
rect 37154 32510 37156 32562
rect 37100 32498 37156 32510
rect 37324 31892 37380 32732
rect 38108 32722 38164 32732
rect 38220 32452 38276 34972
rect 38220 32386 38276 32396
rect 38108 32228 38164 32238
rect 37324 31836 37828 31892
rect 37324 31750 37380 31762
rect 37324 31698 37326 31750
rect 37378 31698 37380 31750
rect 37324 31220 37380 31698
rect 37324 31164 37716 31220
rect 36764 30604 37380 30660
rect 36876 30324 36932 30334
rect 35868 30210 35924 30222
rect 35868 30158 35870 30210
rect 35922 30158 35924 30210
rect 35868 29428 35924 30158
rect 35980 29652 36036 29662
rect 35980 29453 36036 29596
rect 35980 29401 35982 29453
rect 36034 29401 36036 29453
rect 35980 29389 36036 29401
rect 36876 29428 36932 30268
rect 37324 30175 37380 30604
rect 37660 30324 37716 31164
rect 37548 30268 37716 30324
rect 37324 30123 37326 30175
rect 37378 30123 37380 30175
rect 35868 28756 35924 29372
rect 35868 28690 35924 28700
rect 36036 28868 36092 28878
rect 36036 28754 36092 28812
rect 36036 28702 36038 28754
rect 36090 28702 36092 28754
rect 36036 28690 36092 28702
rect 36876 28868 36932 29372
rect 36484 28644 36540 28654
rect 36484 28550 36540 28588
rect 36876 28532 36932 28812
rect 36876 28466 36932 28476
rect 36988 29540 37044 29550
rect 36764 28420 36820 28430
rect 36148 28084 36204 28094
rect 35980 28028 36148 28084
rect 35868 26852 35924 26862
rect 35868 26758 35924 26796
rect 35868 25508 35924 25518
rect 35868 25414 35924 25452
rect 35420 24444 35588 24500
rect 35196 24332 35460 24342
rect 34972 24276 35028 24286
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 34972 24162 35028 24220
rect 34972 24110 34974 24162
rect 35026 24110 35028 24162
rect 34972 24098 35028 24110
rect 34860 23650 34916 23660
rect 35308 23938 35364 23950
rect 35308 23886 35310 23938
rect 35362 23886 35364 23938
rect 34916 23492 34972 23502
rect 34468 23380 34524 23390
rect 34468 23286 34524 23324
rect 34916 23380 34972 23436
rect 35308 23492 35364 23886
rect 35420 23940 35476 23950
rect 35420 23846 35476 23884
rect 35084 23380 35140 23390
rect 34916 23378 35028 23380
rect 34916 23326 34918 23378
rect 34970 23326 35028 23378
rect 34916 23314 35028 23326
rect 34636 22484 34692 22494
rect 34636 22342 34692 22428
rect 34300 22036 34356 22204
rect 34188 21980 34356 22036
rect 34412 22314 34468 22326
rect 34412 22262 34414 22314
rect 34466 22262 34468 22314
rect 34636 22290 34638 22342
rect 34690 22290 34692 22342
rect 34636 22278 34692 22290
rect 34860 22372 34916 22382
rect 34860 22290 34862 22316
rect 34914 22290 34916 22316
rect 34860 22278 34916 22290
rect 34972 22335 35028 23314
rect 34972 22283 34974 22335
rect 35026 22283 35028 22335
rect 35308 23380 35364 23436
rect 35308 23324 35476 23380
rect 35084 22372 35140 23324
rect 35308 23044 35364 23054
rect 35308 22950 35364 22988
rect 35420 22932 35476 23324
rect 35420 22866 35476 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35420 22372 35476 22382
rect 35084 22354 35308 22372
rect 35084 22316 35254 22354
rect 35252 22302 35254 22316
rect 35306 22302 35308 22354
rect 35252 22290 35308 22302
rect 35420 22290 35422 22316
rect 35474 22290 35476 22316
rect 34188 21140 34244 21980
rect 34412 21812 34468 22262
rect 34972 21924 35028 22283
rect 35420 22278 35476 22290
rect 34972 21858 35028 21868
rect 34412 21746 34468 21756
rect 35308 21474 35364 21486
rect 35308 21422 35310 21474
rect 35362 21422 35364 21474
rect 35308 21364 35364 21422
rect 35308 21298 35364 21308
rect 34188 21074 34244 21084
rect 34300 21252 34356 21262
rect 34300 21026 34356 21196
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 34300 20974 34302 21026
rect 34354 20974 34356 21026
rect 34300 20962 34356 20974
rect 34860 21028 34916 21038
rect 33964 20750 33966 20802
rect 34018 20750 34020 20802
rect 33964 20738 34020 20750
rect 34748 20914 34804 20926
rect 34748 20862 34750 20914
rect 34802 20862 34804 20914
rect 33744 20700 33800 20712
rect 34356 20244 34412 20254
rect 33628 20022 33630 20074
rect 33682 20022 33684 20074
rect 33628 19908 33684 20022
rect 33068 18454 33070 18506
rect 33122 18454 33124 18506
rect 33292 19852 33684 19908
rect 33852 20132 33908 20142
rect 33852 20046 33908 20076
rect 34356 20130 34412 20188
rect 34356 20078 34358 20130
rect 34410 20078 34412 20130
rect 34356 20066 34412 20078
rect 34748 20132 34804 20862
rect 34860 20787 34916 20972
rect 35532 21028 35588 24444
rect 35756 24162 35812 25116
rect 35756 24110 35758 24162
rect 35810 24110 35812 24162
rect 35756 24098 35812 24110
rect 35868 23044 35924 23054
rect 35644 22484 35700 22494
rect 35644 22342 35700 22428
rect 35644 22290 35646 22342
rect 35698 22290 35700 22342
rect 35644 22278 35700 22290
rect 35868 22314 35924 22988
rect 35868 22262 35870 22314
rect 35922 22262 35924 22314
rect 35868 21364 35924 22262
rect 35868 21298 35924 21308
rect 35532 20962 35588 20972
rect 34860 20735 34862 20787
rect 34914 20735 34916 20787
rect 34860 20723 34916 20735
rect 35196 20802 35252 20814
rect 35196 20750 35198 20802
rect 35250 20750 35252 20802
rect 35196 20580 35252 20750
rect 35420 20804 35476 20814
rect 35420 20802 35588 20804
rect 35420 20750 35422 20802
rect 35474 20750 35588 20802
rect 35420 20748 35588 20750
rect 35420 20738 35476 20748
rect 35196 20514 35252 20524
rect 34748 20066 34804 20076
rect 33852 19994 33854 20046
rect 33906 19994 33908 20046
rect 33292 18497 33348 19852
rect 33852 19796 33908 19994
rect 33516 19740 33908 19796
rect 34076 20046 34132 20058
rect 34076 19994 34078 20046
rect 34130 19994 34132 20046
rect 33516 18564 33572 19740
rect 33852 19124 33908 19134
rect 34076 19124 34132 19994
rect 34636 20018 34692 20030
rect 34636 19966 34638 20018
rect 34690 19966 34692 20018
rect 34636 19572 34692 19966
rect 34860 20018 34916 20030
rect 34860 19966 34862 20018
rect 34914 19966 34916 20018
rect 34860 19796 34916 19966
rect 35140 20020 35196 20030
rect 35140 19926 35196 19964
rect 34860 19730 34916 19740
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 34636 19506 34692 19516
rect 33068 18442 33124 18454
rect 33236 18485 33348 18497
rect 33236 18433 33238 18485
rect 33290 18433 33348 18485
rect 33460 18508 33572 18564
rect 33740 19122 34132 19124
rect 33740 19070 33854 19122
rect 33906 19070 34132 19122
rect 33740 19068 34132 19070
rect 33460 18506 33516 18508
rect 33460 18454 33462 18506
rect 33514 18454 33516 18506
rect 33460 18442 33516 18454
rect 33628 18478 33684 18490
rect 33628 18452 33630 18478
rect 33682 18452 33684 18478
rect 33236 18396 33348 18433
rect 33628 18386 33684 18396
rect 33740 17780 33796 19068
rect 33852 19058 33908 19068
rect 33908 18676 33964 18686
rect 33908 18450 33964 18620
rect 35532 18676 35588 20748
rect 35756 20580 35812 20590
rect 35756 20578 35924 20580
rect 35756 20526 35758 20578
rect 35810 20526 35924 20578
rect 35756 20524 35924 20526
rect 35756 20514 35812 20524
rect 35756 19348 35812 19358
rect 35756 19254 35812 19292
rect 35532 18610 35588 18620
rect 35868 18676 35924 20524
rect 35980 20045 36036 28028
rect 36148 27990 36204 28028
rect 36596 28084 36652 28094
rect 36764 28084 36820 28364
rect 36596 28082 36820 28084
rect 36596 28030 36598 28082
rect 36650 28030 36820 28082
rect 36596 28028 36820 28030
rect 36596 28018 36652 28028
rect 36764 27858 36820 28028
rect 36764 27806 36766 27858
rect 36818 27806 36820 27858
rect 36764 27794 36820 27806
rect 36988 27858 37044 29484
rect 37212 28644 37268 28654
rect 37212 28550 37268 28588
rect 36988 27806 36990 27858
rect 37042 27806 37044 27858
rect 36988 27412 37044 27806
rect 37324 27860 37380 30123
rect 37436 30212 37492 30222
rect 37436 30130 37438 30156
rect 37490 30130 37492 30156
rect 37436 30118 37492 30130
rect 37548 28868 37604 30268
rect 37660 30154 37716 30166
rect 37660 30102 37662 30154
rect 37714 30102 37716 30154
rect 37660 30100 37716 30102
rect 37660 30034 37716 30044
rect 37772 29428 37828 31836
rect 38108 31052 38164 32172
rect 38108 30996 38220 31052
rect 37996 30772 38052 30782
rect 37884 30324 37940 30334
rect 37884 30182 37940 30268
rect 37884 30130 37886 30182
rect 37938 30130 37940 30182
rect 37884 30118 37940 30130
rect 37436 28812 37604 28868
rect 37660 29372 37828 29428
rect 37436 28084 37492 28812
rect 37548 28644 37604 28654
rect 37548 28550 37604 28588
rect 37436 28018 37492 28028
rect 37324 27804 37492 27860
rect 37268 27636 37324 27646
rect 37268 27542 37324 27580
rect 36876 27356 37044 27412
rect 36484 26964 36540 27002
rect 36484 26898 36540 26908
rect 36876 26740 36932 27356
rect 37436 27300 37492 27804
rect 37324 27188 37380 27198
rect 37156 27132 37324 27188
rect 36988 27076 37044 27086
rect 36988 26908 37044 27020
rect 37156 27074 37212 27132
rect 37324 27122 37380 27132
rect 37156 27022 37158 27074
rect 37210 27022 37212 27074
rect 37156 27010 37212 27022
rect 37436 26908 37492 27244
rect 37660 27076 37716 29372
rect 37772 29204 37828 29214
rect 37772 28603 37828 29148
rect 37884 28756 37940 28766
rect 37884 28662 37940 28700
rect 37772 28551 37774 28603
rect 37826 28551 37828 28603
rect 37772 28539 37828 28551
rect 37884 28084 37940 28094
rect 37772 28026 37828 28038
rect 37772 27974 37774 28026
rect 37826 27974 37828 28026
rect 37772 27860 37828 27974
rect 37772 27794 37828 27804
rect 37884 27858 37940 28028
rect 37884 27806 37886 27858
rect 37938 27806 37940 27858
rect 37884 27794 37940 27806
rect 37996 27524 38052 30716
rect 38164 30322 38220 30996
rect 38164 30270 38166 30322
rect 38218 30270 38220 30322
rect 38164 30258 38220 30270
rect 38332 29876 38388 35644
rect 38556 35634 38612 35644
rect 38780 36258 39060 36260
rect 38780 36206 39006 36258
rect 39058 36206 39060 36258
rect 38780 36204 39060 36206
rect 38780 35026 38836 36204
rect 39004 36194 39060 36204
rect 39340 36260 39396 36430
rect 39676 36372 39732 36382
rect 39676 36370 39956 36372
rect 39676 36318 39678 36370
rect 39730 36318 39956 36370
rect 39676 36316 39956 36318
rect 39676 36306 39732 36316
rect 39340 36194 39396 36204
rect 39620 35924 39676 35934
rect 39620 35830 39676 35868
rect 39228 35700 39284 35710
rect 39004 35698 39284 35700
rect 39004 35646 39230 35698
rect 39282 35646 39284 35698
rect 39004 35644 39284 35646
rect 38892 35476 38948 35486
rect 38892 35382 38948 35420
rect 38780 34974 38782 35026
rect 38834 34974 38836 35026
rect 38780 34962 38836 34974
rect 38444 34916 38500 34926
rect 38444 31106 38500 34860
rect 38892 34804 38948 34814
rect 38892 34186 38948 34748
rect 39004 34468 39060 35644
rect 39228 35634 39284 35644
rect 39900 35698 39956 36316
rect 40236 35866 40292 36988
rect 40236 35814 40238 35866
rect 40290 35814 40292 35866
rect 40348 35924 40404 37286
rect 40572 37156 40628 37996
rect 40348 35858 40404 35868
rect 40460 37100 40628 37156
rect 40684 37156 40740 39340
rect 41244 39396 41300 40908
rect 41524 40898 41580 40908
rect 41692 40964 41748 40974
rect 41692 40852 41748 40908
rect 41972 40962 42028 40974
rect 41972 40910 41974 40962
rect 42026 40910 42028 40962
rect 41972 40852 42028 40910
rect 42364 40964 42420 41078
rect 42364 40898 42420 40908
rect 42588 41130 42644 41142
rect 42588 41078 42590 41130
rect 42642 41078 42644 41130
rect 41692 40796 42028 40852
rect 41524 40740 41580 40750
rect 41524 40626 41580 40684
rect 41524 40574 41526 40626
rect 41578 40574 41580 40626
rect 41524 40562 41580 40574
rect 41356 40404 41412 40414
rect 41356 40310 41412 40348
rect 41692 40180 41748 40796
rect 42588 40740 42644 41078
rect 41972 40684 42644 40740
rect 42812 41130 42868 41142
rect 42924 41132 43092 41188
rect 42812 41078 42814 41130
rect 42866 41078 42868 41130
rect 41972 40626 42028 40684
rect 41972 40574 41974 40626
rect 42026 40574 42028 40626
rect 41972 40562 42028 40574
rect 41804 40516 41860 40526
rect 42812 40516 42868 41078
rect 41804 40402 41860 40460
rect 42700 40460 42868 40516
rect 42924 40516 42980 40526
rect 41804 40350 41806 40402
rect 41858 40350 41860 40402
rect 41804 40338 41860 40350
rect 42588 40404 42644 40414
rect 42700 40404 42756 40460
rect 42644 40348 42756 40404
rect 42924 40458 42980 40460
rect 42924 40406 42926 40458
rect 42978 40406 42980 40458
rect 42924 40394 42980 40406
rect 42588 40310 42644 40348
rect 42812 40346 42868 40358
rect 42812 40294 42814 40346
rect 42866 40294 42868 40346
rect 42420 40180 42476 40190
rect 42812 40180 42868 40294
rect 41692 40124 41860 40180
rect 41244 39330 41300 39340
rect 41636 39394 41692 39406
rect 41636 39342 41638 39394
rect 41690 39342 41692 39394
rect 41636 39284 41692 39342
rect 41636 39218 41692 39228
rect 40796 38834 40852 38846
rect 40796 38782 40798 38834
rect 40850 38782 40852 38834
rect 40796 37268 40852 38782
rect 41580 38724 41636 38734
rect 41580 38722 41748 38724
rect 41580 38670 41582 38722
rect 41634 38670 41748 38722
rect 41580 38668 41748 38670
rect 41580 38658 41636 38668
rect 41692 38162 41748 38668
rect 41692 38110 41694 38162
rect 41746 38110 41748 38162
rect 41692 38098 41748 38110
rect 41244 38052 41300 38062
rect 41244 37958 41300 37996
rect 41580 38052 41636 38062
rect 41580 37983 41582 37996
rect 41634 37983 41636 37996
rect 41580 37958 41636 37983
rect 40796 37202 40852 37212
rect 41020 37492 41076 37502
rect 41020 37266 41076 37436
rect 41356 37492 41412 37502
rect 41020 37214 41022 37266
rect 41074 37214 41076 37266
rect 41020 37202 41076 37214
rect 41244 37293 41300 37305
rect 41244 37241 41246 37293
rect 41298 37241 41300 37293
rect 40236 35802 40292 35814
rect 39900 35646 39902 35698
rect 39954 35646 39956 35698
rect 39004 34412 39284 34468
rect 38556 34160 38612 34172
rect 38556 34108 38558 34160
rect 38610 34108 38612 34160
rect 38892 34134 38894 34186
rect 38946 34134 38948 34186
rect 38892 34122 38948 34134
rect 39060 34244 39116 34254
rect 39060 34186 39116 34188
rect 39060 34134 39062 34186
rect 39114 34134 39116 34186
rect 39060 34122 39116 34134
rect 38556 33684 38612 34108
rect 38556 33618 38612 33628
rect 39004 32900 39060 32910
rect 38668 32676 38724 32686
rect 38668 32002 38724 32620
rect 39004 32676 39060 32844
rect 39004 32674 39172 32676
rect 39004 32622 39006 32674
rect 39058 32622 39172 32674
rect 39004 32620 39172 32622
rect 39004 32610 39060 32620
rect 38668 31950 38670 32002
rect 38722 31950 38724 32002
rect 38668 31948 38724 31950
rect 38444 31054 38446 31106
rect 38498 31054 38500 31106
rect 38444 30324 38500 31054
rect 38444 30258 38500 30268
rect 38556 31892 38724 31948
rect 38780 32004 38836 32014
rect 38220 28644 38276 28654
rect 38220 28550 38276 28588
rect 38332 28420 38388 29820
rect 38556 29652 38612 31892
rect 38780 31780 38836 31948
rect 38668 31724 38836 31780
rect 39004 31892 39060 31902
rect 38668 30884 38724 31724
rect 38780 31220 38836 31230
rect 38780 31108 38836 31164
rect 38780 31052 38873 31108
rect 38817 31050 38873 31052
rect 38817 30998 38819 31050
rect 38871 30998 38873 31050
rect 38817 30986 38873 30998
rect 39004 31022 39060 31836
rect 39116 31556 39172 32620
rect 39228 31668 39284 34412
rect 39900 34356 39956 35646
rect 40236 35713 40292 35725
rect 40236 35661 40238 35713
rect 40290 35661 40292 35713
rect 40236 35476 40292 35661
rect 40236 35410 40292 35420
rect 40460 35252 40516 37100
rect 40684 37090 40740 37100
rect 41244 37044 41300 37241
rect 41244 36978 41300 36988
rect 41020 36260 41076 36270
rect 40572 36036 40628 36046
rect 40572 35364 40628 35980
rect 41020 35866 41076 36204
rect 41356 35924 41412 37436
rect 41692 37434 41748 37446
rect 41692 37382 41694 37434
rect 41746 37382 41748 37434
rect 41580 37268 41636 37278
rect 41020 35814 41022 35866
rect 41074 35814 41076 35866
rect 41020 35802 41076 35814
rect 41132 35868 41412 35924
rect 41468 37266 41636 37268
rect 41468 37214 41582 37266
rect 41634 37214 41636 37266
rect 41468 37212 41636 37214
rect 41020 35700 41076 35710
rect 41132 35700 41188 35868
rect 41468 35812 41524 37212
rect 41580 37202 41636 37212
rect 41580 36482 41636 36494
rect 41580 36430 41582 36482
rect 41634 36430 41636 36482
rect 41580 35924 41636 36430
rect 41580 35858 41636 35868
rect 41468 35746 41524 35756
rect 41020 35698 41188 35700
rect 41020 35646 41022 35698
rect 41074 35646 41188 35698
rect 41020 35644 41188 35646
rect 41244 35725 41300 35737
rect 41244 35673 41246 35725
rect 41298 35673 41300 35725
rect 41020 35634 41076 35644
rect 41244 35476 41300 35673
rect 41692 35700 41748 37382
rect 41804 37380 41860 40124
rect 42420 40178 42868 40180
rect 42420 40126 42422 40178
rect 42474 40126 42868 40178
rect 42420 40124 42868 40126
rect 42420 40114 42476 40124
rect 42532 39732 42588 39742
rect 42084 39394 42140 39406
rect 42084 39342 42086 39394
rect 42138 39342 42140 39394
rect 42084 39060 42140 39342
rect 42532 39396 42588 39676
rect 42812 39618 42868 40124
rect 42812 39566 42814 39618
rect 42866 39566 42868 39618
rect 42812 39554 42868 39566
rect 43036 39450 43092 41132
rect 44380 41186 44436 41198
rect 44380 41134 44382 41186
rect 44434 41134 44436 41186
rect 44380 41076 44436 41134
rect 44380 41010 44436 41020
rect 43876 40964 43932 40974
rect 43876 40870 43932 40908
rect 44212 40962 44268 40974
rect 44212 40910 44214 40962
rect 44266 40910 44268 40962
rect 44212 40516 44268 40910
rect 44212 40458 44268 40460
rect 43372 40404 43428 40414
rect 43036 39398 43038 39450
rect 43090 39398 43092 39450
rect 43036 39386 43092 39398
rect 43260 39562 43316 39574
rect 43260 39510 43262 39562
rect 43314 39510 43316 39562
rect 42532 39302 42588 39340
rect 43260 39172 43316 39510
rect 43260 39106 43316 39116
rect 42084 38994 42140 39004
rect 43372 38724 43428 40348
rect 43652 40404 43708 40414
rect 43988 40404 44044 40414
rect 43652 40402 44044 40404
rect 43652 40350 43654 40402
rect 43706 40350 43990 40402
rect 44042 40350 44044 40402
rect 44212 40406 44214 40458
rect 44266 40406 44268 40458
rect 44212 40394 44268 40406
rect 44492 40430 44548 40442
rect 44492 40404 44494 40430
rect 44546 40404 44548 40430
rect 43652 40348 44044 40350
rect 43652 40338 43708 40348
rect 43988 40338 44044 40348
rect 44492 40338 44548 40348
rect 43484 40290 43540 40302
rect 43484 40238 43486 40290
rect 43538 40238 43540 40290
rect 43484 39844 43540 40238
rect 44604 40180 44660 42140
rect 44716 41970 44772 43036
rect 45052 42756 45108 43820
rect 45164 43652 45220 43662
rect 45164 43594 45220 43596
rect 45164 43542 45166 43594
rect 45218 43542 45220 43594
rect 45164 43530 45220 43542
rect 45164 42756 45220 42766
rect 45052 42754 45220 42756
rect 45052 42702 45166 42754
rect 45218 42702 45220 42754
rect 45052 42700 45220 42702
rect 45164 42690 45220 42700
rect 44716 41918 44718 41970
rect 44770 41918 44772 41970
rect 44716 41906 44772 41918
rect 45164 41972 45220 41982
rect 45276 41972 45332 44044
rect 45724 43538 45780 43550
rect 45724 43486 45726 43538
rect 45778 43486 45780 43538
rect 45444 43316 45500 43326
rect 45724 43316 45780 43486
rect 45444 43314 45780 43316
rect 45444 43262 45446 43314
rect 45498 43262 45780 43314
rect 45444 43260 45780 43262
rect 45444 43250 45500 43260
rect 45388 42868 45444 42878
rect 45388 42715 45444 42812
rect 45388 42663 45390 42715
rect 45442 42663 45444 42715
rect 45724 42754 45780 43260
rect 45724 42702 45726 42754
rect 45778 42702 45780 42754
rect 45724 42690 45780 42702
rect 45388 42651 45444 42663
rect 45612 42586 45668 42598
rect 45612 42534 45614 42586
rect 45666 42534 45668 42586
rect 45276 41916 45556 41972
rect 45164 41878 45220 41916
rect 44884 41748 44940 41758
rect 45332 41748 45388 41758
rect 44884 41746 45220 41748
rect 44884 41694 44886 41746
rect 44938 41694 45220 41746
rect 44884 41692 45220 41694
rect 44884 41682 44940 41692
rect 44940 41524 44996 41534
rect 44940 41186 44996 41468
rect 44940 41134 44942 41186
rect 44994 41134 44996 41186
rect 44940 41122 44996 41134
rect 45164 41186 45220 41692
rect 45332 41746 45444 41748
rect 45332 41694 45334 41746
rect 45386 41694 45444 41746
rect 45332 41682 45444 41694
rect 45164 41134 45166 41186
rect 45218 41134 45220 41186
rect 45164 41122 45220 41134
rect 45052 40516 45108 40526
rect 45108 40460 45145 40516
rect 45052 40458 45145 40460
rect 45052 40450 45091 40458
rect 43484 39778 43540 39788
rect 44492 40124 44660 40180
rect 44716 40430 44772 40442
rect 44716 40378 44718 40430
rect 44770 40378 44772 40430
rect 44492 39732 44548 40124
rect 43484 39620 43540 39630
rect 43484 39618 43876 39620
rect 43484 39566 43486 39618
rect 43538 39566 43876 39618
rect 43484 39564 43876 39566
rect 43484 39554 43540 39564
rect 43484 38724 43540 38734
rect 43372 38722 43652 38724
rect 43372 38670 43486 38722
rect 43538 38670 43652 38722
rect 43372 38668 43652 38670
rect 43484 38658 43540 38668
rect 42495 38164 42551 38174
rect 42252 38052 42308 38062
rect 42252 37958 42308 37996
rect 42495 38050 42551 38108
rect 42495 37998 42497 38050
rect 42549 37998 42551 38050
rect 42495 37986 42551 37998
rect 43372 38052 43428 38062
rect 43596 38052 43652 38668
rect 43708 38164 43764 38174
rect 43708 38070 43764 38108
rect 43372 38050 43652 38052
rect 43372 37998 43374 38050
rect 43426 37998 43652 38050
rect 43372 37996 43652 37998
rect 43820 38006 43876 39564
rect 44324 39396 44380 39406
rect 44324 39394 44436 39396
rect 44324 39342 44326 39394
rect 44378 39342 44436 39394
rect 44324 39330 44436 39342
rect 44156 39172 44212 39182
rect 43372 37986 43428 37996
rect 43820 37954 43822 38006
rect 43874 37954 43876 38006
rect 43820 37828 43876 37954
rect 43820 37762 43876 37772
rect 44044 38276 44100 38286
rect 44044 37940 44100 38220
rect 44156 38052 44212 39116
rect 44268 38834 44324 38846
rect 44268 38782 44270 38834
rect 44322 38782 44324 38834
rect 44268 38164 44324 38782
rect 44268 38098 44324 38108
rect 44156 37958 44212 37996
rect 41804 37314 41860 37324
rect 42364 37268 42420 37278
rect 42364 36484 42420 37212
rect 43708 36594 43764 36606
rect 43708 36542 43710 36594
rect 43762 36542 43764 36594
rect 42364 36482 42532 36484
rect 42364 36430 42366 36482
rect 42418 36461 42532 36482
rect 42418 36430 42478 36461
rect 42364 36428 42478 36430
rect 42364 36418 42420 36428
rect 42476 36409 42478 36428
rect 42530 36409 42532 36461
rect 42364 35924 42420 35934
rect 42364 35830 42420 35868
rect 42028 35700 42084 35710
rect 41692 35698 42084 35700
rect 41580 35642 41636 35654
rect 41692 35646 42030 35698
rect 42082 35646 42084 35698
rect 41692 35644 42084 35646
rect 42476 35700 42532 36409
rect 42700 35700 42756 35710
rect 42476 35698 42756 35700
rect 42476 35646 42702 35698
rect 42754 35646 42756 35698
rect 42476 35644 42756 35646
rect 41580 35590 41582 35642
rect 41634 35590 41636 35642
rect 42028 35634 42084 35644
rect 42700 35634 42756 35644
rect 43484 35700 43540 35710
rect 43708 35700 43764 36542
rect 43820 36484 43876 36494
rect 43820 36415 43822 36428
rect 43874 36415 43876 36428
rect 43820 36390 43876 36415
rect 44044 36482 44100 37884
rect 44268 37380 44324 37390
rect 44268 37293 44324 37324
rect 44268 37241 44270 37293
rect 44322 37241 44324 37293
rect 44268 37229 44324 37241
rect 44380 36932 44436 39330
rect 44492 38836 44548 39676
rect 44604 39396 44660 39406
rect 44604 39002 44660 39340
rect 44604 38950 44606 39002
rect 44658 38950 44660 39002
rect 44604 38938 44660 38950
rect 44492 38770 44548 38780
rect 44604 38861 44660 38873
rect 44604 38809 44606 38861
rect 44658 38809 44660 38861
rect 44604 38500 44660 38809
rect 44604 38434 44660 38444
rect 44716 38388 44772 40378
rect 44884 40418 44940 40430
rect 44884 40366 44886 40418
rect 44938 40366 44940 40418
rect 45089 40406 45091 40450
rect 45143 40406 45145 40458
rect 45089 40394 45145 40406
rect 45276 40430 45332 40442
rect 45276 40404 45278 40430
rect 45330 40404 45332 40430
rect 44884 39842 44940 40366
rect 45276 40338 45332 40348
rect 44884 39790 44886 39842
rect 44938 39790 44940 39842
rect 44884 39172 44940 39790
rect 45388 39732 45444 41682
rect 45500 41524 45556 41916
rect 45500 41458 45556 41468
rect 45500 41300 45556 41310
rect 45500 40458 45556 41244
rect 45500 40406 45502 40458
rect 45554 40406 45556 40458
rect 45500 40394 45556 40406
rect 45612 40292 45668 42534
rect 45836 41997 45892 44940
rect 46060 44930 46116 44940
rect 46172 44772 46228 45724
rect 46284 45162 46340 46396
rect 46396 46116 46452 46844
rect 47964 46564 48020 47406
rect 49308 47458 49364 47628
rect 49308 47406 49310 47458
rect 49362 47406 49364 47458
rect 49308 47394 49364 47406
rect 48132 47236 48188 47246
rect 48132 47234 48356 47236
rect 48132 47182 48134 47234
rect 48186 47182 48356 47234
rect 48132 47180 48356 47182
rect 48132 47170 48188 47180
rect 48076 46564 48132 46574
rect 47964 46562 48132 46564
rect 47964 46510 48078 46562
rect 48130 46510 48132 46562
rect 47964 46508 48132 46510
rect 48076 46452 48132 46508
rect 48076 46386 48132 46396
rect 46396 46060 46788 46116
rect 46284 45110 46286 45162
rect 46338 45110 46340 45162
rect 46284 45098 46340 45110
rect 46396 45890 46452 45902
rect 46396 45838 46398 45890
rect 46450 45838 46452 45890
rect 46396 44772 46452 45838
rect 46564 44884 46620 44894
rect 46564 44882 46676 44884
rect 46564 44830 46566 44882
rect 46618 44830 46676 44882
rect 46564 44818 46676 44830
rect 45948 44716 46228 44772
rect 45948 44322 46004 44716
rect 46172 44436 46228 44716
rect 46172 44370 46228 44380
rect 46284 44716 46452 44772
rect 45948 44270 45950 44322
rect 46002 44270 46004 44322
rect 45948 44258 46004 44270
rect 46060 44322 46116 44334
rect 46060 44270 46062 44322
rect 46114 44270 46116 44322
rect 46060 44212 46116 44270
rect 46060 44146 46116 44156
rect 46284 43708 46340 44716
rect 46396 44548 46452 44558
rect 46396 44434 46452 44492
rect 46396 44382 46398 44434
rect 46450 44382 46452 44434
rect 46396 44370 46452 44382
rect 46508 44436 46564 44446
rect 46508 44307 46564 44380
rect 46508 44255 46510 44307
rect 46562 44255 46564 44307
rect 46508 44243 46564 44255
rect 46508 43876 46564 43886
rect 46620 43876 46676 44818
rect 46564 43820 46676 43876
rect 46732 44772 46788 46060
rect 47180 45890 47236 45902
rect 47180 45838 47182 45890
rect 47234 45838 47236 45890
rect 47180 45556 47236 45838
rect 47180 45490 47236 45500
rect 47292 45332 47348 45342
rect 46508 43810 46564 43820
rect 46284 43652 46452 43708
rect 45948 43540 46004 43550
rect 45948 43446 46004 43484
rect 46228 43316 46284 43326
rect 45836 41945 45838 41997
rect 45890 41945 45892 41997
rect 45836 41933 45892 41945
rect 46060 43314 46284 43316
rect 46060 43262 46230 43314
rect 46282 43262 46284 43314
rect 46060 43260 46284 43262
rect 45724 41188 45780 41198
rect 45724 41094 45780 41132
rect 45948 41186 46004 41198
rect 45948 41134 45950 41186
rect 46002 41134 46004 41186
rect 45948 41076 46004 41134
rect 45948 41010 46004 41020
rect 46060 40516 46116 43260
rect 46228 43250 46284 43260
rect 46396 42754 46452 43652
rect 46396 42702 46398 42754
rect 46450 42702 46452 42754
rect 46396 41972 46452 42702
rect 46396 41906 46452 41916
rect 46732 43540 46788 44716
rect 47180 45108 47236 45118
rect 46844 44660 46900 44670
rect 46844 44322 46900 44604
rect 46844 44270 46846 44322
rect 46898 44270 46900 44322
rect 46844 44212 46900 44270
rect 47180 44324 47236 45052
rect 47292 45106 47348 45276
rect 47516 45274 47572 45286
rect 47516 45222 47518 45274
rect 47570 45222 47572 45274
rect 47292 45054 47294 45106
rect 47346 45054 47348 45106
rect 47292 45042 47348 45054
rect 47404 45108 47460 45118
rect 47292 44324 47348 44334
rect 47180 44322 47348 44324
rect 47180 44270 47294 44322
rect 47346 44270 47348 44322
rect 47180 44268 47348 44270
rect 47292 44258 47348 44268
rect 46844 44146 46900 44156
rect 47292 43540 47348 43550
rect 46452 41188 46508 41198
rect 46452 40626 46508 41132
rect 46620 41076 46676 41086
rect 46620 40982 46676 41020
rect 46452 40574 46454 40626
rect 46506 40574 46508 40626
rect 46452 40562 46508 40574
rect 45780 40460 46116 40516
rect 45780 40458 45836 40460
rect 45780 40406 45782 40458
rect 45834 40406 45836 40458
rect 45780 40394 45836 40406
rect 46284 40404 46340 40414
rect 46284 40310 46340 40348
rect 45612 40236 45780 40292
rect 45612 39844 45668 39854
rect 45388 39676 45556 39732
rect 44884 39106 44940 39116
rect 45052 39618 45108 39630
rect 45052 39566 45054 39618
rect 45106 39566 45108 39618
rect 44828 38836 44884 38846
rect 45052 38836 45108 39566
rect 45500 39620 45556 39676
rect 45500 39554 45556 39564
rect 45612 39618 45668 39788
rect 45612 39566 45614 39618
rect 45666 39566 45668 39618
rect 45612 39554 45668 39566
rect 45724 39396 45780 40236
rect 46004 40178 46060 40190
rect 46004 40126 46006 40178
rect 46058 40126 46060 40178
rect 46004 39844 46060 40126
rect 46004 39778 46060 39788
rect 46396 39732 46452 39742
rect 46396 39638 46452 39676
rect 45948 39620 46004 39630
rect 46508 39618 46564 39630
rect 45948 39526 46004 39564
rect 46172 39562 46228 39574
rect 46172 39510 46174 39562
rect 46226 39510 46228 39562
rect 46172 39396 46228 39510
rect 45724 39340 46228 39396
rect 46508 39566 46510 39618
rect 46562 39566 46564 39618
rect 46508 39172 46564 39566
rect 45948 39116 46564 39172
rect 45836 38948 45892 38958
rect 45574 38871 45630 38883
rect 45276 38836 45332 38846
rect 45052 38780 45276 38836
rect 44828 38742 44884 38780
rect 45276 38742 45332 38780
rect 45388 38834 45444 38846
rect 45388 38782 45390 38834
rect 45442 38782 45444 38834
rect 45388 38668 45444 38782
rect 44716 38322 44772 38332
rect 45164 38612 45444 38668
rect 45574 38819 45576 38871
rect 45628 38819 45630 38871
rect 45574 38668 45630 38819
rect 45574 38612 45780 38668
rect 45164 38164 45220 38612
rect 45108 38108 45220 38164
rect 45276 38500 45332 38510
rect 44492 38052 44548 38062
rect 44716 38052 44772 38062
rect 44548 38050 44772 38052
rect 44548 37998 44718 38050
rect 44770 37998 44772 38050
rect 44548 37996 44772 37998
rect 44492 37986 44548 37996
rect 44716 37986 44772 37996
rect 44940 38052 44996 38062
rect 44940 37958 44996 37996
rect 45108 37490 45164 38108
rect 45276 37950 45332 38444
rect 45220 37938 45332 37950
rect 45220 37886 45222 37938
rect 45274 37886 45332 37938
rect 45220 37884 45332 37886
rect 45220 37874 45276 37884
rect 45108 37438 45110 37490
rect 45162 37438 45164 37490
rect 45108 37426 45164 37438
rect 44940 37268 44996 37278
rect 44996 37212 45108 37268
rect 44940 37174 44996 37212
rect 44380 36866 44436 36876
rect 44940 36650 44996 36662
rect 44940 36598 44942 36650
rect 44994 36598 44996 36650
rect 44044 36430 44046 36482
rect 44098 36430 44100 36482
rect 44044 36260 44100 36430
rect 44044 36194 44100 36204
rect 44828 36482 44884 36494
rect 44828 36430 44830 36482
rect 44882 36430 44884 36482
rect 43484 35698 43764 35700
rect 43484 35646 43486 35698
rect 43538 35646 43764 35698
rect 43484 35644 43764 35646
rect 43484 35634 43540 35644
rect 41580 35588 41636 35590
rect 41244 35410 41300 35420
rect 41356 35532 41636 35588
rect 40572 35298 40628 35308
rect 40460 35186 40516 35196
rect 40684 34916 40740 34926
rect 39900 34290 39956 34300
rect 40572 34860 40684 34916
rect 40236 34130 40292 34142
rect 40236 34078 40238 34130
rect 40290 34078 40292 34130
rect 40236 34020 40292 34078
rect 40124 33964 40236 34020
rect 39340 33906 39396 33918
rect 39340 33854 39342 33906
rect 39394 33854 39396 33906
rect 39340 33348 39396 33854
rect 39900 33906 39956 33918
rect 39900 33854 39902 33906
rect 39954 33854 39956 33906
rect 39900 33796 39956 33854
rect 39900 33730 39956 33740
rect 39676 33346 39732 33358
rect 39340 33282 39396 33292
rect 39452 33318 39508 33330
rect 39452 33266 39454 33318
rect 39506 33266 39508 33318
rect 39452 33236 39508 33266
rect 39452 32788 39508 33180
rect 39452 32722 39508 32732
rect 39676 33294 39678 33346
rect 39730 33294 39732 33346
rect 39452 32597 39508 32609
rect 39452 32545 39454 32597
rect 39506 32545 39508 32597
rect 39452 32004 39508 32545
rect 39452 31938 39508 31948
rect 39564 32590 39620 32602
rect 39564 32538 39566 32590
rect 39618 32538 39620 32590
rect 39564 31892 39620 32538
rect 39676 32228 39732 33294
rect 40012 33124 40068 33134
rect 40012 33030 40068 33068
rect 40012 32788 40068 32798
rect 40012 32618 40068 32732
rect 39844 32597 39900 32609
rect 39844 32545 39846 32597
rect 39898 32564 39900 32597
rect 40012 32566 40014 32618
rect 40066 32566 40068 32618
rect 39898 32545 39956 32564
rect 40012 32554 40068 32566
rect 39844 32508 39956 32545
rect 39900 32452 39956 32508
rect 39900 32396 40068 32452
rect 39676 32162 39732 32172
rect 39564 31826 39620 31836
rect 39900 31778 39956 31790
rect 39900 31726 39902 31778
rect 39954 31726 39956 31778
rect 39228 31612 39788 31668
rect 39116 31500 39508 31556
rect 39004 30970 39006 31022
rect 39058 30970 39060 31022
rect 39228 31108 39284 31118
rect 39228 31022 39284 31052
rect 39228 30996 39230 31022
rect 39004 30884 39060 30970
rect 38668 30828 38836 30884
rect 38668 30212 38724 30222
rect 38668 30118 38724 30156
rect 38780 29988 38836 30828
rect 38892 30828 39004 30884
rect 38892 30212 38948 30828
rect 39004 30790 39060 30828
rect 39116 30970 39230 30996
rect 39282 30970 39284 31022
rect 39452 31050 39508 31500
rect 39452 30998 39454 31050
rect 39506 30998 39508 31050
rect 39732 31106 39788 31612
rect 39732 31054 39734 31106
rect 39786 31054 39788 31106
rect 39732 31042 39788 31054
rect 39452 30986 39508 30998
rect 39116 30940 39284 30970
rect 38892 30146 38948 30156
rect 39004 30210 39060 30222
rect 39004 30158 39006 30210
rect 39058 30158 39060 30210
rect 38556 29586 38612 29596
rect 38668 29932 38836 29988
rect 38892 29988 38948 29998
rect 38556 29428 38612 29438
rect 38556 29334 38612 29372
rect 38332 28354 38388 28364
rect 38444 29258 38500 29270
rect 38444 29206 38446 29258
rect 38498 29206 38500 29258
rect 38332 28084 38388 28094
rect 38108 27897 38164 27909
rect 38108 27845 38110 27897
rect 38162 27845 38164 27897
rect 38108 27636 38164 27845
rect 38108 27570 38164 27580
rect 37660 27010 37716 27020
rect 37772 27468 38052 27524
rect 36988 26852 37156 26908
rect 36988 26740 37044 26750
rect 36876 26684 36988 26740
rect 36204 25282 36260 25294
rect 36204 25230 36206 25282
rect 36258 25230 36260 25282
rect 36204 24948 36260 25230
rect 36204 24882 36260 24892
rect 36372 23714 36428 23726
rect 36372 23662 36374 23714
rect 36426 23662 36428 23714
rect 36372 23492 36428 23662
rect 36372 23426 36428 23436
rect 36988 23380 37044 26684
rect 37100 24164 37156 26852
rect 37212 26852 37268 26862
rect 37212 26290 37268 26796
rect 37212 26238 37214 26290
rect 37266 26238 37268 26290
rect 37212 26226 37268 26238
rect 37324 26852 37492 26908
rect 37212 24948 37268 24958
rect 37212 24722 37268 24892
rect 37212 24670 37214 24722
rect 37266 24670 37268 24722
rect 37212 24658 37268 24670
rect 37100 24070 37156 24108
rect 36988 23314 37044 23324
rect 37324 23156 37380 26852
rect 37604 26850 37660 26862
rect 37604 26798 37606 26850
rect 37658 26798 37660 26850
rect 37604 26740 37660 26798
rect 37604 26674 37660 26684
rect 37436 26516 37492 26526
rect 37436 25730 37492 26460
rect 37772 26292 37828 27468
rect 38332 27310 38388 28028
rect 38444 27860 38500 29206
rect 38444 27766 38500 27804
rect 38220 27300 38276 27310
rect 38332 27298 38444 27310
rect 38332 27246 38390 27298
rect 38442 27246 38444 27298
rect 38332 27244 38444 27246
rect 37772 26226 37828 26236
rect 37884 27188 37940 27198
rect 37884 27074 37940 27132
rect 38108 27188 38164 27198
rect 37884 27022 37886 27074
rect 37938 27022 37940 27074
rect 37436 25678 37438 25730
rect 37490 25678 37492 25730
rect 37436 25666 37492 25678
rect 37772 25508 37828 25546
rect 37772 25442 37828 25452
rect 37772 25284 37828 25294
rect 37772 24162 37828 25228
rect 37772 24110 37774 24162
rect 37826 24110 37828 24162
rect 37772 24098 37828 24110
rect 37324 23090 37380 23100
rect 37436 23938 37492 23950
rect 37436 23886 37438 23938
rect 37490 23886 37492 23938
rect 36988 23044 37044 23054
rect 36148 22372 36204 22382
rect 36876 22372 36932 22382
rect 36148 22370 36932 22372
rect 36148 22318 36150 22370
rect 36202 22318 36878 22370
rect 36930 22318 36932 22370
rect 36148 22316 36932 22318
rect 36148 22306 36204 22316
rect 36876 22306 36932 22316
rect 36988 22036 37044 22988
rect 37212 23042 37268 23054
rect 37212 22990 37214 23042
rect 37266 22990 37268 23042
rect 37212 22594 37268 22990
rect 37436 23044 37492 23886
rect 37436 22978 37492 22988
rect 37212 22542 37214 22594
rect 37266 22542 37268 22594
rect 37212 22530 37268 22542
rect 37324 22932 37380 22942
rect 36988 21970 37044 21980
rect 37212 21924 37268 21934
rect 37324 21924 37380 22876
rect 37548 22370 37604 22382
rect 37548 22318 37550 22370
rect 37602 22318 37604 22370
rect 37548 22260 37604 22318
rect 37884 22372 37940 27022
rect 37996 27076 38052 27086
rect 37996 26290 38052 27020
rect 38108 27074 38164 27132
rect 38108 27022 38110 27074
rect 38162 27022 38164 27074
rect 38108 27010 38164 27022
rect 38220 26908 38276 27244
rect 38388 27234 38444 27244
rect 38668 26908 38724 29932
rect 38780 29426 38836 29438
rect 38780 29374 38782 29426
rect 38834 29374 38836 29426
rect 38780 29316 38836 29374
rect 38780 29250 38836 29260
rect 38892 28868 38948 29932
rect 38780 28812 38948 28868
rect 39004 28980 39060 30158
rect 39116 30100 39172 30940
rect 39228 30212 39284 30222
rect 39228 30118 39284 30156
rect 39900 30212 39956 31726
rect 40012 31108 40068 32396
rect 40012 31042 40068 31052
rect 39900 30146 39956 30156
rect 40012 30210 40068 30222
rect 40012 30158 40014 30210
rect 40066 30158 40068 30210
rect 39116 30034 39172 30044
rect 40012 29652 40068 30158
rect 40124 30100 40180 33964
rect 40236 33954 40292 33964
rect 40572 33348 40628 34860
rect 40684 34822 40740 34860
rect 41356 34804 41412 35532
rect 41804 35476 41860 35486
rect 41580 35364 41636 35374
rect 41076 34748 41412 34804
rect 41468 35028 41524 35038
rect 41076 34242 41132 34748
rect 41076 34190 41078 34242
rect 41130 34190 41132 34242
rect 41076 34178 41132 34190
rect 41468 34244 41524 34972
rect 41580 34692 41636 35308
rect 41692 35028 41748 35038
rect 41692 34914 41748 34972
rect 41692 34862 41694 34914
rect 41746 34862 41748 34914
rect 41692 34850 41748 34862
rect 41580 34636 41748 34692
rect 41356 34132 41412 34142
rect 41468 34132 41524 34188
rect 41356 34130 41524 34132
rect 41356 34078 41358 34130
rect 41410 34078 41524 34130
rect 41356 34076 41524 34078
rect 41580 34132 41636 34142
rect 41356 34066 41412 34076
rect 41580 34038 41636 34076
rect 40516 33292 40628 33348
rect 40908 33348 40964 33358
rect 40516 33290 40572 33292
rect 40516 33238 40518 33290
rect 40570 33238 40572 33290
rect 40516 33226 40572 33238
rect 40684 33290 40740 33302
rect 40684 33238 40686 33290
rect 40738 33238 40740 33290
rect 40908 33255 40910 33292
rect 40962 33255 40964 33292
rect 40908 33243 40964 33255
rect 40292 32564 40348 32574
rect 40292 32470 40348 32508
rect 40684 32452 40740 33238
rect 41468 33234 41524 33246
rect 41468 33182 41470 33234
rect 41522 33182 41524 33234
rect 40796 32564 40852 32574
rect 40796 32470 40852 32508
rect 41468 32564 41524 33182
rect 41692 32676 41748 34636
rect 41804 34018 41860 35420
rect 44156 35364 44212 35374
rect 43596 35252 43652 35262
rect 43596 35138 43652 35196
rect 43596 35086 43598 35138
rect 43650 35086 43652 35138
rect 43596 35074 43652 35086
rect 42140 35028 42196 35038
rect 42028 34858 42084 34870
rect 42028 34806 42030 34858
rect 42082 34806 42084 34858
rect 42028 34804 42084 34806
rect 41916 34244 41972 34254
rect 41916 34174 41972 34188
rect 41916 34122 41918 34174
rect 41970 34122 41972 34174
rect 41916 34110 41972 34122
rect 42028 34132 42084 34748
rect 42140 34746 42196 34972
rect 43260 35028 43316 35038
rect 42140 34694 42142 34746
rect 42194 34694 42196 34746
rect 42140 34682 42196 34694
rect 42252 34914 42308 34926
rect 42252 34862 42254 34914
rect 42306 34862 42308 34914
rect 42252 34356 42308 34862
rect 42588 34916 42644 34926
rect 42588 34822 42644 34860
rect 43260 34914 43316 34972
rect 43260 34862 43262 34914
rect 43314 34862 43316 34914
rect 43260 34850 43316 34862
rect 42756 34804 42812 34814
rect 42756 34746 42812 34748
rect 42756 34694 42758 34746
rect 42810 34694 42812 34746
rect 42756 34682 42812 34694
rect 43092 34356 43148 34366
rect 42252 34354 43148 34356
rect 42252 34302 43094 34354
rect 43146 34302 43148 34354
rect 42252 34300 43148 34302
rect 42140 34132 42196 34142
rect 42084 34130 42196 34132
rect 42084 34078 42142 34130
rect 42194 34078 42196 34130
rect 42084 34076 42196 34078
rect 42028 34038 42084 34076
rect 42140 34066 42196 34076
rect 41804 33966 41806 34018
rect 41858 33966 41860 34018
rect 41804 33954 41860 33966
rect 41972 33684 42028 33694
rect 41972 33570 42028 33628
rect 41972 33518 41974 33570
rect 42026 33518 42028 33570
rect 41972 33506 42028 33518
rect 41804 33346 41860 33358
rect 41804 33294 41806 33346
rect 41858 33294 41860 33346
rect 41804 32900 41860 33294
rect 41804 32834 41860 32844
rect 42028 32788 42084 32798
rect 41692 32620 41860 32676
rect 41468 32498 41524 32508
rect 40460 32396 40740 32452
rect 40460 31780 40516 32396
rect 41132 32340 41188 32350
rect 40684 32338 41188 32340
rect 40684 32286 41134 32338
rect 41186 32286 41188 32338
rect 40684 32284 41188 32286
rect 40684 31890 40740 32284
rect 41132 32274 41188 32284
rect 40684 31838 40686 31890
rect 40738 31838 40740 31890
rect 40684 31826 40740 31838
rect 40292 31724 40516 31780
rect 40292 31218 40348 31724
rect 40292 31166 40294 31218
rect 40346 31166 40348 31218
rect 40292 31154 40348 31166
rect 40460 31164 41412 31220
rect 40460 30994 40516 31164
rect 40460 30942 40462 30994
rect 40514 30942 40516 30994
rect 40460 30930 40516 30942
rect 40908 31029 40964 31041
rect 40908 30996 40910 31029
rect 40962 30996 40964 31029
rect 40908 30930 40964 30940
rect 41020 31022 41076 31034
rect 41020 30970 41022 31022
rect 41074 30970 41076 31022
rect 41020 30884 41076 30970
rect 41244 31022 41300 31034
rect 41244 30996 41246 31022
rect 41298 30996 41300 31022
rect 41356 30996 41412 31164
rect 41804 31108 41860 32620
rect 42028 32562 42084 32732
rect 42028 32510 42030 32562
rect 42082 32510 42084 32562
rect 42028 32004 42084 32510
rect 42252 32562 42308 34300
rect 43092 34290 43148 34300
rect 44156 34354 44212 35308
rect 44828 35150 44884 36430
rect 44940 36484 44996 36598
rect 44940 36418 44996 36428
rect 44828 35138 44940 35150
rect 44828 35086 44886 35138
rect 44938 35086 44940 35138
rect 44828 35084 44940 35086
rect 44884 35074 44940 35084
rect 44324 34692 44380 34702
rect 44324 34690 44436 34692
rect 44324 34638 44326 34690
rect 44378 34638 44436 34690
rect 44324 34626 44436 34638
rect 44156 34302 44158 34354
rect 44210 34302 44212 34354
rect 44156 34290 44212 34302
rect 42476 34130 42532 34142
rect 42476 34078 42478 34130
rect 42530 34078 42532 34130
rect 42476 32788 42532 34078
rect 42924 34132 42980 34142
rect 42644 33908 42700 33918
rect 42644 33906 42756 33908
rect 42644 33854 42646 33906
rect 42698 33854 42756 33906
rect 42644 33842 42756 33854
rect 42588 33684 42644 33694
rect 42588 33311 42644 33628
rect 42588 33259 42590 33311
rect 42642 33259 42644 33311
rect 42700 33348 42756 33842
rect 42924 33684 42980 34076
rect 43652 34132 43708 34142
rect 43652 34038 43708 34076
rect 43820 34130 43876 34142
rect 43820 34078 43822 34130
rect 43874 34078 43876 34130
rect 42924 33618 42980 33628
rect 43148 33460 43204 33470
rect 42700 33311 42812 33348
rect 42700 33292 42758 33311
rect 42588 33247 42644 33259
rect 42756 33259 42758 33292
rect 42810 33259 42812 33311
rect 43148 33318 43204 33404
rect 43820 33460 43876 34078
rect 44380 33684 44436 34626
rect 44716 34160 44772 34172
rect 44716 34108 44718 34160
rect 44770 34108 44772 34160
rect 44380 33628 44548 33684
rect 43820 33394 43876 33404
rect 42756 33247 42812 33259
rect 42924 33290 42980 33302
rect 42924 33238 42926 33290
rect 42978 33238 42980 33290
rect 43148 33266 43150 33318
rect 43202 33266 43204 33318
rect 43148 33254 43204 33266
rect 44044 33346 44100 33358
rect 44044 33294 44046 33346
rect 44098 33294 44100 33346
rect 42924 33236 42980 33238
rect 43428 33236 43484 33246
rect 42924 33170 42980 33180
rect 43260 33234 43484 33236
rect 43260 33182 43430 33234
rect 43482 33182 43484 33234
rect 43260 33180 43484 33182
rect 43260 32788 43316 33180
rect 43428 33170 43484 33180
rect 43876 33236 43932 33246
rect 43876 33178 43932 33180
rect 43876 33126 43878 33178
rect 43930 33126 43932 33178
rect 43876 33114 43932 33126
rect 42476 32722 42532 32732
rect 42998 32732 43316 32788
rect 44044 32788 44100 33294
rect 44492 33124 44548 33628
rect 44492 33058 44548 33068
rect 44044 32732 44436 32788
rect 42998 32600 43054 32732
rect 42700 32564 42756 32574
rect 42252 32510 42254 32562
rect 42306 32510 42308 32562
rect 42252 32498 42308 32510
rect 42364 32562 42756 32564
rect 42364 32510 42702 32562
rect 42754 32510 42756 32562
rect 42364 32508 42756 32510
rect 42252 32394 42308 32406
rect 42252 32342 42254 32394
rect 42306 32342 42308 32394
rect 42252 32340 42308 32342
rect 42364 32340 42420 32508
rect 42700 32498 42756 32508
rect 42812 32564 42868 32574
rect 42998 32548 43000 32600
rect 43052 32548 43054 32600
rect 42998 32536 43054 32548
rect 44268 32562 44324 32574
rect 42812 32470 42868 32508
rect 44268 32510 44270 32562
rect 44322 32510 44324 32562
rect 43372 32452 43428 32462
rect 43372 32358 43428 32396
rect 42252 32284 42420 32340
rect 42028 31938 42084 31948
rect 42588 32004 42644 32014
rect 42588 31890 42644 31948
rect 42588 31838 42590 31890
rect 42642 31838 42644 31890
rect 42588 31826 42644 31838
rect 42924 31780 42980 31790
rect 44156 31780 44212 31790
rect 42700 31778 42980 31780
rect 42700 31726 42926 31778
rect 42978 31726 42980 31778
rect 42700 31724 42980 31726
rect 42252 31108 42308 31118
rect 41804 31052 42084 31108
rect 41506 31010 41562 31022
rect 41506 30996 41508 31010
rect 41356 30958 41508 30996
rect 41560 30996 41562 31010
rect 41560 30958 41972 30996
rect 41356 30940 41972 30958
rect 41244 30930 41300 30940
rect 41020 30818 41076 30828
rect 41748 30772 41804 30782
rect 40124 30034 40180 30044
rect 41132 30770 41804 30772
rect 41132 30718 41750 30770
rect 41802 30718 41804 30770
rect 41132 30716 41804 30718
rect 41132 29988 41188 30716
rect 41748 30706 41804 30716
rect 41916 30322 41972 30940
rect 41916 30270 41918 30322
rect 41970 30270 41972 30322
rect 41916 30258 41972 30270
rect 40460 29932 41188 29988
rect 41356 30212 41412 30222
rect 40124 29652 40180 29662
rect 40012 29650 40180 29652
rect 40012 29598 40126 29650
rect 40178 29598 40180 29650
rect 40012 29596 40180 29598
rect 40124 29586 40180 29596
rect 39452 29426 39508 29438
rect 39452 29374 39454 29426
rect 39506 29374 39508 29426
rect 39284 29204 39340 29214
rect 39284 29110 39340 29148
rect 39452 29204 39508 29374
rect 40460 29426 40516 29932
rect 40460 29374 40462 29426
rect 40514 29374 40516 29426
rect 40460 29362 40516 29374
rect 41076 29428 41132 29438
rect 41076 29334 41132 29372
rect 39452 29138 39508 29148
rect 41020 29204 41076 29214
rect 38780 27188 38836 28812
rect 38892 28644 38948 28654
rect 38892 27858 38948 28588
rect 39004 28308 39060 28924
rect 40796 28644 40852 28654
rect 40796 28550 40852 28588
rect 39004 28242 39060 28252
rect 40236 28420 40292 28430
rect 40236 28082 40292 28364
rect 40236 28030 40238 28082
rect 40290 28030 40292 28082
rect 40236 28018 40292 28030
rect 41020 28094 41076 29148
rect 41356 28644 41412 30156
rect 42028 30100 42084 31052
rect 42252 31014 42308 31052
rect 42588 30996 42644 31006
rect 42700 30996 42756 31724
rect 42924 31714 42980 31724
rect 43932 31778 44212 31780
rect 43932 31726 44158 31778
rect 44210 31726 44212 31778
rect 43932 31724 44212 31726
rect 43260 31556 43316 31566
rect 43820 31556 43876 31566
rect 43260 31554 43540 31556
rect 43260 31502 43262 31554
rect 43314 31502 43540 31554
rect 43260 31500 43540 31502
rect 43260 31490 43316 31500
rect 42476 30994 42756 30996
rect 42476 30942 42590 30994
rect 42642 30942 42756 30994
rect 42476 30940 42756 30942
rect 42812 30994 42868 31006
rect 42812 30942 42814 30994
rect 42866 30942 42868 30994
rect 42252 30212 42308 30222
rect 41804 30044 42084 30100
rect 42140 30210 42308 30212
rect 42140 30158 42254 30210
rect 42306 30158 42308 30210
rect 42140 30156 42308 30158
rect 41468 29652 41524 29662
rect 41468 29453 41524 29596
rect 41468 29401 41470 29453
rect 41522 29401 41524 29453
rect 41468 29389 41524 29401
rect 41580 28644 41636 28654
rect 41356 28642 41636 28644
rect 41356 28590 41582 28642
rect 41634 28590 41636 28642
rect 41356 28588 41636 28590
rect 41020 28084 41132 28094
rect 41020 28028 41076 28084
rect 41076 27990 41132 28028
rect 39150 27972 39206 27982
rect 39150 27896 39206 27916
rect 38892 27806 38894 27858
rect 38946 27806 38948 27858
rect 38892 27794 38948 27806
rect 39004 27860 39060 27870
rect 39150 27844 39152 27896
rect 39204 27844 39206 27896
rect 39900 27860 39956 27870
rect 39150 27832 39206 27844
rect 39676 27858 39956 27860
rect 39004 27766 39060 27804
rect 39676 27806 39902 27858
rect 39954 27806 39956 27858
rect 39676 27804 39956 27806
rect 39564 27636 39620 27646
rect 38780 27122 38836 27132
rect 39116 27634 39620 27636
rect 39116 27582 39566 27634
rect 39618 27582 39620 27634
rect 39116 27580 39620 27582
rect 39004 27074 39060 27086
rect 39004 27022 39006 27074
rect 39058 27022 39060 27074
rect 39004 26964 39060 27022
rect 39116 27074 39172 27580
rect 39564 27570 39620 27580
rect 39676 27412 39732 27804
rect 39900 27794 39956 27804
rect 41356 27860 41412 28588
rect 41580 28578 41636 28588
rect 39396 27356 39732 27412
rect 39396 27298 39452 27356
rect 39396 27246 39398 27298
rect 39450 27246 39452 27298
rect 39396 27234 39452 27246
rect 40796 27188 40852 27198
rect 40796 27094 40852 27132
rect 39116 27022 39118 27074
rect 39170 27022 39172 27074
rect 39116 27010 39172 27022
rect 39676 27074 39732 27086
rect 39676 27022 39678 27074
rect 39730 27022 39732 27074
rect 39676 26908 39732 27022
rect 40460 27074 40516 27086
rect 40460 27022 40462 27074
rect 40514 27022 40516 27074
rect 40460 26908 40516 27022
rect 41132 27076 41188 27086
rect 41356 27076 41412 27804
rect 41188 27020 41412 27076
rect 41132 26982 41188 27020
rect 41804 26908 41860 30044
rect 42028 29652 42084 29662
rect 41916 28868 41972 28878
rect 41916 28642 41972 28812
rect 41916 28590 41918 28642
rect 41970 28590 41972 28642
rect 41916 28578 41972 28590
rect 41916 27188 41972 27198
rect 41916 27094 41972 27132
rect 38220 26852 38444 26908
rect 38668 26852 38836 26908
rect 37996 26238 37998 26290
rect 38050 26238 38052 26290
rect 37996 26226 38052 26238
rect 38108 26628 38164 26638
rect 38108 25471 38164 26572
rect 38388 26514 38444 26852
rect 38388 26462 38390 26514
rect 38442 26462 38444 26514
rect 38388 26450 38444 26462
rect 38780 26516 38836 26852
rect 38780 26450 38836 26460
rect 38780 26066 38836 26078
rect 38780 26014 38782 26066
rect 38834 26014 38836 26066
rect 38780 25732 38836 26014
rect 39004 25956 39060 26908
rect 39564 26852 39732 26908
rect 39340 26516 39396 26526
rect 39116 26404 39172 26414
rect 39116 26346 39172 26348
rect 39116 26294 39118 26346
rect 39170 26294 39172 26346
rect 39116 26282 39172 26294
rect 39340 26346 39396 26460
rect 39340 26294 39342 26346
rect 39394 26294 39396 26346
rect 39340 26282 39396 26294
rect 39452 26318 39508 26330
rect 39452 26292 39454 26318
rect 39506 26292 39508 26318
rect 39452 26226 39508 26236
rect 39004 25900 39172 25956
rect 38108 25419 38110 25471
rect 38162 25419 38164 25471
rect 38108 25284 38164 25419
rect 38108 25218 38164 25228
rect 38220 25676 38836 25732
rect 38948 25732 39004 25742
rect 38220 25450 38276 25676
rect 38948 25638 39004 25676
rect 38668 25508 38724 25518
rect 38220 25398 38222 25450
rect 38274 25398 38276 25450
rect 38500 25480 38556 25483
rect 38500 25471 38612 25480
rect 38500 25419 38502 25471
rect 38554 25419 38612 25471
rect 38500 25407 38612 25419
rect 38668 25426 38670 25452
rect 38722 25426 38724 25452
rect 38668 25414 38724 25426
rect 38220 24948 38276 25398
rect 38108 24892 38276 24948
rect 38332 25284 38388 25294
rect 38556 25284 38612 25407
rect 38556 25228 38836 25284
rect 37996 24722 38052 24734
rect 37996 24670 37998 24722
rect 38050 24670 38052 24722
rect 37996 23940 38052 24670
rect 38108 24500 38164 24892
rect 38332 24768 38388 25228
rect 38500 24778 38556 24790
rect 38500 24768 38502 24778
rect 38220 24724 38276 24734
rect 38332 24726 38502 24768
rect 38554 24726 38556 24778
rect 38332 24712 38556 24726
rect 38220 24630 38276 24668
rect 38668 24610 38724 25228
rect 38780 25172 38836 25228
rect 38780 25106 38836 25116
rect 39116 24768 39172 25900
rect 39564 25732 39620 26852
rect 40012 26850 40068 26862
rect 40012 26798 40014 26850
rect 40066 26798 40068 26850
rect 39900 26404 39956 26414
rect 39900 26346 39956 26348
rect 39732 26325 39788 26337
rect 39732 26273 39734 26325
rect 39786 26292 39788 26325
rect 39900 26294 39902 26346
rect 39954 26294 39956 26346
rect 39786 26273 39844 26292
rect 39900 26282 39956 26294
rect 39732 26236 39844 26273
rect 39564 25666 39620 25676
rect 39228 25508 39284 25518
rect 39228 25506 39396 25508
rect 39228 25454 39230 25506
rect 39282 25454 39396 25506
rect 39228 25452 39396 25454
rect 39228 25442 39284 25452
rect 38668 24558 38670 24610
rect 38722 24558 38724 24610
rect 38108 24444 38276 24500
rect 38220 24052 38276 24444
rect 38556 24164 38612 24174
rect 38444 24052 38500 24062
rect 38220 23996 38444 24052
rect 37996 23156 38052 23884
rect 38108 23940 38164 23950
rect 38108 23938 38276 23940
rect 38108 23886 38110 23938
rect 38162 23886 38276 23938
rect 38444 23910 38500 23996
rect 38108 23884 38276 23886
rect 38108 23874 38164 23884
rect 37996 23154 38164 23156
rect 37996 23102 37998 23154
rect 38050 23102 38164 23154
rect 37996 23100 38164 23102
rect 37996 23090 38052 23100
rect 38108 22372 38164 23100
rect 38220 23044 38276 23884
rect 38332 23882 38388 23894
rect 38332 23830 38334 23882
rect 38386 23830 38388 23882
rect 38444 23858 38446 23910
rect 38498 23858 38500 23910
rect 38444 23846 38500 23858
rect 38332 23828 38388 23830
rect 38332 23378 38388 23772
rect 38332 23326 38334 23378
rect 38386 23326 38388 23378
rect 38332 23314 38388 23326
rect 38220 22978 38276 22988
rect 38444 23156 38500 23166
rect 38220 22372 38276 22382
rect 37884 22316 38052 22372
rect 37548 22194 37604 22204
rect 37884 22148 37940 22158
rect 37268 21868 37380 21924
rect 37660 22146 37940 22148
rect 37660 22094 37886 22146
rect 37938 22094 37940 22146
rect 37660 22092 37940 22094
rect 37212 21810 37268 21868
rect 37212 21758 37214 21810
rect 37266 21758 37268 21810
rect 37212 21746 37268 21758
rect 36092 21588 36148 21626
rect 36092 21522 36148 21532
rect 36204 21586 36260 21598
rect 36204 21534 36206 21586
rect 36258 21534 36260 21586
rect 35980 19993 35982 20045
rect 36034 19993 36036 20045
rect 35980 18788 36036 19993
rect 36092 21364 36148 21374
rect 36092 20020 36148 21308
rect 36204 20244 36260 21534
rect 36428 21588 36484 21598
rect 36428 20804 36484 21532
rect 37436 21588 37492 21598
rect 36540 21364 36596 21374
rect 36540 21362 36708 21364
rect 36540 21310 36542 21362
rect 36594 21310 36708 21362
rect 36540 21308 36708 21310
rect 36540 21298 36596 21308
rect 36428 20748 36596 20804
rect 36372 20580 36428 20590
rect 36372 20486 36428 20524
rect 36204 20178 36260 20188
rect 36092 19964 36260 20020
rect 35980 18722 36036 18732
rect 35868 18610 35924 18620
rect 33908 18398 33910 18450
rect 33962 18398 33964 18450
rect 33908 18386 33964 18398
rect 34524 18452 34580 18462
rect 33740 17714 33796 17724
rect 33404 17668 33460 17678
rect 32956 17164 33124 17220
rect 32732 17052 33012 17108
rect 31612 17042 31668 17052
rect 31276 16930 31332 16940
rect 31948 16996 32004 17006
rect 30940 16658 31108 16660
rect 30940 16606 31054 16658
rect 31106 16606 31108 16658
rect 30940 16604 31108 16606
rect 30784 16324 30840 16334
rect 30784 16060 30840 16268
rect 30784 16008 30786 16060
rect 30838 16008 30840 16060
rect 30784 15996 30840 16008
rect 30940 16100 30996 16604
rect 31052 16594 31108 16604
rect 30940 16006 30996 16044
rect 31724 16100 31780 16110
rect 31724 16098 31892 16100
rect 31724 16046 31726 16098
rect 31778 16046 31892 16098
rect 31724 16044 31892 16046
rect 31724 16034 31780 16044
rect 30604 15820 30772 15876
rect 30604 15652 30660 15662
rect 30492 15540 30548 15550
rect 30492 15426 30548 15484
rect 30492 15374 30494 15426
rect 30546 15374 30548 15426
rect 29820 14310 29822 14362
rect 29874 14310 29876 14362
rect 29820 14298 29876 14310
rect 29932 14756 29988 14766
rect 29932 14530 29988 14700
rect 29932 14478 29934 14530
rect 29986 14478 29988 14530
rect 27580 13636 27636 13646
rect 29484 13636 29540 13646
rect 27580 13634 27860 13636
rect 27580 13582 27582 13634
rect 27634 13582 27860 13634
rect 27580 13580 27860 13582
rect 27580 13570 27636 13580
rect 27468 13234 27524 13244
rect 27804 13188 27860 13580
rect 29484 13634 29652 13636
rect 29484 13582 29486 13634
rect 29538 13582 29652 13634
rect 29484 13580 29652 13582
rect 29484 13570 29540 13580
rect 28364 13300 28420 13310
rect 27916 13188 27972 13198
rect 27804 13186 27972 13188
rect 27804 13134 27918 13186
rect 27970 13134 27972 13186
rect 27804 13132 27972 13134
rect 27916 13122 27972 13132
rect 26684 13076 26796 13086
rect 26740 13074 26796 13076
rect 26740 13022 26742 13074
rect 26794 13022 26796 13074
rect 26740 13020 26796 13022
rect 26684 13010 26796 13020
rect 26684 12982 26740 13010
rect 28252 12964 28308 12974
rect 28252 12870 28308 12908
rect 28364 12962 28420 13244
rect 29484 13300 29540 13310
rect 28364 12910 28366 12962
rect 28418 12910 28420 12962
rect 28364 12898 28420 12910
rect 29260 12964 29316 12974
rect 29260 12794 29316 12908
rect 28364 12740 28420 12750
rect 26572 12460 26796 12516
rect 26740 12402 26796 12460
rect 26740 12350 26742 12402
rect 26794 12350 26796 12402
rect 26740 12338 26796 12350
rect 27580 12292 27636 12302
rect 27580 12198 27636 12236
rect 28364 12222 28420 12684
rect 26572 12180 26628 12190
rect 26236 12178 26628 12180
rect 26236 12126 26574 12178
rect 26626 12126 26628 12178
rect 26236 12124 26628 12126
rect 26292 11956 26348 11966
rect 26292 11862 26348 11900
rect 26572 11732 26628 12124
rect 26124 11442 26180 11452
rect 26236 11676 26628 11732
rect 26684 12180 26740 12190
rect 25788 11394 25956 11396
rect 25788 11342 25790 11394
rect 25842 11342 25956 11394
rect 25788 11340 25956 11342
rect 25564 10108 25732 10164
rect 25564 9940 25620 9950
rect 25452 9938 25620 9940
rect 25452 9886 25566 9938
rect 25618 9886 25620 9938
rect 25452 9884 25620 9886
rect 25564 9874 25620 9884
rect 24724 9266 24836 9278
rect 24724 9214 24726 9266
rect 24778 9214 24836 9266
rect 24724 9212 24836 9214
rect 24724 9202 24780 9212
rect 24108 9042 24164 9054
rect 24108 8990 24110 9042
rect 24162 8990 24164 9042
rect 24108 8932 24164 8990
rect 24108 8866 24164 8876
rect 25116 9042 25172 9054
rect 25116 8990 25118 9042
rect 25170 8990 25172 9042
rect 25116 8932 25172 8990
rect 25116 8866 25172 8876
rect 23324 8390 23380 8428
rect 23772 8818 23828 8830
rect 23772 8766 23774 8818
rect 23826 8766 23828 8818
rect 22092 8206 22094 8258
rect 22146 8206 22148 8258
rect 22092 8194 22148 8206
rect 22316 8260 22372 8270
rect 22316 8178 22318 8204
rect 22370 8178 22372 8204
rect 22316 8166 22372 8178
rect 20860 8148 20916 8158
rect 20860 7489 20916 8092
rect 20860 7437 20862 7489
rect 20914 7437 20916 7489
rect 20860 7425 20916 7437
rect 21084 7588 21140 7598
rect 21084 7474 21140 7532
rect 20636 7410 20692 7420
rect 21084 7422 21086 7474
rect 21138 7422 21140 7474
rect 21084 7410 21140 7422
rect 21756 7476 21812 7486
rect 21756 7382 21812 7420
rect 20748 7362 20804 7374
rect 20748 7310 20750 7362
rect 20802 7310 20804 7362
rect 20748 6804 20804 7310
rect 22540 7364 22596 7374
rect 22540 7362 22820 7364
rect 22540 7310 22542 7362
rect 22594 7310 22820 7362
rect 22540 7308 22820 7310
rect 22540 7298 22596 7308
rect 22764 7028 22820 7308
rect 22764 6972 23156 7028
rect 23100 6914 23156 6972
rect 23100 6862 23102 6914
rect 23154 6862 23156 6914
rect 23100 6850 23156 6862
rect 20748 6738 20804 6748
rect 21196 6690 21252 6702
rect 21196 6638 21198 6690
rect 21250 6638 21252 6690
rect 20412 6514 20468 6524
rect 20580 6580 20636 6590
rect 20580 6578 21140 6580
rect 20580 6526 20582 6578
rect 20634 6526 21140 6578
rect 20580 6524 21140 6526
rect 20580 6514 20636 6524
rect 20076 6412 20244 6468
rect 19068 6188 19460 6244
rect 18340 6132 18396 6142
rect 18340 6038 18396 6076
rect 18732 6132 18788 6142
rect 18732 6130 19348 6132
rect 18732 6078 18734 6130
rect 18786 6078 19348 6130
rect 18732 6076 19348 6078
rect 18732 6066 18788 6076
rect 19292 5933 19348 6076
rect 19068 5908 19124 5918
rect 19292 5881 19294 5933
rect 19346 5881 19348 5933
rect 19292 5869 19348 5881
rect 19404 6020 19460 6188
rect 19068 5814 19124 5852
rect 17836 5618 17892 5628
rect 19068 5684 19124 5694
rect 17500 5236 17556 5246
rect 16604 4340 16660 4350
rect 16716 4340 16772 4956
rect 16604 4338 16772 4340
rect 16604 4286 16606 4338
rect 16658 4286 16772 4338
rect 16604 4284 16772 4286
rect 16604 4274 16660 4284
rect 16492 4162 16548 4172
rect 14028 4114 14084 4126
rect 14028 4062 14030 4114
rect 14082 4062 14084 4114
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 14028 3526 14084 4062
rect 14700 4114 14756 4126
rect 14700 4062 14702 4114
rect 14754 4062 14756 4114
rect 14700 3668 14756 4062
rect 14700 3602 14756 3612
rect 14028 3474 14030 3526
rect 14082 3474 14084 3526
rect 16940 3554 16996 5068
rect 16940 3502 16942 3554
rect 16994 3502 16996 3554
rect 16940 3490 16996 3502
rect 17276 5124 17332 5134
rect 14028 3462 14084 3474
rect 1148 3444 1204 3454
rect 1148 800 1204 3388
rect 1764 3444 1820 3454
rect 1764 3330 1820 3388
rect 4732 3444 4788 3454
rect 3220 3332 3276 3342
rect 1764 3278 1766 3330
rect 1818 3278 1820 3330
rect 1764 3266 1820 3278
rect 2940 3330 3276 3332
rect 2940 3278 3222 3330
rect 3274 3278 3276 3330
rect 2940 3276 3276 3278
rect 2940 800 2996 3276
rect 3220 3266 3276 3276
rect 4732 800 4788 3388
rect 5572 3444 5628 3454
rect 5572 3386 5628 3388
rect 5572 3334 5574 3386
rect 5626 3334 5628 3386
rect 5572 3322 5628 3334
rect 6804 3332 6860 3342
rect 8596 3332 8652 3342
rect 10388 3332 10444 3342
rect 12180 3332 12236 3342
rect 6524 3330 6860 3332
rect 6524 3278 6806 3330
rect 6858 3278 6860 3330
rect 6524 3276 6860 3278
rect 6524 800 6580 3276
rect 6804 3266 6860 3276
rect 8316 3330 8652 3332
rect 8316 3278 8598 3330
rect 8650 3278 8652 3330
rect 8316 3276 8652 3278
rect 8316 800 8372 3276
rect 8596 3266 8652 3276
rect 10108 3330 10444 3332
rect 10108 3278 10390 3330
rect 10442 3278 10444 3330
rect 10108 3276 10444 3278
rect 10108 800 10164 3276
rect 10388 3266 10444 3276
rect 11900 3330 12236 3332
rect 11900 3278 12182 3330
rect 12234 3278 12236 3330
rect 11900 3276 12236 3278
rect 11900 800 11956 3276
rect 12180 3266 12236 3276
rect 13524 3332 13580 3342
rect 15596 3332 15652 3342
rect 13524 3330 13748 3332
rect 13524 3278 13526 3330
rect 13578 3278 13748 3330
rect 13524 3276 13748 3278
rect 13524 3266 13580 3276
rect 13692 800 13748 3276
rect 15484 3330 15652 3332
rect 15484 3278 15598 3330
rect 15650 3278 15652 3330
rect 15484 3276 15652 3278
rect 15484 800 15540 3276
rect 15596 3266 15652 3276
rect 17276 800 17332 5068
rect 17500 5094 17556 5180
rect 17500 5042 17502 5094
rect 17554 5042 17556 5094
rect 18508 5234 18564 5246
rect 18508 5182 18510 5234
rect 18562 5182 18564 5234
rect 18508 5124 18564 5182
rect 18508 5058 18564 5068
rect 18956 5124 19012 5134
rect 17500 5030 17556 5042
rect 18732 5012 18788 5022
rect 17724 4900 17780 4910
rect 17724 4338 17780 4844
rect 18508 4506 18564 4518
rect 18508 4454 18510 4506
rect 18562 4454 18564 4506
rect 17724 4286 17726 4338
rect 17778 4286 17780 4338
rect 17724 4274 17780 4286
rect 17948 4338 18004 4350
rect 17948 4286 17950 4338
rect 18002 4286 18004 4338
rect 17444 4228 17500 4238
rect 17444 4134 17500 4172
rect 17724 3668 17780 3678
rect 17724 3574 17780 3612
rect 17948 3668 18004 4286
rect 18396 4338 18452 4350
rect 18396 4286 18398 4338
rect 18450 4286 18452 4338
rect 18396 4228 18452 4286
rect 18508 4340 18564 4454
rect 18732 4394 18788 4956
rect 18732 4342 18734 4394
rect 18786 4342 18788 4394
rect 18732 4330 18788 4342
rect 18956 4338 19012 5068
rect 18508 4274 18564 4284
rect 18956 4286 18958 4338
rect 19010 4286 19012 4338
rect 18956 4274 19012 4286
rect 18396 4162 18452 4172
rect 17948 3602 18004 3612
rect 19068 800 19124 5628
rect 19404 5124 19460 5964
rect 19404 5058 19460 5068
rect 19628 4338 19684 6412
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 20076 6132 20132 6142
rect 20188 6132 20244 6412
rect 20132 6076 20244 6132
rect 20076 6066 20132 6076
rect 20300 5684 20356 5694
rect 20300 5590 20356 5628
rect 20188 5236 20244 5246
rect 20188 4900 20244 5180
rect 20636 5236 20692 5246
rect 20188 4834 20244 4844
rect 20300 5122 20356 5134
rect 20300 5070 20302 5122
rect 20354 5070 20356 5122
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19628 4286 19630 4338
rect 19682 4286 19684 4338
rect 19628 4274 19684 4286
rect 19628 3668 19684 3678
rect 19628 3574 19684 3612
rect 20300 3668 20356 5070
rect 20636 5107 20692 5180
rect 20636 5055 20638 5107
rect 20690 5055 20692 5107
rect 20748 5234 20804 5246
rect 20748 5182 20750 5234
rect 20802 5182 20804 5234
rect 20748 5124 20804 5182
rect 21084 5124 21140 6524
rect 21196 6468 21252 6638
rect 22428 6692 22484 6702
rect 23436 6692 23492 6702
rect 22428 6690 22596 6692
rect 22428 6638 22430 6690
rect 22482 6638 22596 6690
rect 22428 6636 22596 6638
rect 22428 6626 22484 6636
rect 21196 6402 21252 6412
rect 21532 6468 21588 6478
rect 22092 6468 22148 6478
rect 21532 6374 21588 6412
rect 21644 6466 22148 6468
rect 21644 6414 22094 6466
rect 22146 6414 22148 6466
rect 21644 6412 22148 6414
rect 21196 5124 21252 5134
rect 21084 5122 21252 5124
rect 21084 5070 21198 5122
rect 21250 5070 21252 5122
rect 21084 5068 21252 5070
rect 20748 5058 20804 5068
rect 21196 5058 21252 5068
rect 20636 5043 20692 5055
rect 21532 4900 21588 4910
rect 20412 4898 21588 4900
rect 20412 4846 21534 4898
rect 21586 4846 21588 4898
rect 20412 4844 21588 4846
rect 20412 4338 20468 4844
rect 21532 4834 21588 4844
rect 20412 4286 20414 4338
rect 20466 4286 20468 4338
rect 20412 4274 20468 4286
rect 21644 3780 21700 6412
rect 22092 6402 22148 6412
rect 22186 5908 22242 5918
rect 22428 5908 22484 5918
rect 22186 5814 22242 5852
rect 22316 5906 22484 5908
rect 22316 5854 22430 5906
rect 22482 5854 22484 5906
rect 22316 5852 22484 5854
rect 22186 5010 22242 5022
rect 22186 4958 22188 5010
rect 22240 4958 22242 5010
rect 22186 4564 22242 4958
rect 22186 4498 22242 4508
rect 22316 4450 22372 5852
rect 22428 5842 22484 5852
rect 22316 4398 22318 4450
rect 22370 4398 22372 4450
rect 22316 4386 22372 4398
rect 22428 5122 22484 5134
rect 22428 5070 22430 5122
rect 22482 5070 22484 5122
rect 21420 3724 21700 3780
rect 20300 3602 20356 3612
rect 20860 3668 20916 3678
rect 20132 3444 20188 3454
rect 20132 3386 20188 3388
rect 20132 3334 20134 3386
rect 20186 3334 20188 3386
rect 20132 3322 20188 3334
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20860 800 20916 3612
rect 21420 3526 21476 3724
rect 22092 3668 22148 3678
rect 22092 3574 22148 3612
rect 22428 3668 22484 5070
rect 22540 4564 22596 6636
rect 23436 6598 23492 6636
rect 22932 6468 22988 6478
rect 22932 5962 22988 6412
rect 22932 5910 22934 5962
rect 22986 5910 22988 5962
rect 23772 6020 23828 8766
rect 24332 8820 24388 8830
rect 23996 8148 24052 8158
rect 23884 6692 23940 6702
rect 23884 6522 23940 6636
rect 23996 6692 24052 8092
rect 24332 7364 24388 8764
rect 25452 8820 25508 8830
rect 25116 8484 25172 8494
rect 25004 8260 25060 8270
rect 24444 8258 25060 8260
rect 24444 8206 25006 8258
rect 25058 8206 25060 8258
rect 24444 8204 25060 8206
rect 24444 7586 24500 8204
rect 24444 7534 24446 7586
rect 24498 7534 24500 7586
rect 24444 7522 24500 7534
rect 24332 7308 24500 7364
rect 24332 6692 24388 6703
rect 23996 6690 24276 6692
rect 23996 6638 23998 6690
rect 24050 6638 24276 6690
rect 23996 6636 24276 6638
rect 23996 6626 24052 6636
rect 23884 6470 23886 6522
rect 23938 6470 23940 6522
rect 23884 6458 23940 6470
rect 23772 5954 23828 5964
rect 22932 5178 22988 5910
rect 22932 5126 22934 5178
rect 22986 5126 22988 5178
rect 22932 4676 22988 5126
rect 23100 5906 23156 5918
rect 23100 5854 23102 5906
rect 23154 5854 23156 5906
rect 23100 5124 23156 5854
rect 24220 5908 24276 6636
rect 24444 6692 24500 7308
rect 24556 6692 24612 6702
rect 24444 6690 24612 6692
rect 24444 6638 24558 6690
rect 24610 6638 24612 6690
rect 24444 6636 24612 6638
rect 24332 6611 24334 6636
rect 24386 6611 24388 6636
rect 24556 6626 24612 6636
rect 25004 6690 25060 8204
rect 25116 7474 25172 8428
rect 25452 8484 25508 8764
rect 25452 8418 25508 8428
rect 25228 8260 25284 8270
rect 25228 8258 25396 8260
rect 25228 8206 25230 8258
rect 25282 8206 25396 8258
rect 25228 8204 25396 8206
rect 25228 8194 25284 8204
rect 25116 7422 25118 7474
rect 25170 7422 25172 7474
rect 25116 7410 25172 7422
rect 25004 6638 25006 6690
rect 25058 6638 25060 6690
rect 25004 6626 25060 6638
rect 25340 6804 25396 8204
rect 25508 8148 25564 8158
rect 25508 8054 25564 8092
rect 25676 6916 25732 10108
rect 25788 9044 25844 11340
rect 26124 10612 26180 10622
rect 26236 10612 26292 11676
rect 26572 11394 26628 11406
rect 26572 11342 26574 11394
rect 26626 11342 26628 11394
rect 26572 10836 26628 11342
rect 26572 10770 26628 10780
rect 26124 10610 26292 10612
rect 26124 10558 26126 10610
rect 26178 10558 26292 10610
rect 26124 10556 26292 10558
rect 26348 10612 26404 10622
rect 26124 10546 26180 10556
rect 26348 10518 26404 10556
rect 26516 10500 26572 10510
rect 26516 10442 26572 10444
rect 26516 10390 26518 10442
rect 26570 10390 26572 10442
rect 26516 10378 26572 10390
rect 26012 9044 26068 9054
rect 25788 9042 26068 9044
rect 25788 8990 26014 9042
rect 26066 8990 26068 9042
rect 25788 8988 26068 8990
rect 26012 8978 26068 8988
rect 26684 8932 26740 12124
rect 27244 12180 27300 12190
rect 27244 12086 27300 12124
rect 28140 12180 28196 12190
rect 28140 12178 28308 12180
rect 28140 12126 28142 12178
rect 28194 12126 28308 12178
rect 28364 12170 28366 12222
rect 28418 12170 28420 12222
rect 28364 12158 28420 12170
rect 28812 12740 28868 12750
rect 29260 12742 29262 12794
rect 29314 12742 29316 12794
rect 29260 12730 29316 12742
rect 29372 12962 29428 12974
rect 29372 12910 29374 12962
rect 29426 12910 29428 12962
rect 29372 12740 29428 12910
rect 28140 12124 28308 12126
rect 28140 12114 28196 12124
rect 28252 11396 28308 12124
rect 28476 12066 28532 12078
rect 28476 12014 28478 12066
rect 28530 12014 28532 12066
rect 28476 11508 28532 12014
rect 28476 11442 28532 11452
rect 28252 11340 28420 11396
rect 28364 11284 28420 11340
rect 28476 11284 28532 11294
rect 28364 11282 28644 11284
rect 28364 11230 28478 11282
rect 28530 11230 28644 11282
rect 28364 11228 28644 11230
rect 28476 11218 28532 11228
rect 27804 10836 27860 10846
rect 27804 10742 27860 10780
rect 28140 10612 28196 10622
rect 28140 10518 28196 10556
rect 28588 10610 28644 11228
rect 28588 10558 28590 10610
rect 28642 10558 28644 10610
rect 28588 10546 28644 10558
rect 28812 10610 28868 12684
rect 29372 12674 29428 12684
rect 29148 12404 29204 12414
rect 29148 12205 29204 12348
rect 29148 12153 29150 12205
rect 29202 12153 29204 12205
rect 29148 12141 29204 12153
rect 29484 11956 29540 13244
rect 29596 12964 29652 13580
rect 29932 13524 29988 14478
rect 29932 13458 29988 13468
rect 30044 14532 30100 14542
rect 29596 12898 29652 12908
rect 29708 13076 29764 13086
rect 29708 12935 29764 13020
rect 29708 12883 29710 12935
rect 29762 12883 29764 12935
rect 29708 12871 29764 12883
rect 30044 12962 30100 14476
rect 30492 14530 30548 15374
rect 30492 14478 30494 14530
rect 30546 14478 30548 14530
rect 30492 14466 30548 14478
rect 30604 14530 30660 15596
rect 30604 14478 30606 14530
rect 30658 14478 30660 14530
rect 30604 14466 30660 14478
rect 30492 13524 30548 13534
rect 30380 13076 30436 13086
rect 30380 12982 30436 13020
rect 30044 12910 30046 12962
rect 30098 12910 30100 12962
rect 30044 12292 30100 12910
rect 30492 12947 30548 13468
rect 30716 13188 30772 15820
rect 31724 15652 31780 15662
rect 31388 15482 31444 15494
rect 31388 15430 31390 15482
rect 31442 15430 31444 15482
rect 31052 15314 31108 15326
rect 31052 15262 31054 15314
rect 31106 15262 31108 15314
rect 30884 14756 30940 14766
rect 30884 14662 30940 14700
rect 31052 14532 31108 15262
rect 31052 14466 31108 14476
rect 31388 14532 31444 15430
rect 31500 15353 31556 15365
rect 31500 15301 31502 15353
rect 31554 15301 31556 15353
rect 31500 14644 31556 15301
rect 31724 15314 31780 15596
rect 31724 15262 31726 15314
rect 31778 15262 31780 15314
rect 31724 15250 31780 15262
rect 31836 14868 31892 16044
rect 31948 15876 32004 16940
rect 31948 15820 32116 15876
rect 31836 14802 31892 14812
rect 31948 15316 32004 15326
rect 31612 14644 31668 14654
rect 31500 14642 31668 14644
rect 31500 14590 31614 14642
rect 31666 14590 31668 14642
rect 31500 14588 31668 14590
rect 31612 14578 31668 14588
rect 31724 14644 31780 14654
rect 31388 14466 31444 14476
rect 31724 14515 31780 14588
rect 31724 14463 31726 14515
rect 31778 14463 31780 14515
rect 31948 14530 32004 15260
rect 31948 14478 31950 14530
rect 32002 14478 32004 14530
rect 31948 14466 32004 14478
rect 31724 13748 31780 14463
rect 31388 13692 31780 13748
rect 31052 13300 31108 13310
rect 30716 13132 30884 13188
rect 30492 12895 30494 12947
rect 30546 12895 30548 12947
rect 30492 12883 30548 12895
rect 30716 12964 30772 12974
rect 30716 12870 30772 12908
rect 29820 11956 29876 11966
rect 29484 11954 29876 11956
rect 29484 11902 29822 11954
rect 29874 11902 29876 11954
rect 29484 11900 29876 11902
rect 29372 11396 29428 11406
rect 29148 11394 29428 11396
rect 29148 11342 29374 11394
rect 29426 11342 29428 11394
rect 29148 11340 29428 11342
rect 29148 10734 29204 11340
rect 29372 11330 29428 11340
rect 29092 10722 29204 10734
rect 29092 10670 29094 10722
rect 29146 10670 29204 10722
rect 29092 10658 29204 10670
rect 28812 10558 28814 10610
rect 28866 10558 28868 10610
rect 28812 10546 28868 10558
rect 28140 9938 28196 9950
rect 28140 9886 28142 9938
rect 28194 9886 28196 9938
rect 27580 9828 27636 9838
rect 27580 9826 27972 9828
rect 27580 9774 27582 9826
rect 27634 9774 27972 9826
rect 27580 9772 27972 9774
rect 27580 9762 27636 9772
rect 27244 9604 27300 9614
rect 26796 9602 27300 9604
rect 26796 9550 27246 9602
rect 27298 9550 27300 9602
rect 26796 9548 27300 9550
rect 26796 9042 26852 9548
rect 27244 9538 27300 9548
rect 26796 8990 26798 9042
rect 26850 8990 26852 9042
rect 26796 8978 26852 8990
rect 26684 8866 26740 8876
rect 27132 8484 27188 8494
rect 26572 8258 26628 8270
rect 26572 8206 26574 8258
rect 26626 8206 26628 8258
rect 26236 8036 26292 8046
rect 25900 8034 26292 8036
rect 25900 7982 26238 8034
rect 26290 7982 26292 8034
rect 25900 7980 26292 7982
rect 25900 7474 25956 7980
rect 26236 7970 26292 7980
rect 26572 7700 26628 8206
rect 26964 8260 27020 8270
rect 26964 8166 27020 8204
rect 25900 7422 25902 7474
rect 25954 7422 25956 7474
rect 25900 7410 25956 7422
rect 26124 7644 26628 7700
rect 26124 7140 26180 7644
rect 26124 7084 26404 7140
rect 25676 6860 26012 6916
rect 25340 6675 25396 6748
rect 25340 6623 25342 6675
rect 25394 6623 25396 6675
rect 25452 6802 25508 6814
rect 25452 6750 25454 6802
rect 25506 6750 25508 6802
rect 25452 6692 25508 6750
rect 25956 6692 26012 6860
rect 25452 6626 25508 6636
rect 25844 6690 26012 6692
rect 25844 6638 25958 6690
rect 26010 6638 26012 6690
rect 25844 6636 26012 6638
rect 25340 6611 25396 6623
rect 24332 6599 24388 6611
rect 25396 6468 25452 6478
rect 24556 6132 24612 6142
rect 24444 5908 24500 5918
rect 24220 5906 24500 5908
rect 24220 5854 24446 5906
rect 24498 5854 24500 5906
rect 24220 5852 24500 5854
rect 24444 5842 24500 5852
rect 24556 5906 24612 6076
rect 25396 6132 25452 6412
rect 25844 6132 25900 6636
rect 25956 6626 26012 6636
rect 26348 6522 26404 7084
rect 26460 6804 26516 6814
rect 26460 6690 26516 6748
rect 26460 6638 26462 6690
rect 26514 6638 26516 6690
rect 26460 6626 26516 6638
rect 26796 6692 26852 6702
rect 26796 6611 26798 6636
rect 26850 6611 26852 6636
rect 27132 6690 27188 8428
rect 27468 8258 27524 8270
rect 27468 8206 27470 8258
rect 27522 8206 27524 8258
rect 27468 7476 27524 8206
rect 27804 8202 27860 8214
rect 27804 8150 27806 8202
rect 27858 8150 27860 8202
rect 27804 7924 27860 8150
rect 27916 8090 27972 9772
rect 28028 9044 28084 9054
rect 28028 8484 28084 8988
rect 28028 8258 28084 8428
rect 28028 8206 28030 8258
rect 28082 8206 28084 8258
rect 28028 8194 28084 8206
rect 27916 8038 27918 8090
rect 27970 8038 27972 8090
rect 27916 8026 27972 8038
rect 28140 8036 28196 9886
rect 28252 9828 28308 9838
rect 28252 9759 28254 9772
rect 28306 9759 28308 9772
rect 28252 9734 28308 9759
rect 28588 9826 28644 9838
rect 28588 9774 28590 9826
rect 28642 9774 28644 9826
rect 28588 9156 28644 9774
rect 29148 9828 29204 10658
rect 29260 11226 29316 11238
rect 29260 11174 29262 11226
rect 29314 11174 29316 11226
rect 29260 10612 29316 11174
rect 29260 10546 29316 10556
rect 29372 10612 29428 10622
rect 29484 10612 29540 11900
rect 29820 11890 29876 11900
rect 29596 11508 29652 11518
rect 29596 11355 29652 11452
rect 29596 11303 29598 11355
rect 29650 11303 29652 11355
rect 30044 11394 30100 12236
rect 30492 11396 30548 11406
rect 30044 11342 30046 11394
rect 30098 11342 30100 11394
rect 30044 11330 30100 11342
rect 30380 11394 30548 11396
rect 30380 11342 30494 11394
rect 30546 11342 30548 11394
rect 30380 11340 30548 11342
rect 29596 11291 29652 11303
rect 29372 10610 29540 10612
rect 29372 10558 29374 10610
rect 29426 10558 29540 10610
rect 29372 10556 29540 10558
rect 28700 9156 28756 9166
rect 28588 9154 29092 9156
rect 28588 9102 28702 9154
rect 28754 9102 29092 9154
rect 28588 9100 29092 9102
rect 28700 9090 28756 9100
rect 29036 9042 29092 9100
rect 29036 8990 29038 9042
rect 29090 8990 29092 9042
rect 29036 8978 29092 8990
rect 29148 9044 29204 9772
rect 29260 9044 29316 9054
rect 29148 9042 29316 9044
rect 29148 8990 29262 9042
rect 29314 8990 29316 9042
rect 29148 8988 29316 8990
rect 29260 8978 29316 8988
rect 28028 7980 28196 8036
rect 28924 8932 28980 8942
rect 28028 7924 28084 7980
rect 27804 7868 28084 7924
rect 27804 7476 27860 7486
rect 28140 7476 28196 7486
rect 27524 7420 27636 7476
rect 27468 7410 27524 7420
rect 27132 6638 27134 6690
rect 27186 6638 27188 6690
rect 27132 6626 27188 6638
rect 27468 6802 27524 6814
rect 27468 6750 27470 6802
rect 27522 6750 27524 6802
rect 27468 6692 27524 6750
rect 27468 6626 27524 6636
rect 27580 6675 27636 7420
rect 27804 7474 28196 7476
rect 27804 7422 27806 7474
rect 27858 7422 28142 7474
rect 28194 7422 28196 7474
rect 27804 7420 28196 7422
rect 27804 7410 27860 7420
rect 27580 6623 27582 6675
rect 27634 6623 27636 6675
rect 27916 6690 27972 7420
rect 28140 7410 28196 7420
rect 28364 7476 28420 7486
rect 28364 7382 28420 7420
rect 28924 7474 28980 8876
rect 29372 8428 29428 10556
rect 30156 10498 30212 10510
rect 30156 10446 30158 10498
rect 30210 10446 30212 10498
rect 30156 10052 30212 10446
rect 30380 10276 30436 11340
rect 30492 11330 30548 11340
rect 30828 11396 30884 13132
rect 31052 12962 31108 13244
rect 31052 12910 31054 12962
rect 31106 12910 31108 12962
rect 31052 12180 31108 12910
rect 31052 12114 31108 12124
rect 30828 11330 30884 11340
rect 30940 11508 30996 11518
rect 30940 11355 30996 11452
rect 30940 11303 30942 11355
rect 30994 11303 30996 11355
rect 30940 11291 30996 11303
rect 31164 11394 31220 11406
rect 31164 11342 31166 11394
rect 31218 11342 31220 11394
rect 31164 11284 31220 11342
rect 31164 11218 31220 11228
rect 31276 11226 31332 11238
rect 31276 11174 31278 11226
rect 31330 11174 31332 11226
rect 30380 10220 30660 10276
rect 30492 10052 30548 10062
rect 30156 10050 30548 10052
rect 30156 9998 30494 10050
rect 30546 9998 30548 10050
rect 30156 9996 30548 9998
rect 30492 9986 30548 9996
rect 30604 9044 30660 10220
rect 30828 9828 30884 9838
rect 31276 9828 31332 11174
rect 30828 9826 31332 9828
rect 30828 9774 30830 9826
rect 30882 9774 31332 9826
rect 30828 9772 31332 9774
rect 31388 9828 31444 13692
rect 31724 13524 31780 13534
rect 31948 13524 32004 13534
rect 31500 12964 31556 12974
rect 31500 12178 31556 12908
rect 31500 12126 31502 12178
rect 31554 12126 31556 12178
rect 31500 12114 31556 12126
rect 31724 12178 31780 13468
rect 31836 13468 31948 13524
rect 31836 13074 31892 13468
rect 31948 13458 32004 13468
rect 31836 13022 31838 13074
rect 31890 13022 31892 13074
rect 31836 13010 31892 13022
rect 31724 12126 31726 12178
rect 31778 12126 31780 12178
rect 31724 12114 31780 12126
rect 31948 12740 32004 12750
rect 31948 12190 32004 12684
rect 32060 12404 32116 15820
rect 32620 14868 32676 14878
rect 32620 14754 32676 14812
rect 32620 14702 32622 14754
rect 32674 14702 32676 14754
rect 32620 14690 32676 14702
rect 32284 14532 32340 14542
rect 32284 14438 32340 14476
rect 32620 13748 32676 13758
rect 32620 13654 32676 13692
rect 32284 13524 32340 13534
rect 32284 13430 32340 13468
rect 32060 12338 32116 12348
rect 32564 12404 32620 12414
rect 32956 12404 33012 17052
rect 33068 15988 33124 17164
rect 33236 16996 33292 17006
rect 33236 16212 33292 16940
rect 33404 16882 33460 17612
rect 34524 17668 34580 18396
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35028 17892 35084 17902
rect 35028 17798 35084 17836
rect 35420 17780 35476 17790
rect 34524 17602 34580 17612
rect 35308 17668 35364 17678
rect 35308 17574 35364 17612
rect 35420 17666 35476 17724
rect 35420 17614 35422 17666
rect 35474 17614 35476 17666
rect 35420 17602 35476 17614
rect 35644 17666 35700 17678
rect 35644 17614 35646 17666
rect 35698 17614 35700 17666
rect 33404 16830 33406 16882
rect 33458 16830 33460 16882
rect 33404 16818 33460 16830
rect 34188 17444 34244 17454
rect 34188 16770 34244 17388
rect 34188 16718 34190 16770
rect 34242 16718 34244 16770
rect 34188 16706 34244 16718
rect 34412 17332 34468 17342
rect 34412 16884 34468 17276
rect 33236 16146 33292 16156
rect 34412 16100 34468 16828
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 34524 16100 34580 16110
rect 34412 16098 34580 16100
rect 34412 16046 34526 16098
rect 34578 16046 34580 16098
rect 34412 16044 34580 16046
rect 34524 16034 34580 16044
rect 35084 16098 35140 16110
rect 35084 16046 35086 16098
rect 35138 16046 35140 16098
rect 33068 15932 33460 15988
rect 33124 15652 33180 15662
rect 33124 15426 33180 15596
rect 33124 15374 33126 15426
rect 33178 15374 33180 15426
rect 33124 15362 33180 15374
rect 33404 15314 33460 15932
rect 33404 15262 33406 15314
rect 33458 15262 33460 15314
rect 33404 14644 33460 15262
rect 33628 15986 33684 15998
rect 33628 15934 33630 15986
rect 33682 15934 33684 15986
rect 33628 15316 33684 15934
rect 34188 15876 34244 15886
rect 34076 15874 34244 15876
rect 34076 15822 34190 15874
rect 34242 15822 34244 15874
rect 34076 15820 34244 15822
rect 33628 15222 33684 15260
rect 33964 15314 34020 15326
rect 33964 15262 33966 15314
rect 34018 15262 34020 15314
rect 33740 15204 33796 15214
rect 33964 15148 34020 15262
rect 33740 14644 33796 15148
rect 33404 14578 33460 14588
rect 33628 14588 33796 14644
rect 33852 15092 34020 15148
rect 34076 15204 34132 15820
rect 34188 15810 34244 15820
rect 34076 15138 34132 15148
rect 34188 15314 34244 15326
rect 34188 15262 34190 15314
rect 34242 15262 34244 15314
rect 34188 15148 34244 15262
rect 34916 15316 34972 15326
rect 34916 15222 34972 15260
rect 35084 15204 35140 16046
rect 35532 16042 35588 16054
rect 35532 15990 35534 16042
rect 35586 15990 35588 16042
rect 34188 15092 34356 15148
rect 33628 13746 33684 14588
rect 33852 14530 33908 15092
rect 34300 14868 34356 15092
rect 34468 15092 34524 15102
rect 34468 14998 34524 15036
rect 33852 14478 33854 14530
rect 33906 14478 33908 14530
rect 33628 13694 33630 13746
rect 33682 13694 33684 13746
rect 33516 13524 33572 13534
rect 32564 12310 32620 12348
rect 32844 12348 33012 12404
rect 33068 12852 33124 12862
rect 31948 12178 32060 12190
rect 31948 12126 32006 12178
rect 32058 12126 32060 12178
rect 31948 12124 32060 12126
rect 32004 12114 32060 12124
rect 32620 12068 32676 12078
rect 32620 11618 32676 12012
rect 32620 11566 32622 11618
rect 32674 11566 32676 11618
rect 32620 11554 32676 11566
rect 31724 11508 31780 11518
rect 31724 11414 31780 11452
rect 31836 11396 31892 11406
rect 31836 11327 31838 11340
rect 31890 11327 31892 11340
rect 31836 10724 31892 11327
rect 31836 10658 31892 10668
rect 32172 11394 32228 11406
rect 32172 11342 32174 11394
rect 32226 11342 32228 11394
rect 32060 10612 32116 10622
rect 32172 10612 32228 11342
rect 32844 10836 32900 12348
rect 32956 12180 33012 12190
rect 32956 12086 33012 12124
rect 32956 11396 33012 11406
rect 33068 11396 33124 12796
rect 33516 11508 33572 13468
rect 33628 12852 33684 13694
rect 33740 13914 33796 13926
rect 33740 13862 33742 13914
rect 33794 13862 33796 13914
rect 33740 13748 33796 13862
rect 33740 13682 33796 13692
rect 33740 13076 33796 13086
rect 33852 13076 33908 14478
rect 34076 14812 34356 14868
rect 34076 14515 34132 14812
rect 34300 14756 34356 14812
rect 34300 14700 34916 14756
rect 34076 14463 34078 14515
rect 34130 14463 34132 14515
rect 34076 14451 34132 14463
rect 34188 14642 34244 14654
rect 34188 14590 34190 14642
rect 34242 14590 34244 14642
rect 34188 14196 34244 14590
rect 34076 14140 34244 14196
rect 34300 14532 34356 14542
rect 34076 13802 34132 14140
rect 34076 13750 34078 13802
rect 34130 13750 34132 13802
rect 34076 13738 34132 13750
rect 34300 13746 34356 14476
rect 34300 13694 34302 13746
rect 34354 13694 34356 13746
rect 34300 13682 34356 13694
rect 33740 13074 33908 13076
rect 33740 13022 33742 13074
rect 33794 13022 33908 13074
rect 33740 13020 33908 13022
rect 33740 13010 33796 13020
rect 34188 12962 34244 12974
rect 34188 12910 34190 12962
rect 34242 12910 34244 12962
rect 34860 12962 34916 14700
rect 35084 14532 35140 15148
rect 35196 15314 35252 15326
rect 35196 15262 35198 15314
rect 35250 15262 35252 15314
rect 35196 15092 35252 15262
rect 35420 15314 35476 15326
rect 35420 15262 35422 15314
rect 35474 15262 35476 15314
rect 35420 15092 35476 15262
rect 35532 15204 35588 15990
rect 35644 15930 35700 17614
rect 35980 17444 36036 17454
rect 35980 17350 36036 17388
rect 35756 16772 35812 16782
rect 35756 16098 35812 16716
rect 35756 16046 35758 16098
rect 35810 16046 35812 16098
rect 35756 16034 35812 16046
rect 36092 16770 36148 16782
rect 36092 16718 36094 16770
rect 36146 16718 36148 16770
rect 35644 15878 35646 15930
rect 35698 15878 35700 15930
rect 35644 15866 35700 15878
rect 35756 15329 35812 15392
rect 35756 15316 35758 15329
rect 35810 15316 35812 15329
rect 35644 15204 35700 15214
rect 35532 15202 35700 15204
rect 35532 15150 35646 15202
rect 35698 15150 35700 15202
rect 35532 15148 35700 15150
rect 35644 15138 35700 15148
rect 35420 15036 35588 15092
rect 35196 15026 35252 15036
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35532 14756 35588 15036
rect 35196 14532 35252 14542
rect 35084 14530 35252 14532
rect 35084 14478 35198 14530
rect 35250 14478 35252 14530
rect 35084 14476 35252 14478
rect 35196 14466 35252 14476
rect 35308 13860 35364 13870
rect 35532 13860 35588 14700
rect 35644 14644 35700 14654
rect 35644 14491 35700 14588
rect 35644 14439 35646 14491
rect 35698 14439 35700 14491
rect 35756 14532 35812 15260
rect 36092 15316 36148 16718
rect 36204 16324 36260 19964
rect 36540 19236 36596 20748
rect 36652 19348 36708 21308
rect 37436 20804 37492 21532
rect 37324 20802 37492 20804
rect 37324 20750 37438 20802
rect 37490 20750 37492 20802
rect 37324 20748 37492 20750
rect 37100 20578 37156 20590
rect 37100 20526 37102 20578
rect 37154 20526 37156 20578
rect 36652 19282 36708 19292
rect 36988 19794 37044 19806
rect 36988 19742 36990 19794
rect 37042 19742 37044 19794
rect 36540 19142 36596 19180
rect 36652 18788 36708 18798
rect 36428 18452 36484 18462
rect 36428 18358 36484 18396
rect 36652 17118 36708 18732
rect 36988 18676 37044 19742
rect 37100 19460 37156 20526
rect 37100 19394 37156 19404
rect 36876 18564 36932 18574
rect 36876 17666 36932 18508
rect 36876 17614 36878 17666
rect 36930 17614 36932 17666
rect 36652 17106 36764 17118
rect 36652 17054 36710 17106
rect 36762 17054 36764 17106
rect 36652 17052 36764 17054
rect 36708 17042 36764 17052
rect 36204 16258 36260 16268
rect 36764 16772 36820 16782
rect 36484 16212 36540 16222
rect 36484 16118 36540 16156
rect 36764 15438 36820 16716
rect 36876 16098 36932 17614
rect 36988 16212 37044 18620
rect 37100 19236 37156 19246
rect 37100 18564 37156 19180
rect 37100 18452 37156 18508
rect 37212 18452 37268 18462
rect 37100 18450 37268 18452
rect 37100 18398 37214 18450
rect 37266 18398 37268 18450
rect 37100 18396 37268 18398
rect 37212 18386 37268 18396
rect 37156 17108 37212 17118
rect 37324 17108 37380 20748
rect 37436 20738 37492 20748
rect 37548 21586 37604 21598
rect 37548 21534 37550 21586
rect 37602 21534 37604 21586
rect 37548 21476 37604 21534
rect 37548 20356 37604 21420
rect 37548 20290 37604 20300
rect 37660 20020 37716 22092
rect 37884 22082 37940 22092
rect 37996 21700 38052 22316
rect 37996 21634 38052 21644
rect 38108 22370 38276 22372
rect 38108 22318 38222 22370
rect 38274 22318 38276 22370
rect 38108 22316 38276 22318
rect 37884 21476 37940 21486
rect 37884 21382 37940 21420
rect 37996 20804 38052 20814
rect 38108 20804 38164 22316
rect 38220 22306 38276 22316
rect 38444 21812 38500 23100
rect 38556 22932 38612 24108
rect 38668 23910 38724 24558
rect 38668 23858 38670 23910
rect 38722 23858 38724 23910
rect 38668 23846 38724 23858
rect 38780 24712 39172 24768
rect 38668 23156 38724 23166
rect 38668 23062 38724 23100
rect 38556 22876 38724 22932
rect 38556 21812 38612 21822
rect 38444 21810 38612 21812
rect 38444 21758 38558 21810
rect 38610 21758 38612 21810
rect 38444 21756 38612 21758
rect 38220 21700 38276 21710
rect 38220 21586 38276 21644
rect 38220 21534 38222 21586
rect 38274 21534 38276 21586
rect 38220 21476 38276 21534
rect 38220 21410 38276 21420
rect 37996 20802 38164 20804
rect 37996 20750 37998 20802
rect 38050 20750 38164 20802
rect 37996 20748 38164 20750
rect 37996 20738 38052 20748
rect 37828 20580 37884 20590
rect 38444 20580 38500 21756
rect 38556 21746 38612 21756
rect 37828 20578 38500 20580
rect 37828 20526 37830 20578
rect 37882 20526 38500 20578
rect 37828 20524 38500 20526
rect 37828 20514 37884 20524
rect 37660 19954 37716 19964
rect 38108 20356 38164 20366
rect 37884 19908 37940 19918
rect 37884 19346 37940 19852
rect 37884 19294 37886 19346
rect 37938 19294 37940 19346
rect 37884 19282 37940 19294
rect 37660 18564 37716 18574
rect 37660 18450 37716 18508
rect 37660 18398 37662 18450
rect 37714 18398 37716 18450
rect 37660 18386 37716 18398
rect 38108 18340 38164 20300
rect 38556 20033 38612 20058
rect 38556 20020 38558 20033
rect 38610 20020 38612 20033
rect 38556 19954 38612 19964
rect 38444 19908 38500 19918
rect 38444 19814 38500 19852
rect 38668 19796 38724 22876
rect 38780 21812 38836 24712
rect 39172 24610 39228 24622
rect 39172 24558 39174 24610
rect 39226 24558 39228 24610
rect 39172 24164 39228 24558
rect 39172 24098 39228 24108
rect 39340 23940 39396 25452
rect 39788 25172 39844 26236
rect 40012 25618 40068 26798
rect 40180 26852 40516 26908
rect 41356 26852 41860 26908
rect 40180 26402 40236 26852
rect 40180 26350 40182 26402
rect 40234 26350 40236 26402
rect 40180 26338 40236 26350
rect 40012 25566 40014 25618
rect 40066 25566 40068 25618
rect 40012 25554 40068 25566
rect 41132 26290 41188 26302
rect 41132 26238 41134 26290
rect 41186 26238 41188 26290
rect 39452 24892 39732 24948
rect 39452 24778 39508 24892
rect 39452 24726 39454 24778
rect 39506 24726 39508 24778
rect 39452 24714 39508 24726
rect 39564 24750 39620 24762
rect 39564 24698 39566 24750
rect 39618 24698 39620 24750
rect 39564 24052 39620 24698
rect 39564 23986 39620 23996
rect 39452 23940 39508 23950
rect 38892 23882 38948 23894
rect 39340 23884 39452 23940
rect 38892 23830 38894 23882
rect 38946 23830 38948 23882
rect 39452 23846 39508 23884
rect 38892 22484 38948 23830
rect 39172 23828 39228 23838
rect 39004 23826 39228 23828
rect 39004 23774 39174 23826
rect 39226 23774 39228 23826
rect 39004 23772 39228 23774
rect 39004 23154 39060 23772
rect 39172 23762 39228 23772
rect 39004 23102 39006 23154
rect 39058 23102 39060 23154
rect 39004 23090 39060 23102
rect 39676 23380 39732 24892
rect 39788 24769 39844 25116
rect 40012 25396 40068 25406
rect 40012 24778 40068 25340
rect 39788 24757 39900 24769
rect 39788 24712 39846 24757
rect 39844 24705 39846 24712
rect 39898 24705 39900 24757
rect 40012 24726 40014 24778
rect 40066 24726 40068 24778
rect 40292 25284 40348 25294
rect 40292 24834 40348 25228
rect 41132 25284 41188 26238
rect 41132 25218 41188 25228
rect 40292 24782 40294 24834
rect 40346 24782 40348 24834
rect 40292 24770 40348 24782
rect 41356 24836 41412 26852
rect 42028 26526 42084 29596
rect 42140 28980 42196 30156
rect 42252 30146 42308 30156
rect 42140 28627 42196 28924
rect 42252 28756 42308 28766
rect 42476 28756 42532 30940
rect 42588 30930 42644 30940
rect 42588 29988 42644 29998
rect 42700 29988 42756 29998
rect 42588 29986 42700 29988
rect 42588 29934 42590 29986
rect 42642 29934 42700 29986
rect 42588 29932 42700 29934
rect 42588 29922 42644 29932
rect 42252 28754 42532 28756
rect 42252 28702 42254 28754
rect 42306 28702 42532 28754
rect 42252 28700 42532 28702
rect 42252 28690 42308 28700
rect 42140 28575 42142 28627
rect 42194 28575 42196 28627
rect 42140 28563 42196 28575
rect 42476 28626 42588 28644
rect 42476 28574 42534 28626
rect 42586 28574 42588 28626
rect 42476 28562 42588 28574
rect 42700 28614 42756 29932
rect 42700 28562 42702 28614
rect 42754 28562 42756 28614
rect 42140 28420 42196 28430
rect 42140 26908 42196 28364
rect 42476 27524 42532 28562
rect 42700 28550 42756 28562
rect 42812 29202 42868 30942
rect 42812 29150 42814 29202
rect 42866 29150 42868 29202
rect 42644 28084 42700 28094
rect 42644 27990 42700 28028
rect 42812 27860 42868 29150
rect 42924 30212 42980 30222
rect 43484 30212 43540 31500
rect 43596 31554 43876 31556
rect 43596 31502 43822 31554
rect 43874 31502 43876 31554
rect 43596 31500 43876 31502
rect 43596 30994 43652 31500
rect 43820 31490 43876 31500
rect 43932 31220 43988 31724
rect 44156 31714 44212 31724
rect 44268 31444 44324 32510
rect 44380 32564 44436 32732
rect 44604 32564 44660 32574
rect 44380 32562 44660 32564
rect 44380 32510 44606 32562
rect 44658 32510 44660 32562
rect 44380 32508 44660 32510
rect 44268 31378 44324 31388
rect 43596 30942 43598 30994
rect 43650 30942 43652 30994
rect 43596 30930 43652 30942
rect 43820 31164 43988 31220
rect 44604 31220 44660 32508
rect 44716 32004 44772 34108
rect 44940 34169 44996 34181
rect 44940 34117 44942 34169
rect 44994 34117 44996 34169
rect 44940 33684 44996 34117
rect 44828 33628 44996 33684
rect 44828 33246 44884 33628
rect 44828 33234 44940 33246
rect 44828 33182 44886 33234
rect 44938 33182 44940 33234
rect 44828 33180 44940 33182
rect 44884 33170 44940 33180
rect 45052 33012 45108 37212
rect 45164 36484 45220 36494
rect 45164 36390 45220 36428
rect 45612 36482 45668 36494
rect 45612 36430 45614 36482
rect 45666 36430 45668 36482
rect 45164 35924 45220 35934
rect 45164 35252 45220 35868
rect 45164 34914 45220 35196
rect 45164 34862 45166 34914
rect 45218 34862 45220 34914
rect 45164 34850 45220 34862
rect 45276 35700 45332 35710
rect 45276 35364 45332 35644
rect 45612 35700 45668 36430
rect 45612 35634 45668 35644
rect 45388 35586 45444 35598
rect 45388 35534 45390 35586
rect 45442 35534 45444 35586
rect 45388 35476 45444 35534
rect 45388 35420 45668 35476
rect 45276 34914 45332 35308
rect 45276 34862 45278 34914
rect 45330 34862 45332 34914
rect 45612 35252 45668 35420
rect 45612 34914 45668 35196
rect 45276 34850 45332 34862
rect 45444 34858 45500 34870
rect 45444 34806 45446 34858
rect 45498 34806 45500 34858
rect 45444 34804 45500 34806
rect 45444 34738 45500 34748
rect 45612 34862 45614 34914
rect 45666 34862 45668 34914
rect 45612 34580 45668 34862
rect 45220 34524 45668 34580
rect 45220 34186 45276 34524
rect 45220 34134 45222 34186
rect 45274 34134 45276 34186
rect 45500 34244 45556 34254
rect 45724 34244 45780 38612
rect 45836 38276 45892 38892
rect 45948 38722 46004 39116
rect 45948 38670 45950 38722
rect 46002 38670 46004 38722
rect 45948 38658 46004 38670
rect 46508 38722 46564 38734
rect 46508 38670 46510 38722
rect 46562 38670 46564 38722
rect 45948 38276 46004 38286
rect 45836 38274 46004 38276
rect 45836 38222 45950 38274
rect 46002 38222 46004 38274
rect 45836 38220 46004 38222
rect 45948 38210 46004 38220
rect 46508 38276 46564 38670
rect 46508 38210 46564 38220
rect 46620 38612 46676 38622
rect 46060 38164 46116 38174
rect 45948 37492 46004 37502
rect 46060 37492 46116 38108
rect 46620 38162 46676 38556
rect 46620 38110 46622 38162
rect 46674 38110 46676 38162
rect 46620 38098 46676 38110
rect 46732 38164 46788 43484
rect 47068 43538 47348 43540
rect 47068 43486 47294 43538
rect 47346 43486 47348 43538
rect 47068 43484 47348 43486
rect 46956 43316 47012 43326
rect 46956 43222 47012 43260
rect 46956 41524 47012 41534
rect 46956 40516 47012 41468
rect 46956 40402 47012 40460
rect 46956 40350 46958 40402
rect 47010 40350 47012 40402
rect 46956 40338 47012 40350
rect 47068 40964 47124 43484
rect 47292 43474 47348 43484
rect 47180 43092 47236 43102
rect 47180 42866 47236 43036
rect 47180 42814 47182 42866
rect 47234 42814 47236 42866
rect 47180 42802 47236 42814
rect 47404 40964 47460 45052
rect 47516 44324 47572 45222
rect 47740 45145 47796 45157
rect 47740 45093 47742 45145
rect 47794 45093 47796 45145
rect 47516 44258 47572 44268
rect 47628 44548 47684 44558
rect 47628 44307 47684 44492
rect 47740 44434 47796 45093
rect 47964 45108 48020 45118
rect 47964 45014 48020 45052
rect 48300 44660 48356 47180
rect 48972 47234 49028 47246
rect 48972 47182 48974 47234
rect 49026 47182 49028 47234
rect 48972 47124 49028 47182
rect 48972 47058 49028 47068
rect 48636 46676 48692 46686
rect 48636 46582 48692 46620
rect 48972 46564 49028 46574
rect 48972 46470 49028 46508
rect 49084 45778 49140 45790
rect 49084 45726 49086 45778
rect 49138 45726 49140 45778
rect 49084 45332 49140 45726
rect 49084 45266 49140 45276
rect 48636 45220 48692 45230
rect 48636 45106 48692 45164
rect 48636 45054 48638 45106
rect 48690 45054 48692 45106
rect 48636 45042 48692 45054
rect 48860 45106 48916 45118
rect 48860 45054 48862 45106
rect 48914 45054 48916 45106
rect 48300 44594 48356 44604
rect 48860 44548 48916 45054
rect 49140 45108 49196 45118
rect 49140 45014 49196 45052
rect 48860 44482 48916 44492
rect 47740 44382 47742 44434
rect 47794 44382 47796 44434
rect 47740 44370 47796 44382
rect 47628 44255 47630 44307
rect 47682 44255 47684 44307
rect 47628 44243 47684 44255
rect 48300 44322 48356 44334
rect 48300 44270 48302 44322
rect 48354 44270 48356 44322
rect 47852 43553 47908 43565
rect 47516 43540 47572 43550
rect 47516 43446 47572 43484
rect 47852 43501 47854 43553
rect 47906 43501 47908 43553
rect 47852 43204 47908 43501
rect 47852 43138 47908 43148
rect 47964 43426 48020 43438
rect 47964 43374 47966 43426
rect 48018 43374 48020 43426
rect 47964 43092 48020 43374
rect 47964 43026 48020 43036
rect 47964 41972 48020 41982
rect 47964 41878 48020 41916
rect 48300 41972 48356 44270
rect 48636 43540 48692 43550
rect 48524 43538 48692 43540
rect 48524 43486 48638 43538
rect 48690 43486 48692 43538
rect 48524 43484 48692 43486
rect 48300 41906 48356 41916
rect 48412 43204 48468 43214
rect 48300 41524 48356 41534
rect 47404 40908 47888 40964
rect 47068 40404 47124 40908
rect 47068 40338 47124 40348
rect 47832 40458 47888 40908
rect 47832 40406 47834 40458
rect 47886 40406 47888 40458
rect 48076 40740 48132 40750
rect 48076 40514 48132 40684
rect 48076 40462 48078 40514
rect 48130 40462 48132 40514
rect 48076 40450 48132 40462
rect 47832 40292 47888 40406
rect 47832 40236 48244 40292
rect 46956 39844 47012 39854
rect 46956 39618 47012 39788
rect 46956 39566 46958 39618
rect 47010 39566 47012 39618
rect 46956 39554 47012 39566
rect 47068 39732 47124 39742
rect 47068 39618 47124 39676
rect 47068 39566 47070 39618
rect 47122 39566 47124 39618
rect 47628 39730 47684 39742
rect 47628 39678 47630 39730
rect 47682 39678 47684 39730
rect 47068 39554 47124 39566
rect 47234 39562 47290 39574
rect 47234 39510 47236 39562
rect 47288 39510 47290 39562
rect 47234 39284 47290 39510
rect 47234 39218 47290 39228
rect 47628 39060 47684 39678
rect 48188 39580 48244 40236
rect 48188 39528 48190 39580
rect 48242 39528 48244 39580
rect 48188 39516 48244 39528
rect 48300 39396 48356 41468
rect 48412 40740 48468 43148
rect 48524 41524 48580 43484
rect 48636 43474 48692 43484
rect 48972 43316 49028 43326
rect 48972 43314 49252 43316
rect 48972 43262 48974 43314
rect 49026 43262 49252 43314
rect 48972 43260 49252 43262
rect 48972 43250 49028 43260
rect 49084 42642 49140 42654
rect 49084 42590 49086 42642
rect 49138 42590 49140 42642
rect 48524 41458 48580 41468
rect 48636 41970 48692 41982
rect 48636 41918 48638 41970
rect 48690 41918 48692 41970
rect 48524 41188 48580 41198
rect 48524 41094 48580 41132
rect 48412 40674 48468 40684
rect 48412 40516 48468 40526
rect 48412 39620 48468 40460
rect 48524 39620 48580 39630
rect 48412 39618 48580 39620
rect 48412 39566 48526 39618
rect 48578 39566 48580 39618
rect 48412 39564 48580 39566
rect 48524 39554 48580 39564
rect 48300 39330 48356 39340
rect 48636 39172 48692 41918
rect 48972 41748 49028 41758
rect 48972 41654 49028 41692
rect 48748 41188 48804 41198
rect 48748 40290 48804 41132
rect 48860 41076 48916 41086
rect 48860 40964 48916 41020
rect 48860 40908 49028 40964
rect 48748 40238 48750 40290
rect 48802 40238 48804 40290
rect 48748 40226 48804 40238
rect 48860 40417 48916 40429
rect 48860 40365 48862 40417
rect 48914 40365 48916 40417
rect 48860 39956 48916 40365
rect 48748 39900 48916 39956
rect 48748 39730 48804 39900
rect 48972 39844 49028 40908
rect 49084 40628 49140 42590
rect 49084 40562 49140 40572
rect 48748 39678 48750 39730
rect 48802 39678 48804 39730
rect 48748 39666 48804 39678
rect 48916 39788 49028 39844
rect 49084 40402 49140 40414
rect 49084 40350 49086 40402
rect 49138 40350 49140 40402
rect 49084 40292 49140 40350
rect 48916 39674 48972 39788
rect 48916 39622 48918 39674
rect 48970 39622 48972 39674
rect 48916 39610 48972 39622
rect 48636 39116 49028 39172
rect 47292 39004 47684 39060
rect 47292 38881 47348 39004
rect 47068 38869 47124 38881
rect 46732 38098 46788 38108
rect 46844 38836 46900 38846
rect 46284 38050 46340 38062
rect 46284 37998 46286 38050
rect 46338 37998 46340 38050
rect 46284 37828 46340 37998
rect 46844 37940 46900 38780
rect 47068 38817 47070 38869
rect 47122 38817 47124 38869
rect 47068 38668 47124 38817
rect 47236 38869 47348 38881
rect 47236 38817 47238 38869
rect 47290 38817 47348 38869
rect 47236 38780 47348 38817
rect 47068 38612 47236 38668
rect 46284 37762 46340 37772
rect 46396 37884 46900 37940
rect 45948 37490 46116 37492
rect 45948 37438 45950 37490
rect 46002 37438 46116 37490
rect 45948 37436 46116 37438
rect 45948 37426 46004 37436
rect 46284 37268 46340 37278
rect 46396 37268 46452 37884
rect 46284 37266 46452 37268
rect 46284 37214 46286 37266
rect 46338 37214 46452 37266
rect 46284 37212 46452 37214
rect 46620 37492 46676 37502
rect 47180 37492 47236 38612
rect 47292 37828 47348 38780
rect 47404 38862 47460 38874
rect 47404 38836 47406 38862
rect 47458 38836 47460 38862
rect 47678 38862 47734 38874
rect 47678 38810 47680 38862
rect 47732 38836 47734 38862
rect 47732 38810 48580 38836
rect 47678 38780 48580 38810
rect 47404 38770 47460 38780
rect 48524 38668 48580 38780
rect 48636 38834 48692 38846
rect 48636 38782 48638 38834
rect 48690 38782 48692 38834
rect 48636 38724 48692 38782
rect 48860 38836 48916 39116
rect 48972 39058 49028 39116
rect 48972 39006 48974 39058
rect 49026 39006 49028 39058
rect 48972 38994 49028 39006
rect 48860 38770 48916 38780
rect 48636 38668 48804 38724
rect 47908 38610 47964 38622
rect 47908 38558 47910 38610
rect 47962 38558 47964 38610
rect 47908 38500 47964 38558
rect 47908 38434 47964 38444
rect 48300 38612 48580 38668
rect 48188 37828 48244 37838
rect 47292 37772 47908 37828
rect 47740 37604 47796 37614
rect 46620 37266 46676 37436
rect 47068 37434 47124 37446
rect 47180 37436 47348 37492
rect 47068 37382 47070 37434
rect 47122 37382 47124 37434
rect 46788 37322 46844 37334
rect 46788 37270 46790 37322
rect 46842 37270 46844 37322
rect 46788 37268 46844 37270
rect 46620 37214 46622 37266
rect 46674 37214 46676 37266
rect 46284 37202 46340 37212
rect 46620 37202 46676 37214
rect 46732 37212 46844 37268
rect 45836 36482 45892 36494
rect 45836 36430 45838 36482
rect 45890 36430 45892 36482
rect 45836 35924 45892 36430
rect 45836 35858 45892 35868
rect 45948 36484 46004 36494
rect 45836 35698 45892 35710
rect 45836 35646 45838 35698
rect 45890 35646 45892 35698
rect 45836 35252 45892 35646
rect 45948 35586 46004 36428
rect 46116 36372 46172 36382
rect 46116 36278 46172 36316
rect 46620 36370 46676 36382
rect 46620 36318 46622 36370
rect 46674 36318 46676 36370
rect 45948 35534 45950 35586
rect 46002 35534 46004 35586
rect 45948 35522 46004 35534
rect 46172 35725 46228 35737
rect 46172 35673 46174 35725
rect 46226 35673 46228 35725
rect 45836 35186 45892 35196
rect 46172 34916 46228 35673
rect 46508 35700 46564 35710
rect 46508 35606 46564 35644
rect 46396 34916 46452 34926
rect 46172 34850 46228 34860
rect 46284 34858 46340 34870
rect 46284 34806 46286 34858
rect 46338 34806 46340 34858
rect 46396 34822 46452 34860
rect 46284 34804 46340 34806
rect 46284 34738 46340 34748
rect 46116 34692 46172 34702
rect 45500 34242 45780 34244
rect 45500 34190 45502 34242
rect 45554 34190 45780 34242
rect 45500 34188 45780 34190
rect 45836 34690 46172 34692
rect 45836 34638 46118 34690
rect 46170 34638 46172 34690
rect 45836 34636 46172 34638
rect 45500 34178 45556 34188
rect 45220 34122 45276 34134
rect 45836 33796 45892 34636
rect 46116 34626 46172 34636
rect 45388 33740 45892 33796
rect 45948 34468 46004 34478
rect 46620 34468 46676 36318
rect 46732 36372 46788 37212
rect 46732 35476 46788 36316
rect 46844 35700 46900 35710
rect 46844 35698 47012 35700
rect 46844 35646 46846 35698
rect 46898 35646 47012 35698
rect 46844 35644 47012 35646
rect 46844 35634 46900 35644
rect 46732 35420 46900 35476
rect 46844 34692 46900 35420
rect 46956 35028 47012 35644
rect 46956 34962 47012 34972
rect 47068 34804 47124 37382
rect 47180 37266 47236 37278
rect 47180 37214 47182 37266
rect 47234 37214 47236 37266
rect 47180 35924 47236 37214
rect 47180 35858 47236 35868
rect 47292 35812 47348 37436
rect 47740 37266 47796 37548
rect 47740 37214 47742 37266
rect 47794 37214 47796 37266
rect 47740 37202 47796 37214
rect 47852 37268 47908 37772
rect 48076 37268 48132 37278
rect 47852 37266 48132 37268
rect 47852 37214 48078 37266
rect 48130 37214 48132 37266
rect 47852 37212 48132 37214
rect 48076 37202 48132 37212
rect 48188 37098 48244 37772
rect 48188 37046 48190 37098
rect 48242 37046 48244 37098
rect 48188 37034 48244 37046
rect 47292 35746 47348 35756
rect 47740 36260 47796 36270
rect 47516 35713 47572 35725
rect 47516 35661 47518 35713
rect 47570 35661 47572 35713
rect 47404 35588 47460 35598
rect 47180 35586 47460 35588
rect 47180 35534 47406 35586
rect 47458 35534 47460 35586
rect 47180 35532 47460 35534
rect 47180 35026 47236 35532
rect 47404 35522 47460 35532
rect 47516 35252 47572 35661
rect 47740 35698 47796 36204
rect 47740 35646 47742 35698
rect 47794 35646 47796 35698
rect 47740 35634 47796 35646
rect 47180 34974 47182 35026
rect 47234 34974 47236 35026
rect 47180 34962 47236 34974
rect 47292 35196 47572 35252
rect 47068 34748 47236 34804
rect 46844 34636 47104 34692
rect 46620 34412 46900 34468
rect 45948 34132 46004 34412
rect 46172 34132 46228 34142
rect 45948 34130 46228 34132
rect 45948 34078 46174 34130
rect 46226 34078 46228 34130
rect 45948 34076 46228 34078
rect 45388 33460 45444 33740
rect 45948 33684 46004 34076
rect 46172 34066 46228 34076
rect 45276 33404 45444 33460
rect 45724 33628 46004 33684
rect 44716 31938 44772 31948
rect 44940 32956 45108 33012
rect 45164 33290 45220 33302
rect 45164 33238 45166 33290
rect 45218 33238 45220 33290
rect 44604 31164 44772 31220
rect 43708 30884 43764 30894
rect 43708 30324 43764 30828
rect 43820 30436 43876 31164
rect 44716 30660 44772 31164
rect 44940 30884 44996 32956
rect 44940 30818 44996 30828
rect 45052 32564 45108 32574
rect 44604 30604 44772 30660
rect 44100 30436 44156 30446
rect 43820 30434 44156 30436
rect 43820 30382 44102 30434
rect 44154 30382 44156 30434
rect 43820 30380 44156 30382
rect 44100 30370 44156 30380
rect 43708 30268 43876 30324
rect 43596 30212 43652 30222
rect 42924 28614 42980 30156
rect 43260 30154 43316 30166
rect 43260 30102 43262 30154
rect 43314 30102 43316 30154
rect 43260 30100 43316 30102
rect 43260 30034 43316 30044
rect 43372 30154 43428 30166
rect 43484 30156 43596 30212
rect 43372 30102 43374 30154
rect 43426 30102 43428 30154
rect 43596 30130 43598 30156
rect 43650 30130 43652 30156
rect 43596 30118 43652 30130
rect 43820 30182 43876 30268
rect 43820 30130 43822 30182
rect 43874 30130 43876 30182
rect 43820 30118 43876 30130
rect 43372 29988 43428 30102
rect 43372 29922 43428 29932
rect 44492 29988 44548 29998
rect 44380 29540 44436 29550
rect 44380 29482 44436 29484
rect 44380 29430 44382 29482
rect 44434 29430 44436 29482
rect 44380 29418 44436 29430
rect 44492 29482 44548 29932
rect 44492 29430 44494 29482
rect 44546 29430 44548 29482
rect 44492 29418 44548 29430
rect 43932 28868 43988 28878
rect 43932 28774 43988 28812
rect 42924 28562 42926 28614
rect 42978 28562 42980 28614
rect 42924 28550 42980 28562
rect 43148 28644 43204 28654
rect 44268 28644 44324 28654
rect 43148 28562 43150 28588
rect 43202 28562 43204 28588
rect 43148 28550 43204 28562
rect 43820 28642 44324 28644
rect 43820 28590 44270 28642
rect 44322 28590 44324 28642
rect 43820 28588 44324 28590
rect 43428 28532 43484 28542
rect 42812 27766 42868 27804
rect 43260 28530 43484 28532
rect 43260 28478 43430 28530
rect 43482 28478 43484 28530
rect 43260 28476 43484 28478
rect 42476 27468 43092 27524
rect 42140 26852 42308 26908
rect 42028 26514 42140 26526
rect 42028 26462 42086 26514
rect 42138 26462 42140 26514
rect 42028 26460 42140 26462
rect 42084 26450 42140 26460
rect 42252 26292 42308 26852
rect 42140 26236 42308 26292
rect 42028 26180 42084 26190
rect 41468 26068 41524 26078
rect 41468 26066 41860 26068
rect 41468 26014 41470 26066
rect 41522 26014 41860 26066
rect 41468 26012 41860 26014
rect 41468 26002 41524 26012
rect 41356 24780 41524 24836
rect 40012 24714 40068 24726
rect 41132 24724 41188 24734
rect 41132 24722 41412 24724
rect 39844 24693 39900 24705
rect 41132 24670 41134 24722
rect 41186 24670 41412 24722
rect 41132 24668 41412 24670
rect 41132 24658 41188 24668
rect 40236 24052 40292 24062
rect 40236 23958 40292 23996
rect 41356 23940 41412 24668
rect 39340 22932 39396 22942
rect 38892 22418 38948 22428
rect 39004 22930 39396 22932
rect 39004 22878 39342 22930
rect 39394 22878 39396 22930
rect 39004 22876 39396 22878
rect 39004 22482 39060 22876
rect 39340 22866 39396 22876
rect 39676 22708 39732 23324
rect 40404 23380 40460 23390
rect 40404 23286 40460 23324
rect 40908 23380 40964 23390
rect 40124 23156 40180 23166
rect 39956 23044 40012 23054
rect 39956 22950 40012 22988
rect 39004 22430 39006 22482
rect 39058 22430 39060 22482
rect 39004 22418 39060 22430
rect 39228 22652 39732 22708
rect 39228 22148 39284 22652
rect 40124 22372 40180 23100
rect 40124 22306 40180 22316
rect 40348 22596 40404 22606
rect 38780 21756 39060 21812
rect 38892 21588 38948 21598
rect 38780 21364 38836 21374
rect 38780 20914 38836 21308
rect 38892 21252 38948 21532
rect 38892 21186 38948 21196
rect 38780 20862 38782 20914
rect 38834 20862 38836 20914
rect 38780 20850 38836 20862
rect 39004 20692 39060 21756
rect 39228 21810 39284 22092
rect 39228 21758 39230 21810
rect 39282 21758 39284 21810
rect 39228 21746 39284 21758
rect 39564 21586 39620 21598
rect 39564 21534 39566 21586
rect 39618 21534 39620 21586
rect 39564 21252 39620 21534
rect 39564 21186 39620 21196
rect 39676 21586 39732 21598
rect 39676 21534 39678 21586
rect 39730 21534 39732 21586
rect 39676 21140 39732 21534
rect 40012 21364 40068 21374
rect 40012 21270 40068 21308
rect 39676 21084 40068 21140
rect 38892 20636 39060 20692
rect 38892 20356 38948 20636
rect 38892 20300 39060 20356
rect 39004 20244 39060 20300
rect 39004 20188 39172 20244
rect 38668 19730 38724 19740
rect 38892 20018 38948 20030
rect 38892 19966 38894 20018
rect 38946 19966 38948 20018
rect 38892 19572 38948 19966
rect 38892 19506 38948 19516
rect 39004 20020 39060 20030
rect 37156 17106 37380 17108
rect 37156 17054 37158 17106
rect 37210 17054 37380 17106
rect 37156 17052 37380 17054
rect 37772 18284 38164 18340
rect 37156 17042 37212 17052
rect 37548 16884 37604 16894
rect 37548 16790 37604 16828
rect 36988 16146 37044 16156
rect 36876 16046 36878 16098
rect 36930 16046 36932 16098
rect 36876 16034 36932 16046
rect 37660 16100 37716 16110
rect 37660 16006 37716 16044
rect 37772 15876 37828 18284
rect 37996 18116 38052 18126
rect 37884 17444 37940 17454
rect 37884 17350 37940 17388
rect 37492 15820 37828 15876
rect 37884 17108 37940 17118
rect 37996 17108 38052 18060
rect 38108 17668 38164 18284
rect 38332 18564 38388 18574
rect 38220 17668 38276 17678
rect 38108 17666 38276 17668
rect 38108 17614 38222 17666
rect 38274 17614 38276 17666
rect 38108 17612 38276 17614
rect 38220 17602 38276 17612
rect 38332 17666 38388 18508
rect 38332 17614 38334 17666
rect 38386 17614 38388 17666
rect 38332 17602 38388 17614
rect 38780 18452 38836 18462
rect 37884 17106 38052 17108
rect 37884 17054 37886 17106
rect 37938 17054 38052 17106
rect 37884 17052 38052 17054
rect 37492 15538 37548 15820
rect 37492 15486 37494 15538
rect 37546 15486 37548 15538
rect 37492 15474 37548 15486
rect 36764 15426 36876 15438
rect 36764 15374 36822 15426
rect 36874 15374 36876 15426
rect 36764 15372 36876 15374
rect 36820 15362 36876 15372
rect 36316 15316 36372 15326
rect 36092 15314 36372 15316
rect 36092 15262 36094 15314
rect 36146 15262 36318 15314
rect 36370 15262 36372 15314
rect 36092 15260 36372 15262
rect 36092 15250 36148 15260
rect 36316 15250 36372 15260
rect 36540 15316 36596 15326
rect 37884 15316 37940 17052
rect 38556 16897 38612 16909
rect 38556 16845 38558 16897
rect 38610 16845 38612 16897
rect 38444 16770 38500 16782
rect 38444 16718 38446 16770
rect 38498 16718 38500 16770
rect 38444 16436 38500 16718
rect 38556 16772 38612 16845
rect 38556 16706 38612 16716
rect 38780 16660 38836 18396
rect 39004 17108 39060 19964
rect 39116 18452 39172 20188
rect 40012 20186 40068 21084
rect 40012 20134 40014 20186
rect 40066 20134 40068 20186
rect 40012 20122 40068 20134
rect 39900 20057 39956 20069
rect 39116 18386 39172 18396
rect 39564 20018 39620 20030
rect 39564 19966 39566 20018
rect 39618 19966 39620 20018
rect 39564 18116 39620 19966
rect 39900 20005 39902 20057
rect 39954 20005 39956 20057
rect 39900 19908 39956 20005
rect 40124 20020 40180 20030
rect 40124 20018 40292 20020
rect 40124 19966 40126 20018
rect 40178 19966 40292 20018
rect 40124 19964 40292 19966
rect 40124 19954 40180 19964
rect 39900 19842 39956 19852
rect 40124 19796 40180 19806
rect 39788 19572 39844 19582
rect 39788 19346 39844 19516
rect 39788 19294 39790 19346
rect 39842 19294 39844 19346
rect 39788 19282 39844 19294
rect 39900 19460 39956 19470
rect 39564 18050 39620 18060
rect 39900 18676 39956 19404
rect 39900 18477 39956 18620
rect 39900 18425 39902 18477
rect 39954 18425 39956 18477
rect 39900 18004 39956 18425
rect 40124 18228 40180 19740
rect 40236 19246 40292 19964
rect 40348 19460 40404 22540
rect 40908 22484 40964 23324
rect 41244 23181 41300 23193
rect 41244 23129 41246 23181
rect 41298 23129 41300 23181
rect 40908 22390 40964 22428
rect 41020 22708 41076 22718
rect 40348 19394 40404 19404
rect 40460 21476 40516 21486
rect 40236 19234 40348 19246
rect 40236 19182 40294 19234
rect 40346 19182 40348 19234
rect 40236 19170 40348 19182
rect 40236 18452 40292 19170
rect 40236 18386 40292 18396
rect 40460 18350 40516 21420
rect 41020 21140 41076 22652
rect 41244 22596 41300 23129
rect 41244 22530 41300 22540
rect 41356 22372 41412 23884
rect 41468 22708 41524 24780
rect 41804 24724 41860 26012
rect 41916 25508 41972 25518
rect 41916 25414 41972 25452
rect 41916 24724 41972 24734
rect 41804 24722 41972 24724
rect 41804 24670 41918 24722
rect 41970 24670 41972 24722
rect 41804 24668 41972 24670
rect 41916 24658 41972 24668
rect 41468 22642 41524 22652
rect 41916 23156 41972 23166
rect 41916 22930 41972 23100
rect 41916 22878 41918 22930
rect 41970 22878 41972 22930
rect 41468 22372 41524 22382
rect 41916 22372 41972 22878
rect 42028 22932 42084 26124
rect 42140 24500 42196 26236
rect 42532 26180 42588 26190
rect 42532 26086 42588 26124
rect 43036 26180 43092 27468
rect 43260 26290 43316 28476
rect 43428 28466 43484 28476
rect 43596 27746 43652 27758
rect 43596 27694 43598 27746
rect 43650 27694 43652 27746
rect 43596 26514 43652 27694
rect 43820 27524 43876 28588
rect 44268 28578 44324 28588
rect 44604 28644 44660 30604
rect 44716 30212 44772 30222
rect 44716 29482 44772 30156
rect 44828 30154 44884 30166
rect 44828 30102 44830 30154
rect 44882 30102 44884 30154
rect 44828 29876 44884 30102
rect 44940 30154 44996 30166
rect 44940 30102 44942 30154
rect 44994 30102 44996 30154
rect 44940 29988 44996 30102
rect 44940 29922 44996 29932
rect 44828 29810 44884 29820
rect 45052 29540 45108 32508
rect 45164 32450 45220 33238
rect 45276 32562 45332 33404
rect 45276 32510 45278 32562
rect 45330 32510 45332 32562
rect 45276 32498 45332 32510
rect 45388 33290 45444 33302
rect 45388 33238 45390 33290
rect 45442 33238 45444 33290
rect 45164 32398 45166 32450
rect 45218 32398 45220 32450
rect 45164 32386 45220 32398
rect 45388 32452 45444 33238
rect 45612 33290 45668 33302
rect 45612 33238 45614 33290
rect 45666 33238 45668 33290
rect 45612 33236 45668 33238
rect 45612 33170 45668 33180
rect 45724 33290 45780 33628
rect 46620 33572 46676 33582
rect 46620 33458 46676 33516
rect 46620 33406 46622 33458
rect 46674 33406 46676 33458
rect 46620 33394 46676 33406
rect 46844 33460 46900 34412
rect 47048 34186 47104 34636
rect 47048 34134 47050 34186
rect 47102 34134 47104 34186
rect 47048 34122 47104 34134
rect 47180 34020 47236 34748
rect 47292 34242 47348 35196
rect 47964 34356 48020 34366
rect 47964 34262 48020 34300
rect 47292 34190 47294 34242
rect 47346 34190 47348 34242
rect 47292 34178 47348 34190
rect 47628 34130 47684 34142
rect 47628 34078 47630 34130
rect 47682 34078 47684 34130
rect 47628 34020 47684 34078
rect 47180 33964 47684 34020
rect 45724 33238 45726 33290
rect 45778 33238 45780 33290
rect 45388 32386 45444 32396
rect 45220 32004 45276 32014
rect 45220 31946 45276 31948
rect 45220 31894 45222 31946
rect 45274 31894 45276 31946
rect 45724 32004 45780 33238
rect 45948 33346 46004 33358
rect 45948 33294 45950 33346
rect 46002 33294 46004 33346
rect 45836 33124 45892 33134
rect 45836 32589 45892 33068
rect 45836 32537 45838 32589
rect 45890 32537 45892 32589
rect 45836 32525 45892 32537
rect 45948 32564 46004 33294
rect 46116 33236 46172 33246
rect 46116 33178 46172 33180
rect 46116 33126 46118 33178
rect 46170 33126 46172 33178
rect 46116 33114 46172 33126
rect 45948 32498 46004 32508
rect 46844 32340 46900 33404
rect 46844 32274 46900 32284
rect 47404 33572 47460 33582
rect 47404 32116 47460 33516
rect 48300 32788 48356 38612
rect 48636 38500 48692 38510
rect 48524 38164 48580 38174
rect 48524 38070 48580 38108
rect 48524 36482 48580 36494
rect 48524 36430 48526 36482
rect 48578 36430 48580 36482
rect 48524 34356 48580 36430
rect 48524 34290 48580 34300
rect 47628 32732 48356 32788
rect 48524 33346 48580 33358
rect 48524 33294 48526 33346
rect 48578 33294 48580 33346
rect 48524 32788 48580 33294
rect 48636 32788 48692 38444
rect 48748 37828 48804 38668
rect 48748 37762 48804 37772
rect 49084 37492 49140 40236
rect 49196 38164 49252 43260
rect 49196 38098 49252 38108
rect 49308 41972 49364 41982
rect 49308 41186 49364 41916
rect 49308 41134 49310 41186
rect 49362 41134 49364 41186
rect 49308 38050 49364 41134
rect 49420 41748 49476 41758
rect 49420 40292 49476 41692
rect 49420 40226 49476 40236
rect 49308 37998 49310 38050
rect 49362 37998 49364 38050
rect 49308 37986 49364 37998
rect 49084 37426 49140 37436
rect 49308 37268 49364 37278
rect 48860 37266 49364 37268
rect 48860 37214 49310 37266
rect 49362 37214 49364 37266
rect 48860 37212 49364 37214
rect 48860 36932 48916 37212
rect 49308 37202 49364 37212
rect 48972 37044 49028 37054
rect 48972 37042 49588 37044
rect 48972 36990 48974 37042
rect 49026 36990 49588 37042
rect 48972 36988 49588 36990
rect 48972 36978 49028 36988
rect 48860 36148 48916 36876
rect 49308 36484 49364 36494
rect 49308 36482 49476 36484
rect 49308 36430 49310 36482
rect 49362 36430 49476 36482
rect 49308 36428 49476 36430
rect 49308 36418 49364 36428
rect 48860 36082 48916 36092
rect 48972 36036 49028 36046
rect 48748 35924 48804 35934
rect 48748 35586 48804 35868
rect 48972 35812 49028 35980
rect 48860 35756 49028 35812
rect 48860 35742 48916 35756
rect 48860 35690 48862 35742
rect 48914 35690 48916 35742
rect 48860 35678 48916 35690
rect 49084 35700 49140 35710
rect 49084 35606 49140 35644
rect 48748 35534 48750 35586
rect 48802 35534 48804 35586
rect 48748 35522 48804 35534
rect 49420 34916 49476 36428
rect 49084 34804 49140 34814
rect 49140 34748 49252 34804
rect 49084 34710 49140 34748
rect 48972 34020 49028 34030
rect 48972 33926 49028 33964
rect 48972 32788 49028 32798
rect 48636 32732 48804 32788
rect 47404 32060 47572 32116
rect 45724 31938 45780 31948
rect 45220 31882 45276 31894
rect 45388 31778 45444 31790
rect 45388 31726 45390 31778
rect 45442 31726 45444 31778
rect 45388 31668 45444 31726
rect 45836 31668 45892 31678
rect 45388 31666 45892 31668
rect 45388 31614 45838 31666
rect 45890 31614 45892 31666
rect 45388 31612 45892 31614
rect 45164 30212 45220 30222
rect 45164 30130 45166 30156
rect 45218 30130 45220 30156
rect 45164 30118 45220 30130
rect 45388 30182 45444 31612
rect 45836 31602 45892 31612
rect 47516 31556 47572 32060
rect 47180 31500 47572 31556
rect 46788 31332 46844 31342
rect 46172 31220 46228 31230
rect 46172 31126 46228 31164
rect 46788 31220 46844 31276
rect 46788 31218 46900 31220
rect 46788 31166 46790 31218
rect 46842 31166 46900 31218
rect 46788 31154 46900 31166
rect 45836 30996 45892 31006
rect 45668 30994 45892 30996
rect 45668 30942 45838 30994
rect 45890 30942 45892 30994
rect 45668 30940 45892 30942
rect 45500 30884 45556 30894
rect 45500 30790 45556 30828
rect 45668 30434 45724 30940
rect 45836 30930 45892 30940
rect 45668 30382 45670 30434
rect 45722 30382 45724 30434
rect 45668 30370 45724 30382
rect 45388 30130 45390 30182
rect 45442 30130 45444 30182
rect 45388 30118 45444 30130
rect 46396 30212 46452 30222
rect 46396 30118 46452 30156
rect 46228 29986 46284 29998
rect 46228 29934 46230 29986
rect 46282 29934 46284 29986
rect 46228 29876 46284 29934
rect 46228 29810 46284 29820
rect 44716 29430 44718 29482
rect 44770 29430 44772 29482
rect 44716 29418 44772 29430
rect 44940 29484 45108 29540
rect 46452 29540 46508 29550
rect 44940 29482 45052 29484
rect 44940 29430 44998 29482
rect 45050 29430 45052 29482
rect 46452 29446 46508 29484
rect 44940 29418 45052 29430
rect 45220 29428 45276 29438
rect 45500 29428 45556 29438
rect 45220 29426 45556 29428
rect 44940 28754 44996 29418
rect 45220 29374 45222 29426
rect 45274 29374 45502 29426
rect 45554 29374 45556 29426
rect 45220 29372 45556 29374
rect 45220 29362 45276 29372
rect 45500 29362 45556 29372
rect 45836 29202 45892 29214
rect 45836 29150 45838 29202
rect 45890 29150 45892 29202
rect 45836 28980 45892 29150
rect 46844 29092 46900 31154
rect 47180 30996 47236 31500
rect 47628 31444 47684 32732
rect 48524 32722 48580 32732
rect 47964 32564 48020 32574
rect 48636 32564 48692 32574
rect 47964 32470 48020 32508
rect 48524 32508 48636 32564
rect 48076 32340 48132 32350
rect 47516 31388 47684 31444
rect 47740 31778 47796 31790
rect 47740 31726 47742 31778
rect 47794 31726 47796 31778
rect 47404 31332 47460 31342
rect 47180 30994 47348 30996
rect 47180 30942 47182 30994
rect 47234 30942 47348 30994
rect 47180 30940 47348 30942
rect 47180 30930 47236 30940
rect 47180 30212 47236 30222
rect 47012 30210 47236 30212
rect 47012 30158 47182 30210
rect 47234 30158 47236 30210
rect 47012 30156 47236 30158
rect 47012 29650 47068 30156
rect 47180 30146 47236 30156
rect 47012 29598 47014 29650
rect 47066 29598 47068 29650
rect 47012 29586 47068 29598
rect 47180 29426 47236 29438
rect 47180 29374 47182 29426
rect 47234 29374 47236 29426
rect 47180 29260 47236 29374
rect 47292 29428 47348 30940
rect 47404 30994 47460 31276
rect 47404 30942 47406 30994
rect 47458 30942 47460 30994
rect 47404 30930 47460 30942
rect 47516 30826 47572 31388
rect 47740 31220 47796 31726
rect 47740 31154 47796 31164
rect 47908 31444 47964 31454
rect 47908 31218 47964 31388
rect 47908 31166 47910 31218
rect 47962 31166 47964 31218
rect 47908 31154 47964 31166
rect 47740 30996 47796 31006
rect 48076 30996 48132 32284
rect 47740 30994 48132 30996
rect 47740 30942 47742 30994
rect 47794 30942 48132 30994
rect 47740 30940 48132 30942
rect 48524 31778 48580 32508
rect 48636 32470 48692 32508
rect 48748 32340 48804 32732
rect 48524 31726 48526 31778
rect 48578 31726 48580 31778
rect 47740 30930 47796 30940
rect 47516 30774 47518 30826
rect 47570 30774 47572 30826
rect 47516 30548 47572 30774
rect 47404 30492 47572 30548
rect 47404 29652 47460 30492
rect 48524 30212 48580 31726
rect 48636 32284 48804 32340
rect 48636 30994 48692 32284
rect 48860 32004 48916 32014
rect 48860 31910 48916 31948
rect 48972 31218 49028 32732
rect 49196 31778 49252 34748
rect 49308 34132 49364 34142
rect 49308 34038 49364 34076
rect 49308 33348 49364 33358
rect 49420 33348 49476 34860
rect 49308 33346 49476 33348
rect 49308 33294 49310 33346
rect 49362 33294 49476 33346
rect 49308 33292 49476 33294
rect 49308 32564 49364 33292
rect 49308 32498 49364 32508
rect 49196 31726 49198 31778
rect 49250 31726 49252 31778
rect 49196 31714 49252 31726
rect 48972 31166 48974 31218
rect 49026 31166 49028 31218
rect 48972 31154 49028 31166
rect 48636 30942 48638 30994
rect 48690 30942 48692 30994
rect 48636 30930 48692 30942
rect 48524 30146 48580 30156
rect 49084 30098 49140 30110
rect 49084 30046 49086 30098
rect 49138 30046 49140 30098
rect 47628 29988 47684 29998
rect 47404 29596 47572 29652
rect 47404 29428 47460 29438
rect 47292 29426 47460 29428
rect 47292 29374 47406 29426
rect 47458 29374 47460 29426
rect 47292 29372 47460 29374
rect 47404 29362 47460 29372
rect 47516 29260 47572 29596
rect 47180 29204 47572 29260
rect 46844 29036 47012 29092
rect 45836 28924 46900 28980
rect 44940 28702 44942 28754
rect 44994 28702 44996 28754
rect 44940 28690 44996 28702
rect 46844 28754 46900 28924
rect 46844 28702 46846 28754
rect 46898 28702 46900 28754
rect 46844 28690 46900 28702
rect 44604 28578 44660 28588
rect 45500 28644 45556 28654
rect 45500 27970 45556 28588
rect 45500 27918 45502 27970
rect 45554 27918 45556 27970
rect 45500 27906 45556 27918
rect 44716 27860 44772 27870
rect 43820 27468 43988 27524
rect 43596 26462 43598 26514
rect 43650 26462 43652 26514
rect 43596 26450 43652 26462
rect 43820 26962 43876 26974
rect 43820 26910 43822 26962
rect 43874 26910 43876 26962
rect 43820 26404 43876 26910
rect 43820 26338 43876 26348
rect 43932 26628 43988 27468
rect 44716 27074 44772 27804
rect 44716 27022 44718 27074
rect 44770 27022 44772 27074
rect 44716 27010 44772 27022
rect 45500 27074 45556 27086
rect 45500 27022 45502 27074
rect 45554 27022 45556 27074
rect 45500 26908 45556 27022
rect 46956 26908 47012 29036
rect 47628 28642 47684 29932
rect 48972 29876 49028 29886
rect 47628 28590 47630 28642
rect 47682 28590 47684 28642
rect 47628 28578 47684 28590
rect 47852 29594 47908 29606
rect 47852 29542 47854 29594
rect 47906 29542 47908 29594
rect 47740 27074 47796 27086
rect 47740 27022 47742 27074
rect 47794 27022 47796 27074
rect 45500 26852 46004 26908
rect 43932 26572 44268 26628
rect 43260 26238 43262 26290
rect 43314 26238 43316 26290
rect 43260 26226 43316 26238
rect 43036 26114 43092 26124
rect 42588 25506 42644 25518
rect 42588 25454 42590 25506
rect 42642 25454 42644 25506
rect 42588 25396 42644 25454
rect 43464 25508 43520 25518
rect 43464 25414 43520 25452
rect 42588 25330 42644 25340
rect 43708 25394 43764 25406
rect 43708 25342 43710 25394
rect 43762 25342 43764 25394
rect 43708 24724 43764 25342
rect 43820 25172 43876 25182
rect 43820 24834 43876 25116
rect 43820 24782 43822 24834
rect 43874 24782 43876 24834
rect 43820 24770 43876 24782
rect 43708 24658 43764 24668
rect 42140 24434 42196 24444
rect 42476 24388 42532 24398
rect 42476 23938 42532 24332
rect 42476 23886 42478 23938
rect 42530 23886 42532 23938
rect 42476 23874 42532 23886
rect 42700 23938 42756 23950
rect 42700 23886 42702 23938
rect 42754 23886 42756 23938
rect 42028 22866 42084 22876
rect 42140 23826 42196 23838
rect 42140 23774 42142 23826
rect 42194 23774 42196 23826
rect 42140 23716 42196 23774
rect 42700 23716 42756 23886
rect 42980 23940 43036 23950
rect 42980 23846 43036 23884
rect 43540 23716 43596 23726
rect 42140 23660 42756 23716
rect 43484 23714 43596 23716
rect 43484 23662 43542 23714
rect 43594 23662 43596 23714
rect 41356 22370 41972 22372
rect 41356 22318 41470 22370
rect 41522 22318 41972 22370
rect 41356 22316 41972 22318
rect 41132 21588 41188 21598
rect 41132 21252 41188 21532
rect 41300 21476 41356 21486
rect 41300 21418 41356 21420
rect 41300 21366 41302 21418
rect 41354 21366 41356 21418
rect 41300 21354 41356 21366
rect 41132 21196 41412 21252
rect 41020 21084 41300 21140
rect 40908 21028 40964 21038
rect 40684 20692 40740 20702
rect 40572 20690 40740 20692
rect 40572 20638 40686 20690
rect 40738 20638 40740 20690
rect 40572 20636 40740 20638
rect 40572 20244 40628 20636
rect 40684 20626 40740 20636
rect 40908 20468 40964 20972
rect 41244 20763 41300 21084
rect 41244 20711 41246 20763
rect 41298 20711 41300 20763
rect 41244 20699 41300 20711
rect 40908 20402 40964 20412
rect 41356 20356 41412 21196
rect 41356 20290 41412 20300
rect 40572 20188 41188 20244
rect 40572 19234 40628 20188
rect 41132 20086 41188 20188
rect 41132 20074 41244 20086
rect 40908 20018 40964 20030
rect 40908 19966 40910 20018
rect 40962 19966 40964 20018
rect 41132 20022 41190 20074
rect 41242 20022 41244 20074
rect 41132 20008 41244 20022
rect 40572 19182 40574 19234
rect 40626 19182 40628 19234
rect 40572 19170 40628 19182
rect 40684 19572 40740 19582
rect 40908 19572 40964 19966
rect 41356 19908 41412 19918
rect 41356 19814 41412 19852
rect 40740 19516 40964 19572
rect 40684 19234 40740 19516
rect 40684 19182 40686 19234
rect 40738 19182 40740 19234
rect 40684 19170 40740 19182
rect 41020 19234 41076 19246
rect 41020 19182 41022 19234
rect 41074 19182 41076 19234
rect 40404 18338 40516 18350
rect 40404 18286 40406 18338
rect 40458 18286 40516 18338
rect 40404 18284 40516 18286
rect 41020 18676 41076 19182
rect 41468 19234 41524 22316
rect 42140 22148 42196 23660
rect 43484 23650 43596 23662
rect 43484 23044 43540 23650
rect 42252 22372 42308 22382
rect 42252 22370 42532 22372
rect 42252 22318 42254 22370
rect 42306 22318 42532 22370
rect 42252 22316 42532 22318
rect 42252 22306 42308 22316
rect 42140 22092 42420 22148
rect 42252 21700 42308 21710
rect 41916 21586 41972 21598
rect 41916 21534 41918 21586
rect 41970 21534 41972 21586
rect 41748 21364 41804 21374
rect 41748 21270 41804 21308
rect 41748 20746 41804 20758
rect 41748 20694 41750 20746
rect 41802 20694 41804 20746
rect 41748 20692 41804 20694
rect 41468 19182 41470 19234
rect 41522 19182 41524 19234
rect 41468 19170 41524 19182
rect 41580 20636 41804 20692
rect 41188 19012 41244 19022
rect 41580 19012 41636 20636
rect 41804 20468 41860 20478
rect 41804 20020 41860 20412
rect 41916 20244 41972 21534
rect 42140 21476 42196 21486
rect 41916 20178 41972 20188
rect 42028 20746 42084 20758
rect 42028 20694 42030 20746
rect 42082 20694 42084 20746
rect 41916 20020 41972 20030
rect 41804 20018 41972 20020
rect 41804 19966 41918 20018
rect 41970 19966 41972 20018
rect 41804 19964 41972 19966
rect 41916 19954 41972 19964
rect 42028 19908 42084 20694
rect 42028 19842 42084 19852
rect 42140 20020 42196 21420
rect 42252 21474 42308 21644
rect 42364 21630 42420 22092
rect 42476 21924 42532 22316
rect 43372 22260 43428 22270
rect 42476 21868 43316 21924
rect 43260 21810 43316 21868
rect 43260 21758 43262 21810
rect 43314 21758 43316 21810
rect 43260 21746 43316 21758
rect 42364 21578 42366 21630
rect 42418 21578 42420 21630
rect 42364 21566 42420 21578
rect 42700 21586 42756 21598
rect 42252 21422 42254 21474
rect 42306 21422 42308 21474
rect 42252 21410 42308 21422
rect 42700 21534 42702 21586
rect 42754 21534 42756 21586
rect 42700 21476 42756 21534
rect 42364 21364 42420 21374
rect 42364 20767 42420 21308
rect 42252 20746 42308 20758
rect 42252 20694 42254 20746
rect 42306 20694 42308 20746
rect 42364 20715 42366 20767
rect 42418 20715 42420 20767
rect 42364 20703 42420 20715
rect 42588 21252 42644 21262
rect 42252 20580 42308 20694
rect 42252 20524 42420 20580
rect 42364 20132 42420 20524
rect 42364 20066 42420 20076
rect 42252 20020 42308 20030
rect 42140 20018 42308 20020
rect 42140 19966 42254 20018
rect 42306 19966 42308 20018
rect 42140 19964 42308 19966
rect 41188 19010 41636 19012
rect 41188 18958 41190 19010
rect 41242 18958 41636 19010
rect 41188 18956 41636 18958
rect 41188 18946 41244 18956
rect 41020 18620 41636 18676
rect 41020 18450 41076 18620
rect 41020 18398 41022 18450
rect 41074 18398 41076 18450
rect 40124 18172 40292 18228
rect 39900 17938 39956 17948
rect 39116 17668 39172 17678
rect 39116 17666 39396 17668
rect 39116 17614 39118 17666
rect 39170 17614 39396 17666
rect 39116 17612 39396 17614
rect 39116 17602 39172 17612
rect 39340 17108 39396 17612
rect 40124 17108 40180 17118
rect 39340 17106 40180 17108
rect 39340 17054 40126 17106
rect 40178 17054 40180 17106
rect 39340 17052 40180 17054
rect 39004 17042 39060 17052
rect 40124 17042 40180 17052
rect 38892 16884 38948 16894
rect 39228 16884 39284 16894
rect 38892 16882 39284 16884
rect 38892 16830 38894 16882
rect 38946 16830 39230 16882
rect 39282 16830 39284 16882
rect 38892 16828 39284 16830
rect 38892 16818 38948 16828
rect 38780 16604 38948 16660
rect 38444 16380 38836 16436
rect 38780 15370 38836 16380
rect 38332 15316 38388 15326
rect 37884 15314 38388 15316
rect 37884 15262 38334 15314
rect 38386 15262 38388 15314
rect 38780 15318 38782 15370
rect 38834 15318 38836 15370
rect 38780 15306 38836 15318
rect 37884 15260 38388 15262
rect 36540 15222 36596 15260
rect 37100 15092 37156 15102
rect 36988 14644 37044 14654
rect 36988 14550 37044 14588
rect 35868 14532 35924 14542
rect 35756 14530 35924 14532
rect 35756 14478 35870 14530
rect 35922 14478 35924 14530
rect 35756 14476 35924 14478
rect 35868 14466 35924 14476
rect 35980 14532 36036 14542
rect 35644 14427 35700 14439
rect 35980 14362 36036 14476
rect 37100 14515 37156 15036
rect 38332 15092 38388 15260
rect 38332 15026 38388 15036
rect 37100 14463 37102 14515
rect 37154 14463 37156 14515
rect 37324 14756 37380 14766
rect 37324 14530 37380 14700
rect 37324 14478 37326 14530
rect 37378 14478 37380 14530
rect 37324 14466 37380 14478
rect 37660 14532 37716 14542
rect 37100 14451 37156 14463
rect 37660 14438 37716 14476
rect 38668 14532 38724 14542
rect 35980 14310 35982 14362
rect 36034 14310 36036 14362
rect 35980 14298 36036 14310
rect 37996 14308 38052 14318
rect 37212 14306 38052 14308
rect 35308 13858 35588 13860
rect 35308 13806 35310 13858
rect 35362 13806 35588 13858
rect 35308 13804 35588 13806
rect 37212 14254 37998 14306
rect 38050 14254 38052 14306
rect 37212 14252 38052 14254
rect 35308 13794 35364 13804
rect 37212 13746 37268 14252
rect 37996 14242 38052 14252
rect 38220 14084 38276 14094
rect 37212 13694 37214 13746
rect 37266 13694 37268 13746
rect 37212 13682 37268 13694
rect 37996 13746 38052 13758
rect 37996 13694 37998 13746
rect 38050 13694 38052 13746
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 37772 13076 37828 13086
rect 37772 12982 37828 13020
rect 34188 12852 34244 12910
rect 34468 12906 34524 12918
rect 33628 12796 34244 12852
rect 34300 12852 34356 12862
rect 34468 12854 34470 12906
rect 34522 12854 34524 12906
rect 34468 12852 34524 12854
rect 34300 12794 34356 12796
rect 34300 12742 34302 12794
rect 34354 12742 34356 12794
rect 34300 12730 34356 12742
rect 34412 12796 34524 12852
rect 34860 12910 34862 12962
rect 34914 12910 34916 12962
rect 34412 12628 34468 12796
rect 33852 12572 34468 12628
rect 33740 12068 33796 12078
rect 33740 11974 33796 12012
rect 33516 11452 33796 11508
rect 32956 11394 33124 11396
rect 32956 11342 32958 11394
rect 33010 11342 33124 11394
rect 32956 11340 33124 11342
rect 33628 11350 33684 11362
rect 32956 11330 33012 11340
rect 33628 11298 33630 11350
rect 33682 11298 33684 11350
rect 33628 11284 33684 11298
rect 33460 11228 33628 11284
rect 32844 10780 33124 10836
rect 32956 10612 33012 10622
rect 32060 10610 33012 10612
rect 32060 10558 32062 10610
rect 32114 10558 32958 10610
rect 33010 10558 33012 10610
rect 32060 10556 33012 10558
rect 32060 10546 32116 10556
rect 32956 10546 33012 10556
rect 32508 10388 32564 10398
rect 32508 9838 32564 10332
rect 31612 9828 31668 9838
rect 31388 9826 31668 9828
rect 31388 9774 31614 9826
rect 31666 9774 31668 9826
rect 31388 9772 31668 9774
rect 30828 9762 30884 9772
rect 31612 9716 31668 9772
rect 32488 9826 32564 9838
rect 32488 9774 32490 9826
rect 32542 9774 32564 9826
rect 32488 9772 32564 9774
rect 33068 9828 33124 10780
rect 33180 10724 33236 10734
rect 33180 10610 33236 10668
rect 33460 10722 33516 11228
rect 33628 11218 33684 11228
rect 33460 10670 33462 10722
rect 33514 10670 33516 10722
rect 33460 10658 33516 10670
rect 33180 10558 33182 10610
rect 33234 10558 33236 10610
rect 33180 9940 33236 10558
rect 33628 10388 33684 10398
rect 33180 9884 33572 9940
rect 33068 9772 33180 9828
rect 33516 9787 33572 9884
rect 32488 9762 32544 9772
rect 33124 9770 33180 9772
rect 31612 9650 31668 9660
rect 32732 9714 32788 9726
rect 32732 9662 32734 9714
rect 32786 9662 32788 9714
rect 31500 9057 31556 9069
rect 30604 8978 30660 8988
rect 30828 9044 30884 9054
rect 30828 9042 31220 9044
rect 30828 8990 30830 9042
rect 30882 8990 31220 9042
rect 30828 8988 31220 8990
rect 30828 8978 30884 8988
rect 29540 8818 29596 8830
rect 30492 8820 30548 8830
rect 29540 8766 29542 8818
rect 29594 8766 29596 8818
rect 29540 8428 29596 8766
rect 29260 8372 29428 8428
rect 29484 8372 29596 8428
rect 30044 8818 30548 8820
rect 30044 8766 30494 8818
rect 30546 8766 30548 8818
rect 30044 8764 30548 8766
rect 29260 8258 29316 8372
rect 29260 8206 29262 8258
rect 29314 8206 29316 8258
rect 29260 8194 29316 8206
rect 29260 7588 29316 7598
rect 29260 7494 29316 7532
rect 28924 7422 28926 7474
rect 28978 7422 28980 7474
rect 28924 7410 28980 7422
rect 29484 7476 29540 8372
rect 30044 8370 30100 8764
rect 30492 8754 30548 8764
rect 30044 8318 30046 8370
rect 30098 8318 30100 8370
rect 30044 8306 30100 8318
rect 31164 7642 31220 8988
rect 31500 9005 31502 9057
rect 31554 9005 31556 9057
rect 31164 7590 31166 7642
rect 31218 7590 31220 7642
rect 31388 8930 31444 8942
rect 31388 8878 31390 8930
rect 31442 8878 31444 8930
rect 31164 7578 31220 7590
rect 31276 7588 31332 7598
rect 31052 7501 31108 7513
rect 29484 7410 29540 7420
rect 30716 7476 30772 7486
rect 28644 7250 28700 7262
rect 28644 7198 28646 7250
rect 28698 7198 28700 7250
rect 28644 6804 28700 7198
rect 28644 6738 28700 6748
rect 29372 6804 29428 6814
rect 27916 6638 27918 6690
rect 27970 6638 27972 6690
rect 27916 6626 27972 6638
rect 27580 6611 27636 6623
rect 26796 6598 26852 6611
rect 26348 6470 26350 6522
rect 26402 6470 26404 6522
rect 26348 6458 26404 6470
rect 27020 6580 27076 6590
rect 25396 6038 25452 6076
rect 25788 6076 25844 6132
rect 25788 6038 25900 6076
rect 26516 6132 26572 6142
rect 26516 6038 26572 6076
rect 24556 5854 24558 5906
rect 24610 5854 24612 5906
rect 24556 5842 24612 5854
rect 23604 5794 23660 5806
rect 23604 5742 23606 5794
rect 23658 5742 23660 5794
rect 23604 5684 23660 5742
rect 24164 5684 24220 5694
rect 23604 5628 23828 5684
rect 23660 5124 23716 5134
rect 23100 5030 23156 5068
rect 23212 5122 23716 5124
rect 23212 5070 23662 5122
rect 23714 5070 23716 5122
rect 23212 5068 23716 5070
rect 22932 4610 22988 4620
rect 22540 4498 22596 4508
rect 22858 4452 22914 4462
rect 22858 4358 22914 4396
rect 23100 4340 23156 4350
rect 23212 4340 23268 5068
rect 23660 5058 23716 5068
rect 23772 5124 23828 5628
rect 24164 5682 24276 5684
rect 24164 5630 24166 5682
rect 24218 5630 24276 5682
rect 24164 5618 24276 5630
rect 23100 4338 23268 4340
rect 23100 4286 23102 4338
rect 23154 4286 23268 4338
rect 23604 4676 23660 4686
rect 23604 4394 23660 4620
rect 23604 4342 23606 4394
rect 23658 4342 23660 4394
rect 23772 4452 23828 5068
rect 23772 4358 23828 4396
rect 23604 4330 23660 4342
rect 24220 4338 24276 5618
rect 24444 5124 24500 5134
rect 24444 4564 24500 5068
rect 25564 5124 25620 5134
rect 25564 5030 25620 5068
rect 25396 4676 25452 4686
rect 24556 4564 24612 4574
rect 24444 4562 24612 4564
rect 24444 4510 24558 4562
rect 24610 4510 24612 4562
rect 24444 4508 24612 4510
rect 24556 4498 24612 4508
rect 25228 4452 25284 4462
rect 25228 4358 25284 4396
rect 25396 4394 25452 4620
rect 23100 4284 23268 4286
rect 24220 4286 24222 4338
rect 24274 4286 24276 4338
rect 25396 4342 25398 4394
rect 25450 4342 25452 4394
rect 25788 4452 25844 6038
rect 26348 5124 26404 5134
rect 26348 5030 26404 5068
rect 26908 5124 26964 5134
rect 26684 4900 26740 4910
rect 26684 4898 26852 4900
rect 26684 4846 26686 4898
rect 26738 4846 26852 4898
rect 26684 4844 26852 4846
rect 26684 4834 26740 4844
rect 25788 4386 25844 4396
rect 26142 4564 26198 4574
rect 26142 4450 26198 4508
rect 26142 4398 26144 4450
rect 26196 4398 26198 4450
rect 26142 4386 26198 4398
rect 26628 4506 26684 4518
rect 26628 4454 26630 4506
rect 26682 4454 26684 4506
rect 25396 4330 25452 4342
rect 25900 4340 25956 4350
rect 23100 4274 23156 4284
rect 24220 4274 24276 4286
rect 25900 4246 25956 4284
rect 26628 4004 26684 4454
rect 26572 3948 26684 4004
rect 22428 3602 22484 3612
rect 24780 3668 24836 3678
rect 24780 3574 24836 3612
rect 21420 3474 21422 3526
rect 21474 3474 21476 3526
rect 21420 3462 21476 3474
rect 22652 3444 22708 3454
rect 22652 800 22708 3388
rect 23940 3330 23996 3342
rect 23940 3278 23942 3330
rect 23994 3278 23996 3330
rect 23940 2770 23996 3278
rect 26572 2996 26628 3948
rect 26684 3668 26740 3678
rect 26796 3668 26852 4844
rect 26908 4338 26964 5068
rect 27020 5122 27076 6524
rect 29260 6466 29316 6478
rect 29260 6414 29262 6466
rect 29314 6414 29316 6466
rect 27020 5070 27022 5122
rect 27074 5070 27076 5122
rect 27020 5058 27076 5070
rect 27132 5906 27188 5918
rect 27132 5854 27134 5906
rect 27186 5854 27188 5906
rect 27132 5124 27188 5854
rect 27916 5908 27972 5918
rect 27916 5814 27972 5852
rect 29260 5908 29316 6414
rect 29260 5842 29316 5852
rect 29372 5246 29428 6748
rect 30268 6802 30324 6814
rect 30268 6750 30270 6802
rect 30322 6750 30324 6802
rect 29596 6690 29652 6702
rect 29596 6638 29598 6690
rect 29650 6638 29652 6690
rect 29596 6132 29652 6638
rect 29596 6066 29652 6076
rect 29932 6692 29988 6702
rect 29820 6020 29876 6030
rect 29932 6020 29988 6636
rect 30156 6646 30212 6658
rect 30156 6594 30158 6646
rect 30210 6594 30212 6646
rect 30156 6580 30212 6594
rect 30156 6514 30212 6524
rect 30268 6356 30324 6750
rect 30492 6692 30548 6702
rect 30492 6598 30548 6636
rect 30716 6690 30772 7420
rect 31052 7449 31054 7501
rect 31106 7449 31108 7501
rect 31052 7252 31108 7449
rect 31276 7474 31332 7532
rect 31276 7422 31278 7474
rect 31330 7422 31332 7474
rect 31276 7410 31332 7422
rect 31388 7252 31444 8878
rect 31500 8484 31556 9005
rect 31500 8418 31556 8428
rect 31836 9042 31892 9054
rect 31836 8990 31838 9042
rect 31890 8990 31892 9042
rect 31836 8372 31892 8990
rect 32732 8708 32788 9662
rect 33124 9718 33126 9770
rect 33178 9718 33180 9770
rect 33124 9156 33180 9718
rect 33292 9770 33348 9782
rect 33292 9718 33294 9770
rect 33346 9718 33348 9770
rect 33516 9735 33518 9787
rect 33570 9735 33572 9787
rect 33516 9723 33572 9735
rect 33292 9716 33348 9718
rect 33292 9650 33348 9660
rect 33628 9604 33684 10332
rect 33404 9548 33684 9604
rect 33124 9100 33236 9156
rect 32732 8652 33124 8708
rect 33068 8428 33124 8652
rect 33180 8596 33236 9100
rect 33404 9154 33460 9548
rect 33740 9492 33796 11452
rect 33852 11226 33908 12572
rect 34300 11844 34356 11854
rect 33964 11396 34020 11406
rect 34300 11396 34356 11788
rect 34692 11620 34748 11630
rect 34860 11620 34916 12910
rect 35980 12964 36036 12974
rect 37324 12964 37380 12974
rect 35980 12962 36148 12964
rect 35980 12910 35982 12962
rect 36034 12910 36148 12962
rect 35980 12908 36148 12910
rect 35980 12898 36036 12908
rect 35980 12178 36036 12190
rect 35980 12126 35982 12178
rect 36034 12126 36036 12178
rect 35644 12066 35700 12078
rect 35644 12014 35646 12066
rect 35698 12014 35700 12066
rect 35644 11956 35700 12014
rect 35644 11890 35700 11900
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 34692 11618 34916 11620
rect 34692 11566 34694 11618
rect 34746 11566 34916 11618
rect 34692 11564 34916 11566
rect 34692 11554 34748 11564
rect 35980 11508 36036 12126
rect 35980 11442 36036 11452
rect 33964 11394 34356 11396
rect 33964 11342 33966 11394
rect 34018 11342 34302 11394
rect 34354 11342 34356 11394
rect 33964 11340 34356 11342
rect 33964 11330 34020 11340
rect 34300 11330 34356 11340
rect 34412 11394 34468 11406
rect 34412 11342 34414 11394
rect 34466 11342 34468 11394
rect 33852 11174 33854 11226
rect 33906 11174 33908 11226
rect 34412 11284 34468 11342
rect 36092 11294 36148 12908
rect 36988 12962 37380 12964
rect 36988 12910 37326 12962
rect 37378 12910 37380 12962
rect 36988 12908 37380 12910
rect 36316 12740 36372 12750
rect 36316 12738 36820 12740
rect 36316 12686 36318 12738
rect 36370 12686 36820 12738
rect 36316 12684 36820 12686
rect 36316 12674 36372 12684
rect 36764 12178 36820 12684
rect 36764 12126 36766 12178
rect 36818 12126 36820 12178
rect 36764 12114 36820 12126
rect 36540 11956 36596 11966
rect 34412 11218 34468 11228
rect 36036 11282 36148 11294
rect 36036 11230 36038 11282
rect 36090 11230 36148 11282
rect 36036 11228 36148 11230
rect 36204 11396 36260 11406
rect 36036 11218 36092 11228
rect 33852 11162 33908 11174
rect 35252 11172 35308 11182
rect 35700 11172 35756 11182
rect 35252 11170 35756 11172
rect 35252 11118 35254 11170
rect 35306 11118 35702 11170
rect 35754 11118 35756 11170
rect 35252 11116 35756 11118
rect 35252 11106 35308 11116
rect 34356 10948 34412 10958
rect 34356 10834 34412 10892
rect 34356 10782 34358 10834
rect 34410 10782 34412 10834
rect 34356 10164 34412 10782
rect 35700 10724 35756 11116
rect 36204 10948 36260 11340
rect 35700 10658 35756 10668
rect 36092 10892 36260 10948
rect 36316 11394 36372 11406
rect 36316 11342 36318 11394
rect 36370 11342 36372 11394
rect 34972 10625 35028 10637
rect 34356 10098 34412 10108
rect 34636 10610 34692 10622
rect 34636 10558 34638 10610
rect 34690 10558 34692 10610
rect 33404 9102 33406 9154
rect 33458 9102 33460 9154
rect 33404 9090 33460 9102
rect 33516 9436 33796 9492
rect 34076 9714 34132 9726
rect 34076 9662 34078 9714
rect 34130 9662 34132 9714
rect 33180 8530 33236 8540
rect 33516 8428 33572 9436
rect 34076 8428 34132 9662
rect 34636 9268 34692 10558
rect 34972 10573 34974 10625
rect 35026 10573 35028 10625
rect 34860 10052 34916 10062
rect 34972 10052 35028 10573
rect 35308 10610 35364 10622
rect 35308 10558 35310 10610
rect 35362 10558 35364 10610
rect 34860 10050 35028 10052
rect 34860 9998 34862 10050
rect 34914 9998 35028 10050
rect 34860 9996 35028 9998
rect 35084 10498 35140 10510
rect 35084 10446 35086 10498
rect 35138 10446 35140 10498
rect 34860 9986 34916 9996
rect 35084 9604 35140 10446
rect 35308 10388 35364 10558
rect 35308 10322 35364 10332
rect 35476 10388 35532 10398
rect 35476 10386 35588 10388
rect 35476 10334 35478 10386
rect 35530 10334 35588 10386
rect 35476 10322 35588 10334
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35252 10052 35308 10062
rect 35252 9826 35308 9996
rect 35252 9774 35254 9826
rect 35306 9774 35308 9826
rect 35252 9762 35308 9774
rect 35420 9940 35476 9950
rect 35420 9826 35476 9884
rect 35420 9774 35422 9826
rect 35474 9774 35476 9826
rect 35420 9762 35476 9774
rect 35532 9826 35588 10322
rect 35532 9774 35534 9826
rect 35586 9774 35588 9826
rect 35532 9604 35588 9774
rect 35868 10052 35924 10062
rect 35868 9826 35924 9996
rect 35868 9774 35870 9826
rect 35922 9774 35924 9826
rect 35084 9548 35364 9604
rect 35532 9548 35812 9604
rect 33068 8372 33328 8428
rect 31836 8316 32004 8372
rect 31948 8148 32004 8316
rect 32396 8260 32452 8270
rect 31948 8146 32228 8148
rect 31948 8094 31950 8146
rect 32002 8094 32228 8146
rect 31948 8092 32228 8094
rect 31948 8082 32004 8092
rect 31052 7196 31444 7252
rect 31612 7588 31668 7598
rect 30716 6638 30718 6690
rect 30770 6638 30772 6690
rect 30716 6580 30772 6638
rect 30996 6580 31052 6590
rect 30716 6514 30772 6524
rect 30940 6578 31052 6580
rect 30940 6526 30998 6578
rect 31050 6526 31052 6578
rect 30940 6514 31052 6526
rect 30268 6300 30548 6356
rect 29820 6018 29988 6020
rect 29820 5966 29822 6018
rect 29874 5966 29988 6018
rect 30380 6132 30436 6142
rect 30380 6074 30436 6076
rect 30380 6022 30382 6074
rect 30434 6022 30436 6074
rect 30380 6010 30436 6022
rect 29820 5964 29988 5966
rect 30492 5974 30548 6300
rect 29820 5954 29876 5964
rect 30492 5962 30604 5974
rect 30268 5908 30324 5918
rect 30492 5910 30550 5962
rect 30602 5910 30604 5962
rect 30492 5891 30604 5910
rect 30940 5908 30996 6514
rect 30716 5906 30996 5908
rect 30268 5796 30324 5852
rect 28196 5236 28252 5246
rect 27132 5058 27188 5068
rect 27468 5124 27524 5134
rect 26908 4286 26910 4338
rect 26962 4286 26964 4338
rect 26908 4274 26964 4286
rect 26684 3666 26852 3668
rect 26684 3614 26686 3666
rect 26738 3614 26852 3666
rect 26684 3612 26852 3614
rect 26684 3602 26740 3612
rect 27468 3554 27524 5068
rect 27916 5122 27972 5134
rect 27916 5070 27918 5122
rect 27970 5070 27972 5122
rect 27916 5012 27972 5070
rect 27916 4946 27972 4956
rect 28196 5122 28252 5180
rect 28196 5070 28198 5122
rect 28250 5070 28252 5122
rect 27580 4898 27636 4910
rect 27580 4846 27582 4898
rect 27634 4846 27636 4898
rect 27580 4340 27636 4846
rect 28196 4900 28252 5070
rect 28476 5236 28532 5246
rect 28476 5122 28532 5180
rect 28924 5180 29204 5236
rect 28476 5070 28478 5122
rect 28530 5070 28532 5122
rect 28476 5058 28532 5070
rect 28700 5124 28756 5134
rect 28924 5124 28980 5180
rect 28700 5122 28980 5124
rect 28700 5070 28702 5122
rect 28754 5070 28980 5122
rect 28700 5068 28980 5070
rect 28700 5058 28756 5068
rect 29036 5012 29092 5022
rect 28196 4834 28252 4844
rect 28812 4900 28868 4910
rect 27692 4340 27748 4350
rect 27580 4338 27748 4340
rect 27580 4286 27694 4338
rect 27746 4286 27748 4338
rect 27580 4284 27748 4286
rect 27692 4274 27748 4284
rect 27468 3502 27470 3554
rect 27522 3502 27524 3554
rect 27468 3490 27524 3502
rect 28812 3556 28868 4844
rect 28812 3490 28868 3500
rect 27748 3444 27804 3454
rect 27748 3386 27804 3388
rect 27748 3334 27750 3386
rect 27802 3334 27804 3386
rect 29036 3386 29092 4956
rect 29148 4564 29204 5180
rect 29316 5234 29428 5246
rect 29316 5182 29318 5234
rect 29370 5182 29428 5234
rect 29316 5180 29428 5182
rect 29708 5740 30324 5796
rect 30716 5854 30942 5906
rect 30994 5854 30996 5906
rect 30716 5852 30996 5854
rect 29316 5170 29372 5180
rect 29484 5124 29540 5134
rect 29484 5030 29540 5068
rect 29148 4508 29652 4564
rect 29596 4450 29652 4508
rect 29596 4398 29598 4450
rect 29650 4398 29652 4450
rect 29484 3668 29540 3678
rect 29148 3556 29204 3566
rect 29148 3462 29204 3500
rect 29484 3527 29540 3612
rect 29484 3475 29486 3527
rect 29538 3475 29540 3527
rect 29596 3556 29652 4398
rect 29596 3490 29652 3500
rect 29708 3554 29764 5740
rect 30716 5236 30772 5852
rect 30940 5842 30996 5852
rect 31500 6466 31556 6478
rect 31500 6414 31502 6466
rect 31554 6414 31556 6466
rect 30492 5124 30548 5134
rect 30492 5030 30548 5068
rect 30716 4900 30772 5180
rect 31388 5460 31444 5470
rect 30492 4844 30772 4900
rect 31164 5124 31220 5134
rect 29708 3502 29710 3554
rect 29762 3502 29764 3554
rect 29708 3490 29764 3502
rect 30156 3556 30212 3566
rect 29484 3463 29540 3475
rect 30156 3462 30212 3500
rect 30492 3539 30548 4844
rect 31164 4562 31220 5068
rect 31164 4510 31166 4562
rect 31218 4510 31220 4562
rect 31164 4498 31220 4510
rect 31276 5122 31332 5134
rect 31276 5070 31278 5122
rect 31330 5070 31332 5122
rect 31052 3780 31108 3790
rect 31276 3780 31332 5070
rect 31052 3778 31332 3780
rect 31052 3726 31054 3778
rect 31106 3726 31332 3778
rect 31052 3724 31332 3726
rect 31052 3714 31108 3724
rect 30604 3668 30660 3678
rect 30604 3574 30660 3612
rect 30492 3487 30494 3539
rect 30546 3487 30548 3539
rect 31388 3554 31444 5404
rect 31500 4900 31556 6414
rect 31612 5908 31668 7532
rect 31780 7476 31836 7486
rect 31780 7382 31836 7420
rect 32060 7474 32116 7486
rect 32060 7422 32062 7474
rect 32114 7422 32116 7474
rect 32060 7252 32116 7422
rect 32172 7474 32228 8092
rect 32172 7422 32174 7474
rect 32226 7422 32228 7474
rect 32172 7410 32228 7422
rect 32396 7252 32452 8204
rect 33272 8258 33328 8372
rect 33272 8206 33274 8258
rect 33326 8206 33328 8258
rect 33272 8194 33328 8206
rect 33404 8372 33572 8428
rect 33852 8372 34132 8428
rect 34188 9212 34692 9268
rect 33236 7364 33292 7374
rect 33236 7362 33348 7364
rect 33236 7310 33238 7362
rect 33290 7310 33348 7362
rect 33236 7298 33348 7310
rect 32060 7196 32452 7252
rect 33180 7140 33236 7150
rect 33180 6802 33236 7084
rect 33180 6750 33182 6802
rect 33234 6750 33236 6802
rect 33180 6738 33236 6750
rect 31836 6692 31892 6702
rect 31836 6598 31892 6636
rect 32340 6692 32396 6702
rect 32340 6598 32396 6636
rect 32620 6690 32676 6702
rect 32620 6638 32622 6690
rect 32674 6638 32676 6690
rect 31612 5814 31668 5852
rect 31724 6074 31780 6086
rect 31724 6022 31726 6074
rect 31778 6022 31780 6074
rect 31724 5460 31780 6022
rect 32060 5945 32116 5957
rect 32060 5893 32062 5945
rect 32114 5893 32116 5945
rect 32060 5796 32116 5893
rect 32284 5908 32340 5918
rect 32620 5908 32676 6638
rect 32844 6692 32900 6702
rect 32844 6598 32900 6636
rect 33292 6692 33348 7298
rect 33404 6804 33460 8372
rect 33852 8258 33908 8372
rect 33852 8206 33854 8258
rect 33906 8206 33908 8258
rect 33852 8194 33908 8206
rect 34188 8260 34244 9212
rect 35308 9042 35364 9548
rect 35308 8990 35310 9042
rect 35362 8990 35364 9042
rect 35308 8978 35364 8990
rect 35644 8820 35700 8830
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 34188 8194 34244 8204
rect 34748 8260 34804 8270
rect 33516 8148 33572 8158
rect 33516 8054 33572 8092
rect 34188 8034 34244 8046
rect 34188 7982 34190 8034
rect 34242 7982 34244 8034
rect 34188 7700 34244 7982
rect 34188 7634 34244 7644
rect 34748 7476 34804 8204
rect 34916 8260 34972 8270
rect 34916 8166 34972 8204
rect 35644 8260 35700 8764
rect 35756 8260 35812 9548
rect 35868 8820 35924 9774
rect 35868 8754 35924 8764
rect 35980 9940 36036 9950
rect 35980 9826 36036 9884
rect 35980 9774 35982 9826
rect 36034 9774 36036 9826
rect 35868 8260 35924 8270
rect 35756 8258 35924 8260
rect 35756 8206 35870 8258
rect 35922 8206 35924 8258
rect 35756 8204 35924 8206
rect 35980 8260 36036 9774
rect 36092 9044 36148 10892
rect 36316 10062 36372 11342
rect 36540 11394 36596 11900
rect 36540 11342 36542 11394
rect 36594 11342 36596 11394
rect 36540 11330 36596 11342
rect 36876 11396 36932 11406
rect 36764 10836 36820 10846
rect 36876 10836 36932 11340
rect 36764 10834 36932 10836
rect 36764 10782 36766 10834
rect 36818 10782 36932 10834
rect 36764 10780 36932 10782
rect 36764 10770 36820 10780
rect 36988 10164 37044 12908
rect 37324 12898 37380 12908
rect 37660 12918 37716 12930
rect 37660 12866 37662 12918
rect 37714 12866 37716 12918
rect 37660 12404 37716 12866
rect 37660 12348 37940 12404
rect 36988 10098 37044 10108
rect 37772 11508 37828 11518
rect 36260 10050 36372 10062
rect 36260 9998 36262 10050
rect 36314 9998 36372 10050
rect 36260 9996 36372 9998
rect 37156 10052 37212 10062
rect 36260 9986 36316 9996
rect 37156 9938 37212 9996
rect 37772 10052 37828 11452
rect 37772 9986 37828 9996
rect 37156 9886 37158 9938
rect 37210 9886 37212 9938
rect 37156 9874 37212 9886
rect 37660 9828 37716 9838
rect 37884 9828 37940 12348
rect 37996 11396 38052 13694
rect 37996 11330 38052 11340
rect 38108 13076 38164 13086
rect 37660 9826 37940 9828
rect 37660 9774 37662 9826
rect 37714 9774 37940 9826
rect 37660 9772 37940 9774
rect 37660 9762 37716 9772
rect 37884 9604 37940 9772
rect 37996 11172 38052 11182
rect 37996 9826 38052 11116
rect 38108 10276 38164 13020
rect 38220 11508 38276 14028
rect 38668 13748 38724 14476
rect 38780 13748 38836 13758
rect 38668 13746 38836 13748
rect 38668 13694 38782 13746
rect 38834 13694 38836 13746
rect 38668 13692 38836 13694
rect 38780 13682 38836 13692
rect 38892 13746 38948 16604
rect 39228 16212 39284 16828
rect 39340 16882 39396 16894
rect 39340 16830 39342 16882
rect 39394 16830 39396 16882
rect 39340 16772 39396 16830
rect 40124 16884 40180 16894
rect 39340 16706 39396 16716
rect 40012 16772 40068 16782
rect 39620 16660 39676 16670
rect 39620 16658 39844 16660
rect 39620 16606 39622 16658
rect 39674 16606 39844 16658
rect 39620 16604 39844 16606
rect 39620 16594 39676 16604
rect 39564 16212 39620 16222
rect 39228 16210 39620 16212
rect 39228 16158 39566 16210
rect 39618 16158 39620 16210
rect 39228 16156 39620 16158
rect 39564 16146 39620 16156
rect 39116 15540 39172 15550
rect 39116 15482 39172 15484
rect 39116 15430 39118 15482
rect 39170 15430 39172 15482
rect 39116 15418 39172 15430
rect 39340 15484 39732 15540
rect 39004 15316 39060 15326
rect 39340 15316 39396 15484
rect 39004 15314 39396 15316
rect 39004 15262 39006 15314
rect 39058 15262 39396 15314
rect 39004 15260 39396 15262
rect 39004 15250 39060 15260
rect 39228 15092 39284 15102
rect 39228 14530 39284 15036
rect 39060 14474 39116 14486
rect 39060 14422 39062 14474
rect 39114 14422 39116 14474
rect 39228 14478 39230 14530
rect 39282 14478 39284 14530
rect 39228 14466 39284 14478
rect 39060 14420 39116 14422
rect 39060 14364 39172 14420
rect 38892 13694 38894 13746
rect 38946 13694 38948 13746
rect 38500 13524 38556 13534
rect 38500 13430 38556 13468
rect 38892 13076 38948 13694
rect 39116 13636 39172 14364
rect 39228 14362 39284 14374
rect 39228 14310 39230 14362
rect 39282 14310 39284 14362
rect 39228 14308 39284 14310
rect 39228 14242 39284 14252
rect 39340 13790 39396 15260
rect 39564 15314 39620 15326
rect 39564 15262 39566 15314
rect 39618 15262 39620 15314
rect 39564 15148 39620 15262
rect 39676 15316 39732 15484
rect 39788 15316 39844 16604
rect 39900 16098 39956 16110
rect 39900 16046 39902 16098
rect 39954 16046 39956 16098
rect 39900 15540 39956 16046
rect 40012 15764 40068 16716
rect 40124 15876 40180 16828
rect 40236 16772 40292 18172
rect 40404 17892 40460 18284
rect 40404 17826 40460 17836
rect 41020 17778 41076 18398
rect 41244 18465 41300 18490
rect 41244 18452 41246 18465
rect 41298 18452 41300 18465
rect 41244 18386 41300 18396
rect 41580 18450 41636 18620
rect 41580 18398 41582 18450
rect 41634 18398 41636 18450
rect 41580 18386 41636 18398
rect 41804 18452 41860 18462
rect 42140 18452 42196 19964
rect 42252 19954 42308 19964
rect 42588 19918 42644 21196
rect 42700 20468 42756 21420
rect 43148 20914 43204 20926
rect 43148 20862 43150 20914
rect 43202 20862 43204 20914
rect 43148 20804 43204 20862
rect 43372 20814 43428 22204
rect 43484 21364 43540 22988
rect 43802 22932 43858 22942
rect 43596 22930 43858 22932
rect 43596 22878 43804 22930
rect 43856 22878 43858 22930
rect 43596 22876 43858 22878
rect 43596 21586 43652 22876
rect 43802 22866 43858 22876
rect 43932 22708 43988 26572
rect 44212 26514 44268 26572
rect 44212 26462 44214 26514
rect 44266 26462 44268 26514
rect 44212 26450 44268 26462
rect 44044 26404 44100 26414
rect 44044 24724 44100 26348
rect 45108 26404 45164 26414
rect 45108 26346 45164 26348
rect 44940 26292 44996 26302
rect 45108 26294 45110 26346
rect 45162 26294 45164 26346
rect 45108 26282 45164 26294
rect 45276 26290 45332 26302
rect 44940 26198 44996 26236
rect 45276 26238 45278 26290
rect 45330 26238 45332 26290
rect 44324 25844 44380 25854
rect 45276 25844 45332 26238
rect 44324 25618 44380 25788
rect 44884 25788 45332 25844
rect 45388 26290 45444 26302
rect 45388 26238 45390 26290
rect 45442 26238 45444 26290
rect 44884 25730 44940 25788
rect 44884 25678 44886 25730
rect 44938 25678 44940 25730
rect 44884 25666 44940 25678
rect 44324 25566 44326 25618
rect 44378 25566 44380 25618
rect 44324 25554 44380 25566
rect 44716 25506 44772 25518
rect 44716 25454 44718 25506
rect 44770 25454 44772 25506
rect 44716 25284 44772 25454
rect 44716 25218 44772 25228
rect 44828 25508 44884 25518
rect 44566 25172 44622 25182
rect 44566 24760 44622 25116
rect 44268 24724 44324 24734
rect 44044 24722 44324 24724
rect 44044 24670 44270 24722
rect 44322 24670 44324 24722
rect 44044 24668 44324 24670
rect 44044 23938 44100 24668
rect 44268 24658 44324 24668
rect 44380 24724 44436 24734
rect 44566 24708 44568 24760
rect 44620 24708 44622 24760
rect 44566 24696 44622 24708
rect 44380 24630 44436 24668
rect 44828 24164 44884 25452
rect 45388 24836 45444 26238
rect 45668 26068 45724 26078
rect 45668 26066 45892 26068
rect 45668 26014 45670 26066
rect 45722 26014 45892 26066
rect 45668 26012 45892 26014
rect 45668 26002 45724 26012
rect 45836 25508 45892 26012
rect 45948 25620 46004 26852
rect 46284 26852 46340 26862
rect 46116 26458 46172 26470
rect 46116 26406 46118 26458
rect 46170 26406 46172 26458
rect 46116 26292 46172 26406
rect 46116 26226 46172 26236
rect 46284 26290 46340 26796
rect 46732 26852 47012 26908
rect 47404 26964 47460 27002
rect 47404 26898 47460 26908
rect 46284 26238 46286 26290
rect 46338 26238 46340 26290
rect 46284 26226 46340 26238
rect 46620 26292 46676 26302
rect 46060 25620 46116 25630
rect 45948 25618 46116 25620
rect 45948 25566 46062 25618
rect 46114 25566 46116 25618
rect 45948 25564 46116 25566
rect 46060 25554 46116 25564
rect 46620 25620 46676 26236
rect 46732 25844 46788 26852
rect 47628 26292 47684 26302
rect 47740 26292 47796 27022
rect 46732 25778 46788 25788
rect 47236 26234 47292 26246
rect 47236 26182 47238 26234
rect 47290 26182 47292 26234
rect 47684 26236 47796 26292
rect 47628 26198 47684 26236
rect 47236 25732 47292 26182
rect 47180 25676 47292 25732
rect 47404 26178 47460 26190
rect 47404 26126 47406 26178
rect 47458 26126 47460 26178
rect 46620 25618 47012 25620
rect 46620 25566 46622 25618
rect 46674 25566 47012 25618
rect 46620 25564 47012 25566
rect 46620 25554 46676 25564
rect 45836 25506 46004 25508
rect 45612 25450 45668 25462
rect 45612 25398 45614 25450
rect 45666 25398 45668 25450
rect 45836 25454 45838 25506
rect 45890 25454 46004 25506
rect 45836 25452 46004 25454
rect 45836 25442 45892 25452
rect 45612 25172 45668 25398
rect 45612 25106 45668 25116
rect 45388 24770 45444 24780
rect 45836 24836 45892 24846
rect 45836 24722 45892 24780
rect 45836 24670 45838 24722
rect 45890 24670 45892 24722
rect 45836 24658 45892 24670
rect 45948 24722 46004 25452
rect 46228 25452 46284 25462
rect 46228 25450 46452 25452
rect 46228 25398 46230 25450
rect 46282 25398 46452 25450
rect 46228 25396 46452 25398
rect 46228 25386 46284 25396
rect 45948 24670 45950 24722
rect 46002 24670 46004 24722
rect 45948 24658 46004 24670
rect 45556 24612 45612 24622
rect 45556 24610 45780 24612
rect 45556 24558 45558 24610
rect 45610 24558 45780 24610
rect 45556 24556 45780 24558
rect 45556 24546 45612 24556
rect 44940 24500 44996 24510
rect 44940 24498 45162 24500
rect 44940 24446 44942 24498
rect 44994 24446 45162 24498
rect 44940 24444 45162 24446
rect 44940 24434 44996 24444
rect 44044 23886 44046 23938
rect 44098 23886 44100 23938
rect 44044 23874 44100 23886
rect 44716 24108 44884 24164
rect 44212 23828 44268 23838
rect 44212 23770 44268 23772
rect 44212 23718 44214 23770
rect 44266 23718 44268 23770
rect 44212 23706 44268 23718
rect 44548 23268 44604 23278
rect 44548 23210 44604 23212
rect 44044 23154 44100 23166
rect 44044 23102 44046 23154
rect 44098 23102 44100 23154
rect 44548 23158 44550 23210
rect 44602 23158 44604 23210
rect 44548 23146 44604 23158
rect 44716 23266 44772 24108
rect 44828 23938 44884 23950
rect 44828 23886 44830 23938
rect 44882 23886 44884 23938
rect 44828 23828 44884 23886
rect 44828 23762 44884 23772
rect 44940 23938 44996 23950
rect 44940 23886 44942 23938
rect 44994 23886 44996 23938
rect 44716 23214 44718 23266
rect 44770 23214 44772 23266
rect 44044 22932 44100 23102
rect 44044 22866 44100 22876
rect 44716 22708 44772 23214
rect 44940 23380 44996 23886
rect 45106 23938 45162 24444
rect 45106 23886 45108 23938
rect 45160 23886 45162 23938
rect 45106 23874 45162 23886
rect 45500 24050 45556 24062
rect 45500 23998 45502 24050
rect 45554 23998 45556 24050
rect 44940 23154 44996 23324
rect 44940 23102 44942 23154
rect 44994 23102 44996 23154
rect 44940 23090 44996 23102
rect 45388 23156 45444 23166
rect 45388 23062 45444 23100
rect 45108 22932 45164 22942
rect 45108 22838 45164 22876
rect 43596 21534 43598 21586
rect 43650 21534 43652 21586
rect 43596 21522 43652 21534
rect 43820 22652 43988 22708
rect 44604 22652 44772 22708
rect 43820 21476 43876 22652
rect 44492 22596 44548 22606
rect 43820 21410 43876 21420
rect 43988 22372 44044 22382
rect 43988 21474 44044 22316
rect 44156 22260 44212 22270
rect 44156 22166 44212 22204
rect 44492 21822 44548 22540
rect 44436 21810 44548 21822
rect 44436 21758 44438 21810
rect 44490 21758 44548 21810
rect 44436 21756 44548 21758
rect 44436 21746 44492 21756
rect 44604 21700 44660 22652
rect 45500 22484 45556 23998
rect 45724 22596 45780 24556
rect 46228 24500 46284 24510
rect 46060 24498 46284 24500
rect 46060 24446 46230 24498
rect 46282 24446 46284 24498
rect 46060 24444 46284 24446
rect 45724 22530 45780 22540
rect 45948 23268 46004 23278
rect 45948 22594 46004 23212
rect 45948 22542 45950 22594
rect 46002 22542 46004 22594
rect 45948 22530 46004 22542
rect 45500 22428 45668 22484
rect 44828 22370 44884 22382
rect 44828 22318 44830 22370
rect 44882 22318 44884 22370
rect 44828 22260 44884 22318
rect 45612 22372 45668 22428
rect 45612 22339 45760 22372
rect 45612 22316 45706 22339
rect 45704 22287 45706 22316
rect 45758 22287 45760 22339
rect 45704 22275 45760 22287
rect 44828 22194 44884 22204
rect 44604 21634 44660 21644
rect 45500 21700 45556 21710
rect 45500 21630 45556 21644
rect 46060 21700 46116 24444
rect 46228 24434 46284 24444
rect 46396 23716 46452 25396
rect 46956 24722 47012 25564
rect 46956 24670 46958 24722
rect 47010 24670 47012 24722
rect 46956 24658 47012 24670
rect 47068 25172 47124 25182
rect 47068 24610 47124 25116
rect 47068 24558 47070 24610
rect 47122 24558 47124 24610
rect 47068 24546 47124 24558
rect 46732 23940 46788 23950
rect 46732 23846 46788 23884
rect 46956 23938 47012 23950
rect 46956 23886 46958 23938
rect 47010 23886 47012 23938
rect 46956 23716 47012 23886
rect 47180 23940 47236 25676
rect 47292 24749 47348 24761
rect 47292 24697 47294 24749
rect 47346 24697 47348 24749
rect 47292 24164 47348 24697
rect 47404 24724 47460 26126
rect 47852 25844 47908 29542
rect 48860 29540 48916 29550
rect 48076 29428 48132 29438
rect 48076 29334 48132 29372
rect 48244 27746 48300 27758
rect 48244 27694 48246 27746
rect 48298 27694 48300 27746
rect 48244 27188 48300 27694
rect 48860 27300 48916 29484
rect 48972 28082 49028 29820
rect 49084 29428 49140 30046
rect 49084 29362 49140 29372
rect 49252 28420 49308 28430
rect 49252 28418 49364 28420
rect 49252 28366 49254 28418
rect 49306 28366 49364 28418
rect 49252 28354 49364 28366
rect 48972 28030 48974 28082
rect 49026 28030 49028 28082
rect 48972 28018 49028 28030
rect 49308 27858 49364 28354
rect 49308 27806 49310 27858
rect 49362 27806 49364 27858
rect 49308 27636 49364 27806
rect 49308 27570 49364 27580
rect 48972 27300 49028 27310
rect 48860 27298 49028 27300
rect 48860 27246 48974 27298
rect 49026 27246 49028 27298
rect 48860 27244 49028 27246
rect 48972 27234 49028 27244
rect 48244 27122 48300 27132
rect 49308 27188 49364 27198
rect 47964 27074 48020 27086
rect 47964 27022 47966 27074
rect 48018 27022 48020 27074
rect 47964 26328 48020 27022
rect 49308 27074 49364 27132
rect 49308 27022 49310 27074
rect 49362 27022 49364 27074
rect 48244 26962 48300 26974
rect 48244 26910 48246 26962
rect 48298 26910 48300 26962
rect 48244 26908 48300 26910
rect 49308 26908 49364 27022
rect 48244 26852 48468 26908
rect 49308 26852 49476 26908
rect 47964 26276 47966 26328
rect 48018 26276 48020 26328
rect 47964 25844 48020 26276
rect 47964 25788 48356 25844
rect 47852 25778 47908 25788
rect 48300 25284 48356 25788
rect 48188 25228 48356 25284
rect 47404 24658 47460 24668
rect 47628 25172 47684 25182
rect 47628 24836 47684 25116
rect 47628 24722 47684 24780
rect 47628 24670 47630 24722
rect 47682 24670 47684 24722
rect 47628 24658 47684 24670
rect 47964 24722 48020 24734
rect 47964 24670 47966 24722
rect 48018 24670 48020 24722
rect 47964 24388 48020 24670
rect 47964 24322 48020 24332
rect 47292 24108 48132 24164
rect 47628 23940 47684 23950
rect 47180 23874 47236 23884
rect 47404 23882 47460 23894
rect 46284 23714 47012 23716
rect 46284 23662 46398 23714
rect 46450 23662 47012 23714
rect 46284 23660 47012 23662
rect 47404 23830 47406 23882
rect 47458 23830 47460 23882
rect 47628 23846 47684 23884
rect 48076 23938 48132 24108
rect 48076 23886 48078 23938
rect 48130 23886 48132 23938
rect 46172 23044 46228 23054
rect 46172 22950 46228 22988
rect 46060 21634 46116 21644
rect 44884 21588 44940 21598
rect 44884 21494 44940 21532
rect 45276 21586 45332 21598
rect 45276 21534 45278 21586
rect 45330 21534 45332 21586
rect 45500 21578 45502 21630
rect 45554 21578 45556 21630
rect 45500 21566 45556 21578
rect 46172 21588 46228 21598
rect 46284 21588 46340 23660
rect 46396 23650 46452 23660
rect 47404 22708 47460 23830
rect 47740 23770 47796 23782
rect 47740 23718 47742 23770
rect 47794 23718 47796 23770
rect 47740 23156 47796 23718
rect 47740 23090 47796 23100
rect 48076 23266 48132 23886
rect 48188 23940 48244 25228
rect 48412 24724 48468 26852
rect 49196 26290 49252 26302
rect 49196 26238 49198 26290
rect 49250 26238 49252 26290
rect 48860 26068 48916 26078
rect 48524 26066 48916 26068
rect 48524 26014 48862 26066
rect 48914 26014 48916 26066
rect 48524 26012 48916 26014
rect 48524 25618 48580 26012
rect 48860 26002 48916 26012
rect 48524 25566 48526 25618
rect 48578 25566 48580 25618
rect 48524 25554 48580 25566
rect 49196 24846 49252 26238
rect 49140 24834 49252 24846
rect 49140 24782 49142 24834
rect 49194 24782 49252 24834
rect 49140 24780 49252 24782
rect 49308 25506 49364 25518
rect 49308 25454 49310 25506
rect 49362 25454 49364 25506
rect 49140 24770 49196 24780
rect 48636 24724 48692 24734
rect 48412 24722 48692 24724
rect 48412 24670 48638 24722
rect 48690 24670 48692 24722
rect 48412 24668 48692 24670
rect 48636 24658 48692 24668
rect 48860 24724 48916 24734
rect 48860 24630 48916 24668
rect 48748 24388 48804 24398
rect 48188 23874 48244 23884
rect 48300 23938 48356 23950
rect 48300 23886 48302 23938
rect 48354 23886 48356 23938
rect 48300 23716 48356 23886
rect 48580 23940 48636 23950
rect 48580 23846 48636 23884
rect 48300 23660 48580 23716
rect 48076 23214 48078 23266
rect 48130 23214 48132 23266
rect 47404 22652 47684 22708
rect 46732 22596 46788 22606
rect 46732 22342 46788 22540
rect 46732 22290 46734 22342
rect 46786 22290 46788 22342
rect 46732 22278 46788 22290
rect 46620 21754 46676 21766
rect 46620 21702 46622 21754
rect 46674 21702 46676 21754
rect 43988 21422 43990 21474
rect 44042 21422 44044 21474
rect 43484 21308 43652 21364
rect 43372 20802 43447 20814
rect 43372 20750 43393 20802
rect 43445 20750 43447 20802
rect 43372 20748 43447 20750
rect 43148 20738 43204 20748
rect 43391 20738 43447 20748
rect 43596 20692 43652 21308
rect 43988 21252 44044 21422
rect 45276 21364 45332 21534
rect 46228 21532 46340 21588
rect 46396 21625 46452 21637
rect 46396 21573 46398 21625
rect 46450 21573 46452 21625
rect 46172 21494 46228 21532
rect 45612 21476 45668 21486
rect 45612 21474 46116 21476
rect 45612 21422 45614 21474
rect 45666 21422 46116 21474
rect 45612 21420 46116 21422
rect 45612 21410 45668 21420
rect 43988 21186 44044 21196
rect 45052 21308 45276 21364
rect 46060 21364 46116 21420
rect 46396 21364 46452 21573
rect 46060 21308 46452 21364
rect 45052 20914 45108 21308
rect 45276 21298 45332 21308
rect 45052 20862 45054 20914
rect 45106 20862 45108 20914
rect 44268 20804 44324 20814
rect 44268 20710 44324 20748
rect 45052 20804 45108 20862
rect 45052 20738 45108 20748
rect 45836 21252 45892 21262
rect 42700 20402 42756 20412
rect 43484 20636 43652 20692
rect 42920 20132 42976 20142
rect 42920 20056 42976 20076
rect 42920 20004 42922 20056
rect 42974 20004 42976 20056
rect 42588 19908 42700 19918
rect 42588 19852 42644 19908
rect 42644 19814 42700 19852
rect 42920 19572 42976 20004
rect 43484 19796 43540 20636
rect 45836 20580 45892 21196
rect 46620 21140 46676 21702
rect 46844 21586 46900 21598
rect 46844 21534 46846 21586
rect 46898 21534 46900 21586
rect 46620 21084 46788 21140
rect 46732 20580 46788 21084
rect 45836 20524 46228 20580
rect 46060 20244 46116 20254
rect 46060 20150 46116 20188
rect 43596 20132 43652 20142
rect 43596 20018 43652 20076
rect 45332 20132 45388 20142
rect 45332 20038 45388 20076
rect 45948 20132 46004 20142
rect 43596 19966 43598 20018
rect 43650 19966 43652 20018
rect 43596 19954 43652 19966
rect 43708 20020 43764 20030
rect 44044 20020 44100 20030
rect 43708 19850 43764 19964
rect 43708 19798 43710 19850
rect 43762 19798 43764 19850
rect 43708 19786 43764 19798
rect 43932 20018 44100 20020
rect 43932 19966 44046 20018
rect 44098 19966 44100 20018
rect 43932 19964 44100 19966
rect 43484 19730 43540 19740
rect 42920 19506 42976 19516
rect 43484 19460 43540 19470
rect 42252 19236 42308 19246
rect 42252 19234 42532 19236
rect 42252 19182 42254 19234
rect 42306 19182 42532 19234
rect 42252 19180 42532 19182
rect 42252 19170 42308 19180
rect 41804 18358 41860 18396
rect 41916 18396 42196 18452
rect 42364 18450 42420 18462
rect 42364 18398 42366 18450
rect 42418 18398 42420 18450
rect 41356 18340 41412 18350
rect 41356 18338 41524 18340
rect 41356 18286 41358 18338
rect 41410 18286 41524 18338
rect 41356 18284 41524 18286
rect 41356 18274 41412 18284
rect 41020 17726 41022 17778
rect 41074 17726 41076 17778
rect 41020 17714 41076 17726
rect 41356 18116 41412 18126
rect 41356 17668 41412 18060
rect 41468 17892 41524 18284
rect 41804 18228 41860 18238
rect 41468 17836 41748 17892
rect 41468 17668 41524 17678
rect 41356 17666 41524 17668
rect 41356 17614 41470 17666
rect 41522 17614 41524 17666
rect 41356 17612 41524 17614
rect 41692 17668 41748 17836
rect 41804 17780 41860 18172
rect 41916 18004 41972 18396
rect 42364 18340 42420 18398
rect 42364 18274 42420 18284
rect 42084 18228 42140 18238
rect 42084 18226 42308 18228
rect 42084 18174 42086 18226
rect 42138 18174 42308 18226
rect 42084 18172 42308 18174
rect 42084 18162 42140 18172
rect 41916 17948 42084 18004
rect 41804 17724 41972 17780
rect 41692 17612 41804 17668
rect 41468 17602 41524 17612
rect 41748 17610 41804 17612
rect 41748 17558 41750 17610
rect 41802 17558 41804 17610
rect 41748 17546 41804 17558
rect 41580 17498 41636 17510
rect 41580 17446 41582 17498
rect 41634 17446 41636 17498
rect 41580 17220 41636 17446
rect 40460 17164 41636 17220
rect 41692 17444 41748 17454
rect 40460 16882 40516 17164
rect 41076 16996 41132 17006
rect 41076 16902 41132 16940
rect 41692 16899 41748 17388
rect 41916 16996 41972 17724
rect 40460 16830 40462 16882
rect 40514 16830 40516 16882
rect 40460 16818 40516 16830
rect 41244 16884 41300 16894
rect 40236 16706 40292 16716
rect 41132 16212 41188 16222
rect 41244 16212 41300 16828
rect 41132 16210 41300 16212
rect 41132 16158 41134 16210
rect 41186 16158 41300 16210
rect 41132 16156 41300 16158
rect 41468 16843 41748 16899
rect 41804 16940 41972 16996
rect 41132 16146 41188 16156
rect 40236 16100 40292 16110
rect 40236 16006 40292 16044
rect 40124 15820 40292 15876
rect 40012 15708 40180 15764
rect 39900 15474 39956 15484
rect 39676 15314 39844 15316
rect 39676 15262 39678 15314
rect 39730 15262 39844 15314
rect 39676 15260 39844 15262
rect 39676 15250 39732 15260
rect 39564 15092 39844 15148
rect 39788 14644 39844 15092
rect 39340 13738 39342 13790
rect 39394 13738 39396 13790
rect 39340 13726 39396 13738
rect 39676 14642 39844 14644
rect 39676 14590 39790 14642
rect 39842 14590 39844 14642
rect 39676 14588 39844 14590
rect 39676 13746 39732 14588
rect 39788 14578 39844 14588
rect 39956 15090 40012 15102
rect 39956 15038 39958 15090
rect 40010 15038 40012 15090
rect 39956 14532 40012 15038
rect 40124 14756 40180 15708
rect 40124 14690 40180 14700
rect 39956 14466 40012 14476
rect 39676 13694 39678 13746
rect 39730 13694 39732 13746
rect 39676 13682 39732 13694
rect 39900 14308 39956 14318
rect 39900 13746 39956 14252
rect 40236 14196 40292 15820
rect 39900 13694 39902 13746
rect 39954 13694 39956 13746
rect 39900 13682 39956 13694
rect 40012 14140 40292 14196
rect 39228 13636 39284 13646
rect 39116 13634 39284 13636
rect 39116 13582 39230 13634
rect 39282 13582 39284 13634
rect 39116 13580 39284 13582
rect 39228 13570 39284 13580
rect 38892 13010 38948 13020
rect 39396 13076 39452 13086
rect 39396 12982 39452 13020
rect 39900 13076 39956 13086
rect 39900 12982 39956 13020
rect 38220 11442 38276 11452
rect 38332 12962 38388 12974
rect 38332 12910 38334 12962
rect 38386 12910 38388 12962
rect 38108 10210 38164 10220
rect 38220 11284 38276 11294
rect 38332 11284 38388 12910
rect 38220 11282 38388 11284
rect 38220 11230 38222 11282
rect 38274 11230 38388 11282
rect 38220 11228 38388 11230
rect 38556 12962 38612 12974
rect 38556 12910 38558 12962
rect 38610 12910 38612 12962
rect 38220 10612 38276 11228
rect 37996 9774 37998 9826
rect 38050 9774 38052 9826
rect 37996 9762 38052 9774
rect 38220 9787 38276 10556
rect 38444 10637 38500 10649
rect 38444 10585 38446 10637
rect 38498 10585 38500 10637
rect 38332 9940 38388 9950
rect 38332 9846 38388 9884
rect 38220 9735 38222 9787
rect 38274 9735 38276 9787
rect 38220 9723 38276 9735
rect 37884 9548 38388 9604
rect 36204 9044 36260 9054
rect 36092 9042 36260 9044
rect 36092 8990 36094 9042
rect 36146 8990 36206 9042
rect 36258 8990 36260 9042
rect 36092 8988 36260 8990
rect 36092 8978 36148 8988
rect 36204 8978 36260 8988
rect 36988 8930 37044 8942
rect 36988 8878 36990 8930
rect 37042 8878 37044 8930
rect 36988 8484 37044 8878
rect 37548 8708 37604 8718
rect 37212 8484 37268 8494
rect 36988 8482 37268 8484
rect 36988 8430 37214 8482
rect 37266 8430 37268 8482
rect 36988 8428 37268 8430
rect 37212 8418 37268 8428
rect 36316 8370 36372 8382
rect 36316 8318 36318 8370
rect 36370 8318 36372 8370
rect 35980 8228 36204 8260
rect 35980 8204 36150 8228
rect 35644 8166 35700 8204
rect 35868 8194 35924 8204
rect 36148 8176 36150 8204
rect 36202 8176 36204 8228
rect 36148 8164 36204 8176
rect 35308 8036 35364 8046
rect 35308 8034 35588 8036
rect 35308 7982 35310 8034
rect 35362 7982 35588 8034
rect 35308 7980 35588 7982
rect 35308 7970 35364 7980
rect 34860 7476 34916 7486
rect 34748 7420 34860 7476
rect 34860 7382 34916 7420
rect 34972 7476 35028 7486
rect 35196 7476 35252 7486
rect 34972 7474 35252 7476
rect 34972 7422 34974 7474
rect 35026 7422 35198 7474
rect 35250 7422 35252 7474
rect 34972 7420 35252 7422
rect 33684 7362 33740 7374
rect 33684 7310 33686 7362
rect 33738 7310 33740 7362
rect 33684 7252 33740 7310
rect 34244 7364 34300 7374
rect 34244 7252 34300 7308
rect 33684 7196 34300 7252
rect 34580 7252 34636 7262
rect 34580 7250 34916 7252
rect 34580 7198 34582 7250
rect 34634 7198 34916 7250
rect 34580 7196 34916 7198
rect 33404 6738 33460 6748
rect 33292 6626 33348 6636
rect 33124 5908 33180 5918
rect 32284 5906 33180 5908
rect 32284 5854 32286 5906
rect 32338 5854 33126 5906
rect 33178 5854 33180 5906
rect 32284 5852 33180 5854
rect 32284 5842 32340 5852
rect 33124 5842 33180 5852
rect 33404 5908 33460 5918
rect 33404 5814 33460 5852
rect 33516 5908 33572 5918
rect 33852 5908 33908 5918
rect 33516 5906 33908 5908
rect 33516 5854 33518 5906
rect 33570 5854 33854 5906
rect 33906 5854 33908 5906
rect 33516 5852 33908 5854
rect 32060 5730 32116 5740
rect 31724 5394 31780 5404
rect 33180 5236 33236 5246
rect 33516 5236 33572 5852
rect 33852 5842 33908 5852
rect 33180 5234 33572 5236
rect 33180 5182 33182 5234
rect 33234 5182 33572 5234
rect 33180 5180 33572 5182
rect 33180 5170 33236 5180
rect 33628 5124 33684 5134
rect 33628 5030 33684 5068
rect 31500 4834 31556 4844
rect 32508 5012 32564 5022
rect 32508 4365 32564 4956
rect 33964 5012 34020 7196
rect 34580 7186 34636 7196
rect 34188 5921 34244 5946
rect 34188 5908 34190 5921
rect 34242 5908 34244 5921
rect 34188 5842 34244 5852
rect 34748 5908 34804 5918
rect 34860 5908 34916 7196
rect 34972 7140 35028 7420
rect 35196 7410 35252 7420
rect 35420 7476 35476 7486
rect 35420 7382 35476 7420
rect 35532 7140 35588 7980
rect 35700 7476 35756 7486
rect 36204 7476 36260 7486
rect 35700 7474 36260 7476
rect 35700 7422 35702 7474
rect 35754 7422 36206 7474
rect 36258 7422 36260 7474
rect 35700 7420 36260 7422
rect 35700 7410 35756 7420
rect 36204 7410 36260 7420
rect 36316 7476 36372 8318
rect 37548 8258 37604 8652
rect 37548 8206 37550 8258
rect 37602 8206 37604 8258
rect 37548 8194 37604 8206
rect 37772 8258 37828 8270
rect 37772 8206 37774 8258
rect 37826 8206 37828 8258
rect 38108 8260 38164 8270
rect 37772 7812 37828 8206
rect 37940 8202 37996 8214
rect 37940 8150 37942 8202
rect 37994 8150 37996 8202
rect 38108 8166 38164 8204
rect 38220 8258 38276 8270
rect 38220 8206 38222 8258
rect 38274 8206 38276 8258
rect 37940 7924 37996 8150
rect 38220 8148 38276 8206
rect 38332 8260 38388 9548
rect 38444 8428 38500 10585
rect 38556 10388 38612 12910
rect 39564 12964 39620 12974
rect 39564 12870 39620 12908
rect 38836 12852 38892 12862
rect 38836 12850 39284 12852
rect 38836 12798 38838 12850
rect 38890 12798 39284 12850
rect 38836 12796 39284 12798
rect 38836 12786 38892 12796
rect 39004 12178 39060 12190
rect 39004 12126 39006 12178
rect 39058 12126 39060 12178
rect 38668 12068 38724 12078
rect 39004 12068 39060 12126
rect 38668 12066 39060 12068
rect 38668 12014 38670 12066
rect 38722 12014 39060 12066
rect 38668 12012 39060 12014
rect 39228 12178 39284 12796
rect 39228 12126 39230 12178
rect 39282 12126 39284 12178
rect 38668 11172 38724 12012
rect 39228 11732 39284 12126
rect 39788 12180 39844 12190
rect 39788 12178 39956 12180
rect 39788 12126 39790 12178
rect 39842 12126 39956 12178
rect 39788 12124 39956 12126
rect 39788 12114 39844 12124
rect 39508 11956 39564 11966
rect 39508 11862 39564 11900
rect 38668 11106 38724 11116
rect 39004 11676 39284 11732
rect 38892 10724 38948 10734
rect 38892 10388 38948 10668
rect 39004 10610 39060 11676
rect 39900 11172 39956 12124
rect 39564 11116 39956 11172
rect 39564 10778 39620 11116
rect 39564 10726 39566 10778
rect 39618 10726 39620 10778
rect 39564 10714 39620 10726
rect 39676 10724 39732 10734
rect 39004 10558 39006 10610
rect 39058 10558 39060 10610
rect 39004 10546 39060 10558
rect 39340 10637 39396 10649
rect 39340 10585 39342 10637
rect 39394 10585 39396 10637
rect 39340 10500 39396 10585
rect 39676 10610 39732 10668
rect 40012 10724 40068 14140
rect 41468 14084 41524 16843
rect 41804 16782 41860 16940
rect 42028 16884 42084 17948
rect 42140 17668 42196 17678
rect 42252 17668 42308 18172
rect 42476 18004 42532 19180
rect 43484 18686 43540 19404
rect 43428 18674 43540 18686
rect 43428 18622 43430 18674
rect 43482 18622 43540 18674
rect 43428 18620 43540 18622
rect 43428 18610 43484 18620
rect 42588 18450 42644 18462
rect 42588 18398 42590 18450
rect 42642 18398 42644 18450
rect 42588 18228 42644 18398
rect 43820 18450 43876 18462
rect 43820 18398 43822 18450
rect 43874 18398 43876 18450
rect 42588 18162 42644 18172
rect 42868 18228 42924 18238
rect 42868 18226 43204 18228
rect 42868 18174 42870 18226
rect 42922 18174 43204 18226
rect 42868 18172 43204 18174
rect 42868 18162 42924 18172
rect 42476 17948 42868 18004
rect 42812 17890 42868 17948
rect 42812 17838 42814 17890
rect 42866 17838 42868 17890
rect 42812 17826 42868 17838
rect 42140 17666 42308 17668
rect 42140 17614 42142 17666
rect 42194 17614 42308 17666
rect 42140 17612 42308 17614
rect 42140 17602 42196 17612
rect 41748 16770 41860 16782
rect 41748 16718 41750 16770
rect 41802 16718 41860 16770
rect 41748 16716 41860 16718
rect 41916 16828 42084 16884
rect 42252 16884 42308 17612
rect 43148 17666 43204 18172
rect 43820 18116 43876 18398
rect 43820 18050 43876 18060
rect 43708 18004 43764 18014
rect 43148 17614 43150 17666
rect 43202 17614 43204 17666
rect 43148 17602 43204 17614
rect 43484 17666 43540 17678
rect 43484 17614 43486 17666
rect 43538 17614 43540 17666
rect 42364 17052 42980 17108
rect 42364 16884 42420 17052
rect 42252 16882 42420 16884
rect 42252 16830 42366 16882
rect 42418 16830 42420 16882
rect 42252 16828 42420 16830
rect 41748 16706 41804 16716
rect 41804 16548 41860 16558
rect 41804 15428 41860 16492
rect 41916 15876 41972 16828
rect 42364 16818 42420 16828
rect 42476 16884 42532 16894
rect 42476 16790 42532 16828
rect 42700 16884 42756 16894
rect 42700 16790 42756 16828
rect 42924 16882 42980 17052
rect 42924 16830 42926 16882
rect 42978 16830 42980 16882
rect 42924 16818 42980 16830
rect 43484 16884 43540 17614
rect 43484 16818 43540 16828
rect 42084 16660 42140 16670
rect 43204 16660 43260 16670
rect 42084 16566 42140 16604
rect 42812 16658 43260 16660
rect 42812 16606 43206 16658
rect 43258 16606 43260 16658
rect 42812 16604 43260 16606
rect 41916 15820 42084 15876
rect 41804 15316 41860 15372
rect 41916 15316 41972 15326
rect 41804 15314 41972 15316
rect 41804 15262 41918 15314
rect 41970 15262 41972 15314
rect 41804 15260 41972 15262
rect 41916 15250 41972 15260
rect 41636 15204 41692 15242
rect 41636 15138 41692 15148
rect 42028 15148 42084 15820
rect 42364 15652 42420 15662
rect 42252 15329 42308 15354
rect 42252 15316 42254 15329
rect 42306 15316 42308 15329
rect 42252 15250 42308 15260
rect 42364 15202 42420 15596
rect 42364 15150 42366 15202
rect 42418 15150 42420 15202
rect 42028 15092 42308 15148
rect 42364 15138 42420 15150
rect 42476 15540 42532 15550
rect 41468 14018 41524 14028
rect 41692 14530 41748 14542
rect 41692 14478 41694 14530
rect 41746 14478 41748 14530
rect 40236 13972 40292 13982
rect 40236 13878 40292 13916
rect 41692 13972 41748 14478
rect 41692 13906 41748 13916
rect 41972 14084 42028 14094
rect 41972 13972 42028 14028
rect 41972 13970 42196 13972
rect 41972 13918 41974 13970
rect 42026 13918 42196 13970
rect 41972 13916 42196 13918
rect 41972 13906 42028 13916
rect 42140 13746 42196 13916
rect 42140 13694 42142 13746
rect 42194 13694 42196 13746
rect 42140 13682 42196 13694
rect 41244 13076 41300 13086
rect 40516 12964 40572 12974
rect 40516 12740 40572 12908
rect 41020 12740 41076 12750
rect 40516 12738 40740 12740
rect 40516 12686 40518 12738
rect 40570 12686 40740 12738
rect 40516 12684 40740 12686
rect 40516 12674 40572 12684
rect 40124 11954 40180 11966
rect 40124 11902 40126 11954
rect 40178 11902 40180 11954
rect 40124 11506 40180 11902
rect 40124 11454 40126 11506
rect 40178 11454 40180 11506
rect 40124 11442 40180 11454
rect 40012 10658 40068 10668
rect 39900 10612 39956 10622
rect 39676 10558 39678 10610
rect 39730 10558 39732 10610
rect 39676 10546 39732 10558
rect 39788 10610 39956 10612
rect 39788 10558 39902 10610
rect 39954 10558 39956 10610
rect 39788 10556 39956 10558
rect 39340 10434 39396 10444
rect 39228 10388 39284 10398
rect 38892 10332 39060 10388
rect 38556 10322 38612 10332
rect 38668 10164 38724 10174
rect 38668 9828 38724 10108
rect 38668 9826 38948 9828
rect 38668 9774 38670 9826
rect 38722 9774 38948 9826
rect 38668 9772 38948 9774
rect 38668 9762 38724 9772
rect 38892 9154 38948 9772
rect 38892 9102 38894 9154
rect 38946 9102 38948 9154
rect 38780 9044 38836 9054
rect 38444 8372 38724 8428
rect 38500 8260 38556 8270
rect 38332 8204 38500 8260
rect 38500 8166 38556 8204
rect 38220 8082 38276 8092
rect 38556 8036 38612 8046
rect 37940 7868 38500 7924
rect 37772 7756 38164 7812
rect 36316 7410 36372 7420
rect 36540 7476 36596 7486
rect 36540 7382 36596 7420
rect 37044 7476 37100 7486
rect 37436 7476 37492 7486
rect 37044 7362 37100 7420
rect 36092 7306 36148 7318
rect 36092 7254 36094 7306
rect 36146 7254 36148 7306
rect 34972 7074 35028 7084
rect 35196 7084 35460 7094
rect 35532 7084 35812 7140
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 34804 5852 34916 5908
rect 34972 6804 35028 6814
rect 34972 5950 35028 6748
rect 34972 5898 34974 5950
rect 35026 5898 35028 5950
rect 34972 5886 35028 5898
rect 35084 6690 35140 6702
rect 35084 6638 35086 6690
rect 35138 6638 35140 6690
rect 34748 5814 34804 5852
rect 34300 5796 34356 5806
rect 34300 5702 34356 5740
rect 35084 5794 35140 6638
rect 35756 6692 35812 7084
rect 36092 6804 36148 7254
rect 37044 7310 37046 7362
rect 37098 7310 37100 7362
rect 37044 6916 37100 7310
rect 37044 6850 37100 6860
rect 37156 7474 37492 7476
rect 37156 7422 37438 7474
rect 37490 7422 37492 7474
rect 37156 7420 37492 7422
rect 37156 6914 37212 7420
rect 37436 7410 37492 7420
rect 37156 6862 37158 6914
rect 37210 6862 37212 6914
rect 37156 6850 37212 6862
rect 37660 7028 37716 7038
rect 38108 7028 38164 7756
rect 36092 6738 36148 6748
rect 35644 5908 35700 5918
rect 35084 5742 35086 5794
rect 35138 5742 35140 5794
rect 35084 5730 35140 5742
rect 35532 5906 35700 5908
rect 35532 5854 35646 5906
rect 35698 5854 35700 5906
rect 35532 5852 35700 5854
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 33964 4946 34020 4956
rect 34412 5122 34468 5134
rect 34412 5070 34414 5122
rect 34466 5070 34468 5122
rect 34412 4564 34468 5070
rect 35084 4900 35140 4910
rect 35532 4900 35588 5852
rect 35644 5842 35700 5852
rect 34412 4508 35028 4564
rect 32508 4313 32510 4365
rect 32562 4313 32564 4365
rect 32508 4301 32564 4313
rect 33180 4340 33236 4350
rect 33180 4246 33236 4284
rect 34636 4004 34692 4014
rect 33404 3668 33460 3678
rect 31388 3502 31390 3554
rect 31442 3502 31444 3554
rect 31388 3490 31444 3502
rect 31612 3556 31668 3566
rect 30492 3475 30548 3487
rect 27748 3322 27804 3334
rect 28420 3332 28476 3342
rect 28028 3330 28476 3332
rect 26236 2940 26628 2996
rect 28028 3278 28422 3330
rect 28474 3278 28476 3330
rect 29036 3334 29038 3386
rect 29090 3334 29092 3386
rect 29036 3322 29092 3334
rect 29820 3444 29876 3454
rect 28028 3276 28476 3278
rect 23940 2718 23942 2770
rect 23994 2718 23996 2770
rect 23940 2706 23996 2718
rect 24444 2770 24500 2782
rect 24444 2718 24446 2770
rect 24498 2718 24500 2770
rect 24444 800 24500 2718
rect 26236 800 26292 2940
rect 28028 800 28084 3276
rect 28420 3266 28476 3276
rect 29820 800 29876 3388
rect 31612 800 31668 3500
rect 32396 3556 32452 3566
rect 32396 3462 32452 3500
rect 33404 800 33460 3612
rect 34636 3526 34692 3948
rect 34972 3722 35028 4508
rect 35084 4338 35140 4844
rect 35084 4286 35086 4338
rect 35138 4286 35140 4338
rect 35084 4274 35140 4286
rect 35196 4844 35588 4900
rect 35644 5236 35700 5246
rect 35756 5236 35812 6636
rect 35700 5180 35812 5236
rect 35868 6690 35924 6702
rect 36540 6692 36596 6702
rect 35868 6638 35870 6690
rect 35922 6638 35924 6690
rect 35196 4116 35252 4844
rect 35084 4060 35252 4116
rect 35084 3780 35140 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 35644 3780 35700 5180
rect 35868 5124 35924 6638
rect 36316 6690 36596 6692
rect 36316 6638 36542 6690
rect 36594 6638 36596 6690
rect 36316 6636 36596 6638
rect 35868 4340 35924 5068
rect 36204 6466 36260 6478
rect 36204 6414 36206 6466
rect 36258 6414 36260 6466
rect 35980 4340 36036 4350
rect 35868 4338 36036 4340
rect 35868 4286 35870 4338
rect 35922 4286 35982 4338
rect 36034 4286 36036 4338
rect 35868 4284 36036 4286
rect 35868 4274 35924 4284
rect 35980 4274 36036 4284
rect 35084 3724 35252 3780
rect 34972 3670 34974 3722
rect 35026 3670 35028 3722
rect 34972 3658 35028 3670
rect 34636 3474 34638 3526
rect 34690 3474 34692 3526
rect 34636 3462 34692 3474
rect 35084 3556 35140 3566
rect 35084 3462 35140 3500
rect 35196 800 35252 3724
rect 35420 3724 35700 3780
rect 35420 3554 35476 3724
rect 35420 3502 35422 3554
rect 35474 3502 35476 3554
rect 35420 3490 35476 3502
rect 36204 3526 36260 6414
rect 36316 5234 36372 6636
rect 36540 6626 36596 6636
rect 37324 6692 37380 6702
rect 37548 6692 37604 6702
rect 37324 6690 37548 6692
rect 37324 6638 37326 6690
rect 37378 6638 37548 6690
rect 37324 6636 37548 6638
rect 37324 6626 37380 6636
rect 37548 6598 37604 6636
rect 37660 6690 37716 6972
rect 37940 6972 38164 7028
rect 38312 7700 38368 7710
rect 38312 7474 38368 7644
rect 38312 7422 38314 7474
rect 38366 7422 38368 7474
rect 38312 7028 38368 7422
rect 37940 6914 37996 6972
rect 38312 6962 38368 6972
rect 37940 6862 37942 6914
rect 37994 6862 37996 6914
rect 37940 6850 37996 6862
rect 37660 6638 37662 6690
rect 37714 6638 37716 6690
rect 37660 6626 37716 6638
rect 37436 6468 37492 6478
rect 36316 5182 36318 5234
rect 36370 5182 36372 5234
rect 36316 5170 36372 5182
rect 37156 5236 37212 5246
rect 37156 5142 37212 5180
rect 37436 5122 37492 6412
rect 37884 5933 37940 5945
rect 37884 5881 37886 5933
rect 37938 5881 37940 5933
rect 37884 5236 37940 5881
rect 38108 5236 38164 5246
rect 37884 5180 38052 5236
rect 37436 5070 37438 5122
rect 37490 5070 37492 5122
rect 37436 5058 37492 5070
rect 37884 5066 37940 5078
rect 37884 5014 37886 5066
rect 37938 5014 37940 5066
rect 36764 4340 36820 4350
rect 36764 4246 36820 4284
rect 37884 4228 37940 5014
rect 37884 4162 37940 4172
rect 36988 3668 37044 3678
rect 36988 3574 37044 3612
rect 37996 3668 38052 5180
rect 38108 5122 38164 5180
rect 38108 5070 38110 5122
rect 38162 5070 38164 5122
rect 38108 5058 38164 5070
rect 38444 5124 38500 7868
rect 38556 7586 38612 7980
rect 38556 7534 38558 7586
rect 38610 7534 38612 7586
rect 38556 7140 38612 7534
rect 38668 7364 38724 8372
rect 38668 7298 38724 7308
rect 38556 7084 38724 7140
rect 38556 6692 38612 6702
rect 38556 6598 38612 6636
rect 38668 6020 38724 7084
rect 38556 5964 38724 6020
rect 38556 5962 38612 5964
rect 38556 5910 38558 5962
rect 38610 5910 38612 5962
rect 38556 5898 38612 5910
rect 38220 4954 38276 4966
rect 38220 4902 38222 4954
rect 38274 4902 38276 4954
rect 38220 4676 38276 4902
rect 38444 4900 38500 5068
rect 38556 5684 38612 5694
rect 38556 5122 38612 5628
rect 38556 5070 38558 5122
rect 38610 5070 38612 5122
rect 38556 5058 38612 5070
rect 38444 4844 38724 4900
rect 38220 4610 38276 4620
rect 38668 4450 38724 4844
rect 38668 4398 38670 4450
rect 38722 4398 38724 4450
rect 38668 4386 38724 4398
rect 38780 4228 38836 8988
rect 38892 8258 38948 9102
rect 39004 9826 39060 10332
rect 39004 9774 39006 9826
rect 39058 9774 39060 9826
rect 39004 9492 39060 9774
rect 39004 8484 39060 9436
rect 39116 9658 39172 9670
rect 39116 9606 39118 9658
rect 39170 9606 39172 9658
rect 39116 8708 39172 9606
rect 39116 8642 39172 8652
rect 39228 8494 39284 10332
rect 39340 10276 39396 10286
rect 39340 9799 39396 10220
rect 39340 9747 39342 9799
rect 39394 9747 39396 9799
rect 39676 10164 39732 10174
rect 39676 9826 39732 10108
rect 39676 9774 39678 9826
rect 39730 9774 39732 9826
rect 39676 9762 39732 9774
rect 39340 9735 39396 9747
rect 39788 9604 39844 10556
rect 39900 10546 39956 10556
rect 40236 10388 40292 10398
rect 40124 10386 40292 10388
rect 40124 10334 40238 10386
rect 40290 10334 40292 10386
rect 40124 10332 40292 10334
rect 39508 9548 39844 9604
rect 40012 9716 40068 9726
rect 39508 9154 39564 9548
rect 39508 9102 39510 9154
rect 39562 9102 39564 9154
rect 39508 9090 39564 9102
rect 40012 9054 40068 9660
rect 40124 9268 40180 10332
rect 40236 10322 40292 10332
rect 40684 10052 40740 12684
rect 41020 12646 41076 12684
rect 41244 12068 41300 13020
rect 41356 12962 41412 12974
rect 41356 12910 41358 12962
rect 41410 12910 41412 12962
rect 41356 12852 41412 12910
rect 41356 12786 41412 12796
rect 41692 12962 41748 12974
rect 41692 12910 41694 12962
rect 41746 12910 41748 12962
rect 41692 12740 41748 12910
rect 41916 12964 41972 12974
rect 41916 12895 41918 12908
rect 41970 12895 41972 12908
rect 42252 12962 42308 15092
rect 42252 12910 42254 12962
rect 42306 12910 42308 12962
rect 42252 12898 42308 12910
rect 42364 14980 42420 14990
rect 42364 13524 42420 14924
rect 42476 14530 42532 15484
rect 42700 15316 42756 15326
rect 42700 15146 42756 15260
rect 42812 15314 42868 16604
rect 43204 16594 43260 16604
rect 43260 16436 43316 16446
rect 43036 16098 43092 16110
rect 43036 16046 43038 16098
rect 43090 16046 43092 16098
rect 43036 15652 43092 16046
rect 43036 15586 43092 15596
rect 42812 15262 42814 15314
rect 42866 15262 42868 15314
rect 42812 15250 42868 15262
rect 42924 15540 42980 15550
rect 42700 15094 42702 15146
rect 42754 15094 42756 15146
rect 42700 15082 42756 15094
rect 42812 15092 42868 15102
rect 42812 14766 42868 15036
rect 42756 14754 42868 14766
rect 42756 14702 42758 14754
rect 42810 14702 42868 14754
rect 42756 14700 42868 14702
rect 42756 14690 42812 14700
rect 42476 14478 42478 14530
rect 42530 14478 42532 14530
rect 42476 14466 42532 14478
rect 42924 13746 42980 15484
rect 43148 15428 43204 15438
rect 43036 15314 43092 15326
rect 43036 15262 43038 15314
rect 43090 15262 43092 15314
rect 43036 14980 43092 15262
rect 43036 14914 43092 14924
rect 43036 14532 43092 14542
rect 43148 14532 43204 15372
rect 43036 14530 43204 14532
rect 43036 14478 43038 14530
rect 43090 14478 43204 14530
rect 43036 14476 43204 14478
rect 43260 14530 43316 16380
rect 43708 16212 43764 17948
rect 43932 17778 43988 19964
rect 44044 19954 44100 19964
rect 44156 20018 44212 20030
rect 44156 19966 44158 20018
rect 44210 19966 44212 20018
rect 44156 19348 44212 19966
rect 44322 20020 44378 20030
rect 44322 19926 44378 19964
rect 44996 19908 45052 19918
rect 44716 19794 44772 19806
rect 44716 19742 44718 19794
rect 44770 19742 44772 19794
rect 44716 19684 44772 19742
rect 44716 19618 44772 19628
rect 44044 19292 44212 19348
rect 44044 18618 44100 19292
rect 44044 18566 44046 18618
rect 44098 18566 44100 18618
rect 44044 18554 44100 18566
rect 44156 19122 44212 19134
rect 44156 19070 44158 19122
rect 44210 19070 44212 19122
rect 44044 18465 44100 18477
rect 44044 18413 44046 18465
rect 44098 18452 44100 18465
rect 44156 18452 44212 19070
rect 44996 19012 45052 19852
rect 45444 19460 45500 19470
rect 45444 19346 45500 19404
rect 45948 19358 46004 20076
rect 45444 19294 45446 19346
rect 45498 19294 45500 19346
rect 45444 19282 45500 19294
rect 45892 19346 46004 19358
rect 45892 19294 45894 19346
rect 45946 19294 46004 19346
rect 45892 19292 46004 19294
rect 45892 19282 45948 19292
rect 46172 19012 46228 20524
rect 46396 20524 46788 20580
rect 46396 20018 46452 20524
rect 46844 20468 46900 21534
rect 47348 21476 47404 21486
rect 47348 21382 47404 21420
rect 47628 21474 47684 22652
rect 47628 21422 47630 21474
rect 47682 21422 47684 21474
rect 47628 21410 47684 21422
rect 47740 21601 47796 21613
rect 47740 21549 47742 21601
rect 47794 21549 47796 21601
rect 47740 21476 47796 21549
rect 47740 21410 47796 21420
rect 47852 21588 47908 21598
rect 46396 19966 46398 20018
rect 46450 19966 46452 20018
rect 46396 19954 46452 19966
rect 46620 20356 46676 20366
rect 46620 19906 46676 20300
rect 46732 20064 46788 20074
rect 46844 20064 46900 20412
rect 46956 20802 47012 20814
rect 47740 20804 47796 20814
rect 46956 20750 46958 20802
rect 47010 20750 47012 20802
rect 46956 20244 47012 20750
rect 46956 20178 47012 20188
rect 47292 20748 47740 20804
rect 47852 20804 47908 21532
rect 48076 21586 48132 23214
rect 48076 21534 48078 21586
rect 48130 21534 48132 21586
rect 48076 21522 48132 21534
rect 48524 21476 48580 23660
rect 48636 23156 48692 23166
rect 48636 23062 48692 23100
rect 47964 20804 48020 20814
rect 47852 20802 48020 20804
rect 47852 20750 47966 20802
rect 48018 20750 48020 20802
rect 48524 20804 48580 21420
rect 48636 21586 48692 21598
rect 48636 21534 48638 21586
rect 48690 21534 48692 21586
rect 48636 21364 48692 21534
rect 48636 21298 48692 21308
rect 48636 20804 48692 20814
rect 48524 20802 48692 20804
rect 47852 20748 48020 20750
rect 46732 20062 46900 20064
rect 46732 20010 46734 20062
rect 46786 20010 46900 20062
rect 46732 20008 46900 20010
rect 47068 20020 47124 20030
rect 46732 19998 46788 20008
rect 47068 19926 47124 19964
rect 47292 20018 47348 20748
rect 47740 20710 47796 20748
rect 47964 20738 48020 20748
rect 48300 20746 48356 20758
rect 48300 20694 48302 20746
rect 48354 20694 48356 20746
rect 47292 19966 47294 20018
rect 47346 19966 47348 20018
rect 46620 19854 46622 19906
rect 46674 19854 46676 19906
rect 46620 19842 46676 19854
rect 46956 19796 47012 19806
rect 46396 19236 46452 19246
rect 46396 19142 46452 19180
rect 44996 19010 45220 19012
rect 44996 18958 44998 19010
rect 45050 18958 45220 19010
rect 44996 18956 45220 18958
rect 46172 18956 46788 19012
rect 44996 18946 45052 18956
rect 44492 18452 44548 18462
rect 44098 18450 44548 18452
rect 44098 18413 44494 18450
rect 44044 18398 44494 18413
rect 44546 18398 44548 18450
rect 44044 18396 44548 18398
rect 44492 18386 44548 18396
rect 43932 17726 43934 17778
rect 43986 17726 43988 17778
rect 43932 17714 43988 17726
rect 44044 18116 44100 18126
rect 43820 17668 43876 17678
rect 43820 17599 43822 17612
rect 43874 17599 43876 17612
rect 43820 17574 43876 17599
rect 44044 16882 44100 18060
rect 45164 18004 45220 18956
rect 45368 18452 45424 18462
rect 45948 18452 46004 18462
rect 45368 18450 46004 18452
rect 45368 18398 45370 18450
rect 45422 18398 45950 18450
rect 46002 18398 46004 18450
rect 45368 18396 46004 18398
rect 45368 18386 45424 18396
rect 45052 17948 45220 18004
rect 44044 16830 44046 16882
rect 44098 16830 44100 16882
rect 44044 16436 44100 16830
rect 44268 16884 44324 16894
rect 44268 16790 44324 16828
rect 44548 16884 44604 16894
rect 44548 16790 44604 16828
rect 44044 16370 44100 16380
rect 44940 16436 44996 16446
rect 43260 14478 43262 14530
rect 43314 14478 43316 14530
rect 43036 14466 43092 14476
rect 43260 14466 43316 14478
rect 43372 15540 43428 15550
rect 43372 14530 43428 15484
rect 43484 15316 43540 15326
rect 43484 14980 43540 15260
rect 43708 15148 43764 16156
rect 44212 16212 44268 16222
rect 44212 16118 44268 16156
rect 44940 16210 44996 16380
rect 44940 16158 44942 16210
rect 44994 16158 44996 16210
rect 44940 16146 44996 16158
rect 43820 16098 43876 16110
rect 43820 16046 43822 16098
rect 43874 16046 43876 16098
rect 43820 15540 43876 16046
rect 43820 15474 43876 15484
rect 44716 15540 44772 15550
rect 44716 15446 44772 15484
rect 43708 15092 43988 15148
rect 43484 14914 43540 14924
rect 43372 14478 43374 14530
rect 43426 14478 43428 14530
rect 43372 14466 43428 14478
rect 42924 13694 42926 13746
rect 42978 13694 42980 13746
rect 42476 13524 42532 13534
rect 42364 13522 42532 13524
rect 42364 13470 42478 13522
rect 42530 13470 42532 13522
rect 42364 13468 42532 13470
rect 41916 12870 41972 12895
rect 41692 12674 41748 12684
rect 41916 12794 41972 12806
rect 41916 12742 41918 12794
rect 41970 12742 41972 12794
rect 41916 12180 41972 12742
rect 41916 12114 41972 12124
rect 42028 12178 42084 12190
rect 42028 12126 42030 12178
rect 42082 12126 42084 12178
rect 41412 12068 41468 12078
rect 41244 12012 41412 12068
rect 41412 11974 41468 12012
rect 41748 11956 41804 11966
rect 41692 11954 41804 11956
rect 41692 11902 41750 11954
rect 41802 11902 41804 11954
rect 41692 11890 41804 11902
rect 41020 11732 41076 11742
rect 40908 11396 40964 11406
rect 41020 11396 41076 11676
rect 40908 11394 41076 11396
rect 40908 11342 40910 11394
rect 40962 11342 41022 11394
rect 41074 11342 41076 11394
rect 40908 11340 41076 11342
rect 40908 11330 40964 11340
rect 41020 11330 41076 11340
rect 41020 10625 41076 10637
rect 41020 10573 41022 10625
rect 41074 10573 41076 10625
rect 40908 10500 40964 10510
rect 40908 10406 40964 10444
rect 41020 10164 41076 10573
rect 41244 10612 41300 10622
rect 41244 10518 41300 10556
rect 41580 10500 41636 10510
rect 41020 10098 41076 10108
rect 41468 10498 41636 10500
rect 41468 10446 41582 10498
rect 41634 10446 41636 10498
rect 41468 10444 41636 10446
rect 40684 9996 40908 10052
rect 40292 9940 40348 9950
rect 40292 9846 40348 9884
rect 40124 9202 40180 9212
rect 40572 9826 40628 9838
rect 40572 9774 40574 9826
rect 40626 9774 40628 9826
rect 40572 9156 40628 9774
rect 40852 9770 40908 9996
rect 41468 10050 41524 10444
rect 41580 10434 41636 10444
rect 41468 9998 41470 10050
rect 41522 9998 41524 10050
rect 41468 9986 41524 9998
rect 40684 9714 40740 9726
rect 40684 9662 40686 9714
rect 40738 9662 40740 9714
rect 40684 9492 40740 9662
rect 40852 9718 40854 9770
rect 40906 9718 40908 9770
rect 41020 9828 41076 9838
rect 41692 9828 41748 11890
rect 41804 11394 41860 11406
rect 41804 11342 41806 11394
rect 41858 11342 41860 11394
rect 41804 10498 41860 11342
rect 42028 10836 42084 12126
rect 42140 12178 42196 12190
rect 42140 12126 42142 12178
rect 42194 12126 42196 12178
rect 42140 12068 42196 12126
rect 42140 12002 42196 12012
rect 42364 11844 42420 13468
rect 42476 13458 42532 13468
rect 42588 13524 42644 13534
rect 42476 12964 42532 12974
rect 42588 12964 42644 13468
rect 42476 12962 42644 12964
rect 42476 12910 42478 12962
rect 42530 12910 42644 12962
rect 42476 12908 42644 12910
rect 42476 12898 42532 12908
rect 42756 12852 42812 12862
rect 42756 12758 42812 12796
rect 42588 12292 42644 12302
rect 42588 12222 42644 12236
rect 42588 12170 42590 12222
rect 42642 12170 42644 12222
rect 42588 12158 42644 12170
rect 42812 12178 42868 12190
rect 42812 12126 42814 12178
rect 42866 12126 42868 12178
rect 42364 11778 42420 11788
rect 42476 12066 42532 12078
rect 42476 12014 42478 12066
rect 42530 12014 42532 12066
rect 42476 11732 42532 12014
rect 42812 11956 42868 12126
rect 42924 12180 42980 13694
rect 43708 13636 43764 13646
rect 43708 13634 43876 13636
rect 43708 13582 43710 13634
rect 43762 13582 43876 13634
rect 43708 13580 43876 13582
rect 43708 13570 43764 13580
rect 43596 13524 43652 13534
rect 43596 12962 43652 13468
rect 43820 13074 43876 13580
rect 43932 13300 43988 15092
rect 44828 14420 44884 14430
rect 44828 13748 44884 14364
rect 43932 13244 44100 13300
rect 43820 13022 43822 13074
rect 43874 13022 43876 13074
rect 43820 13010 43876 13022
rect 43932 13076 43988 13086
rect 43596 12910 43598 12962
rect 43650 12910 43652 12962
rect 43596 12898 43652 12910
rect 43932 12947 43988 13020
rect 43932 12895 43934 12947
rect 43986 12895 43988 12947
rect 43932 12883 43988 12895
rect 43820 12852 43876 12862
rect 43260 12738 43316 12750
rect 43260 12686 43262 12738
rect 43314 12686 43316 12738
rect 43260 12292 43316 12686
rect 43148 12180 43204 12190
rect 42924 12178 43204 12180
rect 42924 12126 43150 12178
rect 43202 12126 43204 12178
rect 42924 12124 43204 12126
rect 43148 12114 43204 12124
rect 43260 11956 43316 12236
rect 42812 11890 42868 11900
rect 43148 11900 43316 11956
rect 43372 11956 43428 11966
rect 42476 11676 43092 11732
rect 42476 11172 42532 11182
rect 42028 10780 42196 10836
rect 42140 10622 42196 10780
rect 42122 10610 42196 10622
rect 42122 10558 42124 10610
rect 42176 10558 42196 10610
rect 42122 10556 42196 10558
rect 42364 10612 42420 10622
rect 42122 10546 42178 10556
rect 42364 10518 42420 10556
rect 41804 10446 41806 10498
rect 41858 10446 41860 10498
rect 41804 10434 41860 10446
rect 41916 9940 41972 9950
rect 41804 9828 41860 9838
rect 41692 9826 41860 9828
rect 41692 9774 41806 9826
rect 41858 9774 41860 9826
rect 41692 9772 41860 9774
rect 41020 9734 41076 9772
rect 41804 9762 41860 9772
rect 41916 9826 41972 9884
rect 41916 9774 41918 9826
rect 41970 9774 41972 9826
rect 41916 9762 41972 9774
rect 40852 9716 40908 9718
rect 40852 9650 40908 9660
rect 41580 9604 41636 9614
rect 40684 9436 41412 9492
rect 40572 9090 40628 9100
rect 41132 9268 41188 9278
rect 39788 9044 39844 9054
rect 39788 8950 39844 8988
rect 39900 9042 39956 9054
rect 39900 8990 39902 9042
rect 39954 8990 39956 9042
rect 39004 8428 39172 8484
rect 39228 8482 39340 8494
rect 39228 8430 39286 8482
rect 39338 8430 39340 8482
rect 39228 8428 39340 8430
rect 38892 8206 38894 8258
rect 38946 8206 38948 8258
rect 38892 8194 38948 8206
rect 39004 8260 39060 8270
rect 39004 8166 39060 8204
rect 39116 8036 39172 8428
rect 39284 8418 39340 8428
rect 39004 7980 39172 8036
rect 39564 8258 39620 8270
rect 39564 8206 39566 8258
rect 39618 8206 39620 8258
rect 37996 3602 38052 3612
rect 38668 4172 38836 4228
rect 38892 7140 38948 7150
rect 38892 5906 38948 7084
rect 39004 6468 39060 7980
rect 39452 7476 39508 7486
rect 39340 7474 39508 7476
rect 39340 7422 39454 7474
rect 39506 7422 39508 7474
rect 39340 7420 39508 7422
rect 39172 7364 39228 7374
rect 39172 7270 39228 7308
rect 39228 6916 39284 6926
rect 39004 6402 39060 6412
rect 39116 6804 39172 6814
rect 39116 6018 39172 6748
rect 39116 5966 39118 6018
rect 39170 5966 39172 6018
rect 39116 5954 39172 5966
rect 39228 6020 39284 6860
rect 39340 6692 39396 7420
rect 39452 7410 39508 7420
rect 39564 7140 39620 8206
rect 39788 8258 39844 8270
rect 39788 8206 39790 8258
rect 39842 8206 39844 8258
rect 39788 8148 39844 8206
rect 39788 8082 39844 8092
rect 39900 7252 39956 8990
rect 40012 9042 40124 9054
rect 40012 8990 40070 9042
rect 40122 8990 40124 9042
rect 40012 8988 40124 8990
rect 40068 8978 40124 8988
rect 40236 9044 40292 9054
rect 40236 8950 40292 8988
rect 40796 9042 40852 9054
rect 40796 8990 40798 9042
rect 40850 8990 40852 9042
rect 40348 8258 40404 8270
rect 40348 8206 40350 8258
rect 40402 8206 40404 8258
rect 40068 8148 40124 8158
rect 40068 8146 40292 8148
rect 40068 8094 40070 8146
rect 40122 8094 40292 8146
rect 40068 8092 40292 8094
rect 40068 8082 40124 8092
rect 39900 7186 39956 7196
rect 39564 7074 39620 7084
rect 39340 6468 39396 6636
rect 40236 6468 40292 8092
rect 40348 7476 40404 8206
rect 40796 7476 40852 8990
rect 41132 8370 41188 9212
rect 41132 8318 41134 8370
rect 41186 8318 41188 8370
rect 41132 8306 41188 8318
rect 41132 7476 41188 7486
rect 40348 7474 41188 7476
rect 40348 7422 41134 7474
rect 41186 7422 41188 7474
rect 40348 7420 41188 7422
rect 40348 6692 40404 7420
rect 41132 7410 41188 7420
rect 41244 7252 41300 7262
rect 41244 6916 41300 7196
rect 41356 7028 41412 9436
rect 41580 9042 41636 9548
rect 42252 9604 42308 9614
rect 42252 9510 42308 9548
rect 42476 9604 42532 11116
rect 43036 10722 43092 11676
rect 43036 10670 43038 10722
rect 43090 10670 43092 10722
rect 43036 10658 43092 10670
rect 42868 10554 42924 10566
rect 42868 10502 42870 10554
rect 42922 10502 42924 10554
rect 42868 10052 42924 10502
rect 42868 9986 42924 9996
rect 42476 9538 42532 9548
rect 42868 9602 42924 9614
rect 42868 9550 42870 9602
rect 42922 9550 42924 9602
rect 42868 9492 42924 9550
rect 42868 9426 42924 9436
rect 43148 9156 43204 11900
rect 43372 10610 43428 11900
rect 43820 11844 43876 12796
rect 43932 12180 43988 12190
rect 43932 12086 43988 12124
rect 43372 10558 43374 10610
rect 43426 10558 43428 10610
rect 43372 10546 43428 10558
rect 43708 11282 43764 11294
rect 43708 11230 43710 11282
rect 43762 11230 43764 11282
rect 43708 10612 43764 11230
rect 43820 10612 43876 11788
rect 44044 11172 44100 13244
rect 44268 12962 44324 12974
rect 44268 12910 44270 12962
rect 44322 12910 44324 12962
rect 44268 12852 44324 12910
rect 44828 12852 44884 13692
rect 44940 14418 44996 14430
rect 44940 14366 44942 14418
rect 44994 14366 44996 14418
rect 44940 13076 44996 14366
rect 44940 13010 44996 13020
rect 44940 12906 44996 12918
rect 44940 12854 44942 12906
rect 44994 12854 44996 12906
rect 44940 12852 44996 12854
rect 44828 12796 44996 12852
rect 44268 12786 44324 12796
rect 44604 11844 44660 11854
rect 44324 11172 44380 11182
rect 44044 11170 44436 11172
rect 44044 11118 44326 11170
rect 44378 11118 44436 11170
rect 44044 11116 44436 11118
rect 44324 11106 44436 11116
rect 43932 10612 43988 10622
rect 43820 10610 43988 10612
rect 43820 10558 43934 10610
rect 43986 10558 43988 10610
rect 43820 10556 43988 10558
rect 43708 10164 43764 10556
rect 43932 10546 43988 10556
rect 44380 10612 44436 11106
rect 44604 10654 44660 11788
rect 44940 11844 44996 11854
rect 44604 10602 44606 10654
rect 44658 10602 44660 10654
rect 44604 10590 44660 10602
rect 44716 11732 44772 11742
rect 44716 11394 44772 11676
rect 44716 11342 44718 11394
rect 44770 11342 44772 11394
rect 43484 10108 43764 10164
rect 44156 10442 44212 10454
rect 44156 10390 44158 10442
rect 44210 10390 44212 10442
rect 43316 9828 43372 9838
rect 43316 9734 43372 9772
rect 43148 9090 43204 9100
rect 43260 9604 43316 9614
rect 43484 9604 43540 10108
rect 44156 9940 44212 10390
rect 44156 9874 44212 9884
rect 41580 8990 41582 9042
rect 41634 8990 41636 9042
rect 41580 8978 41636 8990
rect 43036 8372 43092 8382
rect 43092 8316 43204 8372
rect 43036 8278 43092 8316
rect 43036 7501 43092 7513
rect 43036 7449 43038 7501
rect 43090 7449 43092 7501
rect 43036 7364 43092 7449
rect 43036 7298 43092 7308
rect 41356 6972 41748 7028
rect 41244 6860 41524 6916
rect 40460 6804 40516 6814
rect 40460 6710 40516 6748
rect 41244 6692 41300 6702
rect 40348 6626 40404 6636
rect 40908 6636 41244 6692
rect 39340 6412 39508 6468
rect 39228 5954 39284 5964
rect 38892 5854 38894 5906
rect 38946 5854 38948 5906
rect 38892 5236 38948 5854
rect 39284 5850 39340 5862
rect 39284 5798 39286 5850
rect 39338 5798 39340 5850
rect 39284 5460 39340 5798
rect 39452 5684 39508 6412
rect 39676 6412 40292 6468
rect 39676 5906 39732 6412
rect 39676 5854 39678 5906
rect 39730 5854 39732 5906
rect 39676 5842 39732 5854
rect 39900 6020 39956 6030
rect 39900 5906 39956 5964
rect 39900 5854 39902 5906
rect 39954 5854 39956 5906
rect 39900 5842 39956 5854
rect 40908 5906 40964 6636
rect 41244 6598 41300 6636
rect 41356 6690 41412 6702
rect 41356 6638 41358 6690
rect 41410 6638 41412 6690
rect 41356 6580 41412 6638
rect 41356 6514 41412 6524
rect 40908 5854 40910 5906
rect 40962 5854 40964 5906
rect 40908 5842 40964 5854
rect 39452 5618 39508 5628
rect 39564 5738 39620 5750
rect 39564 5686 39566 5738
rect 39618 5686 39620 5738
rect 39564 5460 39620 5686
rect 39284 5404 39620 5460
rect 41356 5684 41412 5694
rect 36204 3474 36206 3526
rect 36258 3474 36260 3526
rect 38668 3556 38724 4172
rect 38892 3790 38948 5180
rect 39340 5236 39396 5246
rect 39340 5142 39396 5180
rect 39452 5124 39508 5134
rect 38836 3778 38948 3790
rect 38836 3726 38838 3778
rect 38890 3726 38948 3778
rect 38836 3724 38948 3726
rect 39004 4900 39060 4910
rect 38836 3714 38892 3724
rect 38668 3490 38724 3500
rect 36204 3462 36260 3474
rect 36988 3444 37044 3454
rect 36988 800 37044 3388
rect 39004 2548 39060 4844
rect 39228 4452 39284 4462
rect 39228 4382 39284 4396
rect 39228 4330 39230 4382
rect 39282 4330 39284 4382
rect 39116 4228 39172 4238
rect 39116 4134 39172 4172
rect 39116 3556 39172 3566
rect 39228 3556 39284 4330
rect 39452 4338 39508 5068
rect 41244 5124 41300 5134
rect 41244 5030 41300 5068
rect 39452 4286 39454 4338
rect 39506 4286 39508 4338
rect 39116 3554 39284 3556
rect 39116 3502 39118 3554
rect 39170 3502 39284 3554
rect 39116 3500 39284 3502
rect 39340 3556 39396 3566
rect 39452 3556 39508 4286
rect 39788 4676 39844 4686
rect 39788 4338 39844 4620
rect 40964 4506 41020 4518
rect 40964 4454 40966 4506
rect 41018 4454 41020 4506
rect 39788 4286 39790 4338
rect 39842 4286 39844 4338
rect 39788 4274 39844 4286
rect 40124 4340 40180 4350
rect 40124 4246 40180 4284
rect 40964 4004 41020 4454
rect 41356 4338 41412 5628
rect 41468 5348 41524 6860
rect 41580 5684 41636 6972
rect 41692 6690 41748 6972
rect 41692 6638 41694 6690
rect 41746 6638 41748 6690
rect 41692 6626 41748 6638
rect 42588 6690 42644 6702
rect 42588 6638 42590 6690
rect 42642 6638 42644 6690
rect 42252 6468 42308 6478
rect 42028 6466 42308 6468
rect 42028 6414 42254 6466
rect 42306 6414 42308 6466
rect 42028 6412 42308 6414
rect 42028 6132 42084 6412
rect 42252 6402 42308 6412
rect 42588 6244 42644 6638
rect 43148 6662 43204 8316
rect 43260 6916 43316 9548
rect 43372 9548 43540 9604
rect 43596 9826 43652 9838
rect 43596 9774 43598 9826
rect 43650 9774 43652 9826
rect 43372 8932 43428 9548
rect 43484 9156 43540 9166
rect 43484 9062 43540 9100
rect 43372 8876 43540 8932
rect 43372 8260 43428 8270
rect 43372 8166 43428 8204
rect 43484 7476 43540 8876
rect 43596 8260 43652 9774
rect 43820 9826 43876 9838
rect 43820 9774 43822 9826
rect 43874 9774 43876 9826
rect 43820 9156 43876 9774
rect 43820 9090 43876 9100
rect 44156 9716 44212 9726
rect 44156 9614 44212 9660
rect 44156 9602 44268 9614
rect 44156 9550 44214 9602
rect 44266 9550 44268 9602
rect 44156 9538 44268 9550
rect 43988 9044 44044 9054
rect 43988 8950 44044 8988
rect 43596 8194 43652 8204
rect 43820 8484 43876 8494
rect 43708 8034 43764 8046
rect 43708 7982 43710 8034
rect 43762 7982 43764 8034
rect 43708 7588 43764 7982
rect 43708 7522 43764 7532
rect 43596 7476 43652 7486
rect 43484 7474 43652 7476
rect 43484 7422 43598 7474
rect 43650 7422 43652 7474
rect 43484 7420 43652 7422
rect 43596 7410 43652 7420
rect 43820 7364 43876 8428
rect 44156 8372 44212 9538
rect 44268 9156 44324 9166
rect 44268 9098 44324 9100
rect 44268 9046 44270 9098
rect 44322 9046 44324 9098
rect 44268 9034 44324 9046
rect 44380 8932 44436 10556
rect 44492 10500 44548 10510
rect 44492 9070 44548 10444
rect 44716 10388 44772 11342
rect 44940 10610 44996 11788
rect 44940 10558 44942 10610
rect 44994 10558 44996 10610
rect 44940 10546 44996 10558
rect 44716 10322 44772 10332
rect 44492 9018 44494 9070
rect 44546 9044 44548 9070
rect 44716 9940 44772 9950
rect 44716 9070 44772 9884
rect 45052 9828 45108 17948
rect 45500 17834 45556 18396
rect 45948 18386 46004 18396
rect 46172 18452 46228 18462
rect 46452 18452 46508 18462
rect 46172 18450 46340 18452
rect 46172 18398 46174 18450
rect 46226 18398 46340 18450
rect 46172 18396 46340 18398
rect 46172 18386 46228 18396
rect 45612 18228 45668 18238
rect 45612 18134 45668 18172
rect 45500 17782 45502 17834
rect 45554 17782 45556 17834
rect 45500 17770 45556 17782
rect 45276 17668 45332 17678
rect 45500 17668 45556 17678
rect 45164 17612 45276 17668
rect 45164 16882 45220 17612
rect 45276 17574 45332 17612
rect 45388 17666 45556 17668
rect 45388 17614 45502 17666
rect 45554 17614 45556 17666
rect 45388 17612 45556 17614
rect 45164 16830 45166 16882
rect 45218 16830 45220 16882
rect 45164 16818 45220 16830
rect 45276 16884 45332 16894
rect 45388 16884 45444 17612
rect 45500 17602 45556 17612
rect 45948 17444 46004 17454
rect 46116 17444 46172 17454
rect 46004 17442 46172 17444
rect 46004 17390 46118 17442
rect 46170 17390 46172 17442
rect 46004 17388 46172 17390
rect 45332 16828 45444 16884
rect 45556 16884 45612 16894
rect 45556 16882 45892 16884
rect 45556 16830 45558 16882
rect 45610 16830 45892 16882
rect 45556 16828 45892 16830
rect 45276 16790 45332 16828
rect 45556 16818 45612 16828
rect 45836 16660 45892 16828
rect 45948 16882 46004 17388
rect 46116 17378 46172 17388
rect 46284 17006 46340 18396
rect 46452 18358 46508 18396
rect 46620 17668 46676 17678
rect 46620 17574 46676 17612
rect 46732 17444 46788 18956
rect 46620 17388 46788 17444
rect 46284 16994 46396 17006
rect 46284 16942 46342 16994
rect 46394 16942 46396 16994
rect 46284 16940 46396 16942
rect 46340 16930 46396 16940
rect 45948 16830 45950 16882
rect 46002 16830 46004 16882
rect 45948 16818 46004 16830
rect 46060 16826 46116 16838
rect 46060 16774 46062 16826
rect 46114 16774 46116 16826
rect 46060 16660 46116 16774
rect 45836 16604 46116 16660
rect 45724 16212 45780 16222
rect 45724 15341 45780 16156
rect 45724 15289 45726 15341
rect 45778 15289 45780 15341
rect 45724 15277 45780 15289
rect 46396 15316 46452 15326
rect 46396 15222 46452 15260
rect 46060 14532 46116 14542
rect 46396 14532 46452 14542
rect 45948 14530 46116 14532
rect 45183 14474 45239 14486
rect 45183 14422 45185 14474
rect 45237 14422 45239 14474
rect 45183 14420 45239 14422
rect 45183 14354 45239 14364
rect 45948 14478 46062 14530
rect 46114 14478 46116 14530
rect 45948 14476 46116 14478
rect 45948 13746 46004 14476
rect 46060 14466 46116 14476
rect 46284 14530 46452 14532
rect 46284 14478 46398 14530
rect 46450 14478 46452 14530
rect 46284 14476 46452 14478
rect 46172 13748 46228 13758
rect 45948 13694 45950 13746
rect 46002 13694 46004 13746
rect 45612 13636 45668 13646
rect 45948 13636 46004 13694
rect 45276 13634 46004 13636
rect 45276 13582 45614 13634
rect 45666 13582 46004 13634
rect 45276 13580 46004 13582
rect 46060 13746 46228 13748
rect 46060 13694 46174 13746
rect 46226 13694 46228 13746
rect 46060 13692 46228 13694
rect 45276 12962 45332 13580
rect 45612 13570 45668 13580
rect 46060 13076 46116 13692
rect 46172 13682 46228 13692
rect 46284 13524 46340 14476
rect 46396 14466 46452 14476
rect 45668 13020 46116 13076
rect 46172 13468 46340 13524
rect 46452 13524 46508 13534
rect 45668 13018 45724 13020
rect 45276 12910 45278 12962
rect 45330 12910 45332 12962
rect 45276 12898 45332 12910
rect 45500 12964 45556 12974
rect 45668 12966 45670 13018
rect 45722 12966 45724 13018
rect 45668 12954 45724 12966
rect 45500 12870 45556 12908
rect 45836 12290 45892 13020
rect 45836 12238 45838 12290
rect 45890 12238 45892 12290
rect 45836 12226 45892 12238
rect 46172 11732 46228 13468
rect 46452 13430 46508 13468
rect 46620 13076 46676 17388
rect 46956 17108 47012 19740
rect 47180 19234 47236 19246
rect 47180 19182 47182 19234
rect 47234 19182 47236 19234
rect 47068 18676 47124 18686
rect 47180 18676 47236 19182
rect 47292 19236 47348 19966
rect 48076 20634 48132 20646
rect 48076 20582 48078 20634
rect 48130 20582 48132 20634
rect 48076 19572 48132 20582
rect 48300 20356 48356 20694
rect 48300 20290 48356 20300
rect 48524 20750 48638 20802
rect 48690 20750 48692 20802
rect 48524 20748 48692 20750
rect 47292 19170 47348 19180
rect 47404 19516 48132 19572
rect 47068 18674 47236 18676
rect 47068 18622 47070 18674
rect 47122 18622 47236 18674
rect 47068 18620 47236 18622
rect 47068 18610 47124 18620
rect 47404 18450 47460 19516
rect 47404 18398 47406 18450
rect 47458 18398 47460 18450
rect 47404 18386 47460 18398
rect 47516 18452 47572 18462
rect 48524 18452 48580 20748
rect 48636 20738 48692 20748
rect 48636 20020 48692 20030
rect 48636 19348 48692 19964
rect 48748 19684 48804 24332
rect 48972 23044 49028 23054
rect 48972 22950 49028 22988
rect 49308 22708 49364 25454
rect 49420 23380 49476 26852
rect 49420 23314 49476 23324
rect 48972 22652 49364 22708
rect 48972 22370 49028 22652
rect 48972 22318 48974 22370
rect 49026 22318 49028 22370
rect 48860 21700 48916 21710
rect 48860 21586 48916 21644
rect 48860 21534 48862 21586
rect 48914 21534 48916 21586
rect 48860 21522 48916 21534
rect 48860 21364 48916 21374
rect 48860 20018 48916 21308
rect 48972 20804 49028 22318
rect 49140 21362 49196 21374
rect 49140 21310 49142 21362
rect 49194 21310 49196 21362
rect 49140 20804 49196 21310
rect 49140 20748 49364 20804
rect 48972 20738 49028 20748
rect 48860 19966 48862 20018
rect 48914 19966 48916 20018
rect 48860 19954 48916 19966
rect 49308 20468 49364 20748
rect 49140 19794 49196 19806
rect 49140 19742 49142 19794
rect 49194 19742 49196 19794
rect 49140 19684 49196 19742
rect 48748 19628 49196 19684
rect 49308 19572 49364 20412
rect 48636 19282 48692 19292
rect 48972 19516 49364 19572
rect 48804 18452 48860 18462
rect 48524 18450 48860 18452
rect 48524 18398 48806 18450
rect 48858 18398 48860 18450
rect 48524 18396 48860 18398
rect 48972 18452 49028 19516
rect 49532 19460 49588 36988
rect 49644 34132 49700 34142
rect 49644 31892 49700 34076
rect 49644 31826 49700 31836
rect 49532 19394 49588 19404
rect 49084 19348 49140 19358
rect 49140 19292 49252 19348
rect 49084 19254 49140 19292
rect 49084 18452 49140 18462
rect 48972 18450 49140 18452
rect 48972 18398 49086 18450
rect 49138 18398 49140 18450
rect 48972 18396 49140 18398
rect 47516 18358 47572 18396
rect 48804 18386 48860 18396
rect 49084 18386 49140 18396
rect 49196 18450 49252 19292
rect 49196 18398 49198 18450
rect 49250 18398 49252 18450
rect 49196 18386 49252 18398
rect 49308 19236 49364 19246
rect 47852 18228 47908 18238
rect 47852 18226 48580 18228
rect 47852 18174 47854 18226
rect 47906 18174 48580 18226
rect 47852 18172 48580 18174
rect 47852 18162 47908 18172
rect 48524 17778 48580 18172
rect 48524 17726 48526 17778
rect 48578 17726 48580 17778
rect 48524 17714 48580 17726
rect 48972 17892 49028 17902
rect 46956 17052 47236 17108
rect 46900 16911 46956 16923
rect 46900 16859 46902 16911
rect 46954 16899 46956 16911
rect 46954 16859 47012 16899
rect 46900 16843 47012 16859
rect 46732 16772 46788 16782
rect 46732 16770 46900 16772
rect 46732 16718 46734 16770
rect 46786 16718 46900 16770
rect 46732 16716 46900 16718
rect 46732 16706 46788 16716
rect 46844 16210 46900 16716
rect 46844 16158 46846 16210
rect 46898 16158 46900 16210
rect 46844 16146 46900 16158
rect 46956 15988 47012 16843
rect 47068 16884 47124 16894
rect 47068 16790 47124 16828
rect 47180 16436 47236 17052
rect 48972 17106 49028 17836
rect 49308 17666 49364 19180
rect 49308 17614 49310 17666
rect 49362 17614 49364 17666
rect 49308 17602 49364 17614
rect 49420 19124 49476 19134
rect 48972 17054 48974 17106
rect 49026 17054 49028 17106
rect 48972 17042 49028 17054
rect 46844 15932 47012 15988
rect 47068 16380 47236 16436
rect 49308 16884 49364 16894
rect 49420 16884 49476 19068
rect 49308 16882 49476 16884
rect 49308 16830 49310 16882
rect 49362 16830 49476 16882
rect 49308 16828 49476 16830
rect 46732 15314 46788 15326
rect 46732 15262 46734 15314
rect 46786 15262 46788 15314
rect 46732 15204 46788 15262
rect 46732 15138 46788 15148
rect 46844 15146 46900 15932
rect 47068 15876 47124 16380
rect 47516 16268 47796 16324
rect 46844 15094 46846 15146
rect 46898 15094 46900 15146
rect 46844 15082 46900 15094
rect 46956 15820 47124 15876
rect 47180 15876 47236 15886
rect 46620 13020 46900 13076
rect 46620 12850 46676 12862
rect 46620 12798 46622 12850
rect 46674 12798 46676 12850
rect 46620 12193 46676 12798
rect 46284 12178 46340 12190
rect 46284 12126 46286 12178
rect 46338 12126 46340 12178
rect 46284 11844 46340 12126
rect 46284 11778 46340 11788
rect 46620 12141 46622 12193
rect 46674 12141 46676 12193
rect 46172 11666 46228 11676
rect 45500 11396 45556 11406
rect 46620 11396 46676 12141
rect 46732 12068 46788 12078
rect 46732 11974 46788 12012
rect 45500 11394 45780 11396
rect 45500 11342 45502 11394
rect 45554 11342 45780 11394
rect 45500 11340 45780 11342
rect 45500 11330 45556 11340
rect 45500 10052 45556 10062
rect 45500 9940 45556 9996
rect 45388 9938 45556 9940
rect 45388 9886 45502 9938
rect 45554 9886 45556 9938
rect 45388 9884 45556 9886
rect 45052 9772 45220 9828
rect 44996 9604 45052 9614
rect 44996 9510 45052 9548
rect 44546 9018 44660 9044
rect 44492 8988 44660 9018
rect 44380 8876 44548 8932
rect 44324 8372 44380 8382
rect 44156 8370 44380 8372
rect 44156 8318 44326 8370
rect 44378 8318 44380 8370
rect 44156 8316 44380 8318
rect 44324 8306 44380 8316
rect 43260 6850 43316 6860
rect 43708 7308 43876 7364
rect 44380 8036 44436 8046
rect 43708 6804 43764 7308
rect 43932 7252 43988 7262
rect 43148 6610 43150 6662
rect 43202 6610 43204 6662
rect 43596 6748 43764 6804
rect 43820 7250 43988 7252
rect 43820 7198 43934 7250
rect 43986 7198 43988 7250
rect 43820 7196 43988 7198
rect 43148 6598 43204 6610
rect 43372 6634 43428 6646
rect 42868 6580 42924 6590
rect 43372 6582 43374 6634
rect 43426 6582 43428 6634
rect 42868 6578 43092 6580
rect 42868 6526 42870 6578
rect 42922 6526 43092 6578
rect 42868 6524 43092 6526
rect 42868 6514 42924 6524
rect 42588 6178 42644 6188
rect 41916 6076 42084 6132
rect 41692 5796 41748 5806
rect 41692 5794 41860 5796
rect 41692 5742 41694 5794
rect 41746 5742 41860 5794
rect 41692 5740 41860 5742
rect 41692 5730 41748 5740
rect 41580 5618 41636 5628
rect 41468 5292 41748 5348
rect 41692 5094 41748 5292
rect 41692 5042 41694 5094
rect 41746 5042 41748 5094
rect 41692 5030 41748 5042
rect 41356 4286 41358 4338
rect 41410 4286 41412 4338
rect 41356 4274 41412 4286
rect 39340 3554 39508 3556
rect 39340 3502 39342 3554
rect 39394 3502 39508 3554
rect 39340 3500 39508 3502
rect 40908 3948 41020 4004
rect 39116 3490 39172 3500
rect 39340 3490 39396 3500
rect 40572 3444 40628 3482
rect 40572 3378 40628 3388
rect 38780 2492 39060 2548
rect 38780 800 38836 2492
rect 40908 2212 40964 3948
rect 41804 3780 41860 5740
rect 41916 5572 41972 6076
rect 41916 5516 42196 5572
rect 41916 5348 41972 5358
rect 41916 5012 41972 5292
rect 41916 4956 42084 5012
rect 41804 3714 41860 3724
rect 42028 4452 42084 4956
rect 42028 3526 42084 4396
rect 42140 4338 42196 5516
rect 43036 5124 43092 6524
rect 43372 6132 43428 6582
rect 43596 6634 43652 6748
rect 43596 6582 43598 6634
rect 43650 6582 43652 6634
rect 43596 6244 43652 6582
rect 43372 6066 43428 6076
rect 43484 6188 43652 6244
rect 43708 6634 43764 6646
rect 43708 6582 43710 6634
rect 43762 6582 43764 6634
rect 43484 5908 43540 6188
rect 43596 6020 43652 6030
rect 43708 6020 43764 6582
rect 43596 6018 43708 6020
rect 43596 5966 43598 6018
rect 43650 5966 43708 6018
rect 43596 5964 43708 5966
rect 43596 5954 43652 5964
rect 43708 5926 43764 5964
rect 43484 5236 43540 5852
rect 43484 5170 43540 5180
rect 43036 5068 43316 5124
rect 43036 4900 43092 4910
rect 43036 4806 43092 4844
rect 42140 4286 42142 4338
rect 42194 4286 42196 4338
rect 42140 4274 42196 4286
rect 42364 4788 42420 4798
rect 42028 3474 42030 3526
rect 42082 3474 42084 3526
rect 42028 3462 42084 3474
rect 40572 2156 40964 2212
rect 40572 800 40628 2156
rect 42364 800 42420 4732
rect 42700 3780 42756 3790
rect 42700 3686 42756 3724
rect 43036 3556 43092 3566
rect 43260 3556 43316 5068
rect 43820 4116 43876 7196
rect 43932 7186 43988 7196
rect 44212 6468 44268 6478
rect 43820 4050 43876 4060
rect 43932 6466 44268 6468
rect 43932 6414 44214 6466
rect 44266 6414 44268 6466
rect 43932 6412 44268 6414
rect 43932 4004 43988 6412
rect 44212 6402 44268 6412
rect 44100 6244 44156 6254
rect 44380 6244 44436 7980
rect 44492 7476 44548 8876
rect 44604 8148 44660 8988
rect 44716 9018 44718 9070
rect 44770 9018 44772 9070
rect 44716 8820 44772 9018
rect 44716 8754 44772 8764
rect 44828 9077 44884 9089
rect 44828 9025 44830 9077
rect 44882 9025 44884 9077
rect 44828 8372 44884 9025
rect 45164 8372 45220 9772
rect 44828 8306 44884 8316
rect 45052 8316 45220 8372
rect 44604 8082 44660 8092
rect 45052 8036 45108 8316
rect 45276 8260 45332 8270
rect 45164 8202 45220 8214
rect 45164 8150 45166 8202
rect 45218 8150 45220 8202
rect 45276 8178 45278 8204
rect 45330 8178 45332 8204
rect 45276 8166 45332 8178
rect 45164 8036 45220 8150
rect 45388 8036 45444 9884
rect 45500 9874 45556 9884
rect 45612 9828 45668 9838
rect 45612 9069 45668 9772
rect 45612 9017 45614 9069
rect 45666 9017 45668 9069
rect 45612 9005 45668 9017
rect 45724 8372 45780 11340
rect 46620 11330 46676 11340
rect 46844 10724 46900 13020
rect 46844 10658 46900 10668
rect 46060 10388 46116 10398
rect 46060 9828 46116 10332
rect 46060 9762 46116 9772
rect 46172 10164 46228 10174
rect 46956 10164 47012 15820
rect 47180 14642 47236 15820
rect 47348 15316 47404 15326
rect 47348 15222 47404 15260
rect 47516 15148 47572 16268
rect 47628 16098 47684 16110
rect 47628 16046 47630 16098
rect 47682 16046 47684 16098
rect 47628 15540 47684 16046
rect 47740 16098 47796 16268
rect 49308 16222 49364 16828
rect 49252 16210 49364 16222
rect 49252 16158 49254 16210
rect 49306 16158 49364 16210
rect 49252 16156 49364 16158
rect 49252 16146 49308 16156
rect 47740 16046 47742 16098
rect 47794 16046 47796 16098
rect 47740 16034 47796 16046
rect 48076 15876 48132 15886
rect 48076 15782 48132 15820
rect 47628 15474 47684 15484
rect 47740 15329 47796 15341
rect 47740 15277 47742 15329
rect 47794 15277 47796 15329
rect 47404 15092 47572 15148
rect 47628 15202 47684 15214
rect 47628 15150 47630 15202
rect 47682 15150 47684 15202
rect 47180 14590 47182 14642
rect 47234 14590 47236 14642
rect 47180 14578 47236 14590
rect 47292 14868 47348 14878
rect 47180 13746 47236 13758
rect 47180 13694 47182 13746
rect 47234 13694 47236 13746
rect 47180 12852 47236 13694
rect 47292 13748 47348 14812
rect 47404 13914 47460 15092
rect 47628 14868 47684 15150
rect 47740 14980 47796 15277
rect 47740 14914 47796 14924
rect 48076 15314 48132 15326
rect 48076 15262 48078 15314
rect 48130 15262 48132 15314
rect 47628 14802 47684 14812
rect 48076 14868 48132 15262
rect 48636 15314 48692 15326
rect 48636 15262 48638 15314
rect 48690 15262 48692 15314
rect 48636 15148 48692 15262
rect 48076 14802 48132 14812
rect 48300 15092 48692 15148
rect 48300 13972 48356 15092
rect 48972 15090 49028 15102
rect 48972 15038 48974 15090
rect 49026 15038 49028 15090
rect 48860 14980 48916 14990
rect 47404 13862 47406 13914
rect 47458 13862 47460 13914
rect 47404 13850 47460 13862
rect 47964 13916 48356 13972
rect 48636 14868 48692 14878
rect 47516 13773 47572 13785
rect 47516 13748 47518 13773
rect 47292 13721 47518 13748
rect 47570 13721 47572 13773
rect 47292 13692 47572 13721
rect 47852 13748 47908 13758
rect 47852 13654 47908 13692
rect 47964 13300 48020 13916
rect 47180 12178 47236 12796
rect 47180 12126 47182 12178
rect 47234 12126 47236 12178
rect 47180 12114 47236 12126
rect 47292 13244 48020 13300
rect 48300 13748 48356 13758
rect 46956 10108 47236 10164
rect 45612 8316 45780 8372
rect 45500 8202 45556 8214
rect 45500 8150 45502 8202
rect 45554 8150 45556 8202
rect 45500 8148 45556 8150
rect 45500 8082 45556 8092
rect 45164 7980 45444 8036
rect 45052 7970 45108 7980
rect 45500 7812 45556 7822
rect 45276 7588 45332 7598
rect 45500 7588 45556 7756
rect 45276 7530 45332 7532
rect 44772 7509 44828 7521
rect 44772 7476 44774 7509
rect 44492 7410 44548 7420
rect 44716 7457 44774 7476
rect 44826 7457 44828 7509
rect 44716 7420 44828 7457
rect 45052 7502 45108 7514
rect 45052 7450 45054 7502
rect 45106 7450 45108 7502
rect 44548 7252 44604 7262
rect 44548 7158 44604 7196
rect 44604 6580 44660 6590
rect 44716 6580 44772 7420
rect 45052 6804 45108 7450
rect 45276 7478 45278 7530
rect 45330 7478 45332 7530
rect 45276 6916 45332 7478
rect 45463 7532 45556 7588
rect 45463 7530 45519 7532
rect 45463 7478 45465 7530
rect 45517 7478 45519 7530
rect 45463 7466 45519 7478
rect 45276 6860 45556 6916
rect 45500 6804 45556 6860
rect 45052 6748 45444 6804
rect 45108 6634 45164 6646
rect 44660 6524 44772 6580
rect 44884 6578 44940 6590
rect 45108 6582 45110 6634
rect 45162 6582 45164 6634
rect 45108 6580 45164 6582
rect 44884 6526 44886 6578
rect 44938 6526 44940 6578
rect 44604 6514 44660 6524
rect 44100 6018 44156 6188
rect 44100 5966 44102 6018
rect 44154 5966 44156 6018
rect 44100 5954 44156 5966
rect 44268 6188 44436 6244
rect 43932 3938 43988 3948
rect 44044 5460 44100 5470
rect 44044 4450 44100 5404
rect 44044 4398 44046 4450
rect 44098 4398 44100 4450
rect 43036 3554 43316 3556
rect 43036 3502 43038 3554
rect 43090 3502 43316 3554
rect 43036 3500 43316 3502
rect 43764 3556 43820 3566
rect 43036 3490 43092 3500
rect 43764 3462 43820 3500
rect 44044 3526 44100 4398
rect 44044 3474 44046 3526
rect 44098 3474 44100 3526
rect 44044 3462 44100 3474
rect 44156 4900 44212 4910
rect 44156 800 44212 4844
rect 44268 3668 44324 6188
rect 44884 6132 44940 6526
rect 44716 6076 44940 6132
rect 45052 6524 45164 6580
rect 45388 6634 45444 6748
rect 45612 6804 45668 8316
rect 45747 8202 45803 8214
rect 45747 8150 45749 8202
rect 45801 8150 45803 8202
rect 45747 8036 45803 8150
rect 46004 8148 46060 8158
rect 46172 8148 46228 10108
rect 47180 9604 47236 10108
rect 46956 9548 47236 9604
rect 46004 8146 46228 8148
rect 46004 8094 46006 8146
rect 46058 8094 46228 8146
rect 46004 8092 46228 8094
rect 46284 8148 46340 8158
rect 46004 8082 46060 8092
rect 45724 7980 45803 8036
rect 45724 7812 45780 7980
rect 45724 7746 45780 7756
rect 45724 7501 45780 7513
rect 45724 7449 45726 7501
rect 45778 7449 45780 7501
rect 45724 7364 45780 7449
rect 45724 7298 45780 7308
rect 45612 6748 45892 6804
rect 45500 6692 45556 6748
rect 45500 6655 45612 6692
rect 45500 6636 45558 6655
rect 45388 6582 45390 6634
rect 45442 6582 45444 6634
rect 45556 6603 45558 6636
rect 45610 6603 45612 6655
rect 45556 6591 45612 6603
rect 45724 6634 45780 6646
rect 44380 6020 44436 6030
rect 44380 5962 44436 5964
rect 44380 5910 44382 5962
rect 44434 5910 44436 5962
rect 44604 6020 44660 6030
rect 44604 5962 44660 5964
rect 44380 5898 44436 5910
rect 44492 5908 44548 5918
rect 44604 5910 44606 5962
rect 44658 5910 44660 5962
rect 44604 5898 44660 5910
rect 44268 3612 44436 3668
rect 44268 3498 44324 3510
rect 44268 3446 44270 3498
rect 44322 3446 44324 3498
rect 44268 3444 44324 3446
rect 44268 3378 44324 3388
rect 44380 3388 44436 3612
rect 44492 3526 44548 5852
rect 44716 5012 44772 6076
rect 44828 5934 44884 5946
rect 44828 5908 44830 5934
rect 44882 5908 44884 5934
rect 44828 5842 44884 5852
rect 44940 5941 44996 5953
rect 44940 5889 44942 5941
rect 44994 5889 44996 5941
rect 44940 5460 44996 5889
rect 44940 5394 44996 5404
rect 44940 5236 44996 5246
rect 44940 5142 44996 5180
rect 44716 4946 44772 4956
rect 45052 4788 45108 6524
rect 45388 6244 45444 6582
rect 45724 6582 45726 6634
rect 45778 6582 45780 6634
rect 45388 6178 45444 6188
rect 45500 6468 45556 6478
rect 44492 3474 44494 3526
rect 44546 3474 44548 3526
rect 44492 3462 44548 3474
rect 44604 4732 45108 4788
rect 45164 6020 45220 6030
rect 44604 4450 44660 4732
rect 44604 4398 44606 4450
rect 44658 4398 44660 4450
rect 44604 3519 44660 4398
rect 44604 3467 44606 3519
rect 44658 3467 44660 3519
rect 44604 3455 44660 3467
rect 45164 3444 45220 5964
rect 45388 5236 45444 5246
rect 45388 3668 45444 5180
rect 45500 4788 45556 6412
rect 45612 5794 45668 5806
rect 45612 5742 45614 5794
rect 45666 5742 45668 5794
rect 45612 5348 45668 5742
rect 45612 4788 45668 5292
rect 45724 5236 45780 6582
rect 45836 6020 45892 6748
rect 46116 6468 46172 6478
rect 46116 6374 46172 6412
rect 45836 5954 45892 5964
rect 46284 5572 46340 8092
rect 46620 8146 46676 8158
rect 46620 8094 46622 8146
rect 46674 8094 46676 8146
rect 46620 7812 46676 8094
rect 46620 7746 46676 7756
rect 46284 5506 46340 5516
rect 46396 6804 46452 6814
rect 46396 5460 46452 6748
rect 46620 6580 46676 6590
rect 46620 6486 46676 6524
rect 46956 6356 47012 9548
rect 47292 7476 47348 13244
rect 48300 12740 48356 13692
rect 48636 13746 48692 14812
rect 48636 13694 48638 13746
rect 48690 13694 48692 13746
rect 48636 13682 48692 13694
rect 48860 13748 48916 14924
rect 48860 13654 48916 13692
rect 48972 13076 49028 15038
rect 49084 14868 49140 14878
rect 49084 14642 49140 14812
rect 49084 14590 49086 14642
rect 49138 14590 49140 14642
rect 49084 14578 49140 14590
rect 49140 13636 49196 13646
rect 49140 13542 49196 13580
rect 48972 13020 49140 13076
rect 48524 12964 48580 12974
rect 48524 12962 49028 12964
rect 48524 12910 48526 12962
rect 48578 12910 49028 12962
rect 48524 12908 49028 12910
rect 48524 12898 48580 12908
rect 47740 12684 48356 12740
rect 47404 12205 47460 12217
rect 47404 12153 47406 12205
rect 47458 12153 47460 12205
rect 47404 12068 47460 12153
rect 47404 12002 47460 12012
rect 47740 12178 47796 12684
rect 48972 12402 49028 12908
rect 47740 12126 47742 12178
rect 47794 12126 47796 12178
rect 47740 11956 47796 12126
rect 47852 12346 47908 12358
rect 47852 12294 47854 12346
rect 47906 12294 47908 12346
rect 48972 12350 48974 12402
rect 49026 12350 49028 12402
rect 48972 12338 49028 12350
rect 47852 12180 47908 12294
rect 48636 12180 48692 12190
rect 47852 12178 48692 12180
rect 47852 12126 48638 12178
rect 48690 12126 48692 12178
rect 47852 12124 48692 12126
rect 48636 12114 48692 12124
rect 47740 11900 48300 11956
rect 48244 11618 48300 11900
rect 48244 11566 48246 11618
rect 48298 11566 48300 11618
rect 48244 11554 48300 11566
rect 48412 11844 48468 11854
rect 47852 11394 47908 11406
rect 47852 11342 47854 11394
rect 47906 11342 47908 11394
rect 47404 11284 47460 11294
rect 47852 11284 47908 11342
rect 47964 11396 48020 11406
rect 47964 11302 48020 11340
rect 47404 11282 47908 11284
rect 47404 11230 47406 11282
rect 47458 11230 47908 11282
rect 47404 11228 47908 11230
rect 47404 11218 47460 11228
rect 47404 10637 47460 10650
rect 47404 10612 47406 10637
rect 47458 10612 47460 10637
rect 47404 10546 47460 10556
rect 47404 10388 47460 10398
rect 47852 10388 47908 11228
rect 48244 10612 48300 10622
rect 48244 10518 48300 10556
rect 47852 10332 48356 10388
rect 47404 9938 47460 10332
rect 47404 9886 47406 9938
rect 47458 9886 47460 9938
rect 47404 9874 47460 9886
rect 48188 9828 48244 9838
rect 48188 9734 48244 9772
rect 48300 9826 48356 10332
rect 48412 9940 48468 11788
rect 48524 11394 48580 11406
rect 48524 11342 48526 11394
rect 48578 11342 48580 11394
rect 48524 10500 48580 11342
rect 48860 11170 48916 11182
rect 48860 11118 48862 11170
rect 48914 11118 48916 11170
rect 48524 10434 48580 10444
rect 48636 10610 48692 10622
rect 48636 10558 48638 10610
rect 48690 10558 48692 10610
rect 48636 10164 48692 10558
rect 48636 10098 48692 10108
rect 48636 9940 48692 9950
rect 48412 9938 48692 9940
rect 48412 9886 48638 9938
rect 48690 9886 48692 9938
rect 48412 9884 48692 9886
rect 48636 9874 48692 9884
rect 48300 9774 48302 9826
rect 48354 9774 48356 9826
rect 48300 9762 48356 9774
rect 48132 9210 48188 9222
rect 48132 9158 48134 9210
rect 48186 9158 48188 9210
rect 48132 8596 48188 9158
rect 48636 9044 48692 9054
rect 48636 9042 48804 9044
rect 48636 8990 48638 9042
rect 48690 8990 48804 9042
rect 48636 8988 48804 8990
rect 48636 8978 48692 8988
rect 47180 7420 47348 7476
rect 47404 8540 48188 8596
rect 48636 8820 48692 8830
rect 47068 7250 47124 7262
rect 47068 7198 47070 7250
rect 47122 7198 47124 7250
rect 47068 6692 47124 7198
rect 47068 6626 47124 6636
rect 46956 6290 47012 6300
rect 47180 6132 47236 7420
rect 47180 6066 47236 6076
rect 47292 7252 47348 7262
rect 46956 5572 47012 5582
rect 46396 5404 46676 5460
rect 45724 5170 45780 5180
rect 46620 5236 46676 5404
rect 45612 4732 46340 4788
rect 45500 4722 45556 4732
rect 45948 4004 46004 4014
rect 45836 3892 45892 3902
rect 45388 3612 45556 3668
rect 45500 3556 45556 3612
rect 45500 3519 45612 3556
rect 45500 3500 45558 3519
rect 44380 3332 44772 3388
rect 45164 3378 45220 3388
rect 45332 3444 45388 3482
rect 45556 3467 45558 3500
rect 45610 3467 45612 3519
rect 45556 3455 45612 3467
rect 45836 3526 45892 3836
rect 45836 3474 45838 3526
rect 45890 3474 45892 3526
rect 45836 3462 45892 3474
rect 45332 3378 45388 3388
rect 44716 2100 44772 3332
rect 44716 2034 44772 2044
rect 45948 800 46004 3948
rect 46284 3556 46340 4732
rect 46508 4226 46564 4238
rect 46508 4174 46510 4226
rect 46562 4174 46564 4226
rect 46508 3780 46564 4174
rect 46508 3714 46564 3724
rect 46620 3556 46676 5180
rect 46844 5122 46900 5134
rect 46844 5070 46846 5122
rect 46898 5070 46900 5122
rect 46228 3538 46340 3556
rect 46060 3498 46116 3510
rect 46060 3446 46062 3498
rect 46114 3446 46116 3498
rect 46228 3486 46230 3538
rect 46282 3500 46340 3538
rect 46396 3500 46676 3556
rect 46732 4788 46788 4798
rect 46282 3486 46284 3500
rect 46228 3474 46284 3486
rect 46060 3388 46116 3446
rect 46396 3388 46452 3500
rect 46060 3332 46452 3388
rect 46732 3444 46788 4732
rect 46844 4228 46900 5070
rect 46844 4162 46900 4172
rect 46956 3554 47012 5516
rect 47292 5460 47348 7196
rect 47404 5572 47460 8540
rect 48524 8260 48580 8270
rect 48412 8258 48580 8260
rect 48412 8206 48526 8258
rect 48578 8206 48580 8258
rect 48412 8204 48580 8206
rect 48300 6692 48356 6702
rect 47852 6468 47908 6478
rect 47740 6132 47796 6142
rect 47516 5908 47572 5918
rect 47516 5814 47572 5852
rect 47404 5516 47572 5572
rect 47292 5404 47460 5460
rect 47068 5124 47124 5134
rect 47292 5124 47348 5134
rect 47124 5068 47236 5124
rect 47068 5058 47124 5068
rect 46956 3502 46958 3554
rect 47010 3502 47012 3554
rect 46956 3490 47012 3502
rect 47180 3556 47236 5068
rect 47292 4338 47348 5068
rect 47292 4286 47294 4338
rect 47346 4286 47348 4338
rect 47292 4274 47348 4286
rect 47404 4338 47460 5404
rect 47404 4286 47406 4338
rect 47458 4286 47460 4338
rect 47404 4274 47460 4286
rect 47516 3892 47572 5516
rect 47628 5124 47684 5134
rect 47628 5030 47684 5068
rect 47740 4562 47796 6076
rect 47852 5087 47908 6412
rect 48300 5908 48356 6636
rect 48412 6132 48468 8204
rect 48524 8194 48580 8204
rect 48636 7474 48692 8764
rect 48748 8260 48804 8988
rect 48748 7700 48804 8204
rect 48860 7924 48916 11118
rect 48972 10388 49028 10398
rect 48972 10294 49028 10332
rect 49084 10164 49140 13020
rect 48972 10108 49140 10164
rect 49308 12962 49364 12974
rect 49308 12910 49310 12962
rect 49362 12910 49364 12962
rect 48972 9380 49028 10108
rect 49308 9828 49364 12910
rect 49308 9762 49364 9772
rect 49140 9604 49196 9614
rect 49140 9602 49588 9604
rect 49140 9550 49142 9602
rect 49194 9550 49588 9602
rect 49140 9548 49588 9550
rect 49140 9538 49196 9548
rect 48972 9324 49140 9380
rect 48972 8818 49028 8830
rect 48972 8766 48974 8818
rect 49026 8766 49028 8818
rect 48972 8484 49028 8766
rect 48972 8418 49028 8428
rect 48860 7858 48916 7868
rect 48972 7700 49028 7710
rect 48748 7698 49028 7700
rect 48748 7646 48974 7698
rect 49026 7646 49028 7698
rect 48748 7644 49028 7646
rect 48972 7634 49028 7644
rect 48636 7422 48638 7474
rect 48690 7422 48692 7474
rect 48636 7410 48692 7422
rect 48524 6692 48580 6702
rect 48524 6690 49028 6692
rect 48524 6638 48526 6690
rect 48578 6638 49028 6690
rect 48524 6636 49028 6638
rect 48524 6626 48580 6636
rect 48412 6066 48468 6076
rect 48636 5908 48692 5918
rect 48300 5906 48692 5908
rect 48300 5854 48302 5906
rect 48354 5854 48638 5906
rect 48690 5854 48692 5906
rect 48300 5852 48692 5854
rect 47852 5035 47854 5087
rect 47906 5035 47908 5087
rect 47852 5023 47908 5035
rect 47964 5236 48020 5246
rect 47964 5094 48020 5180
rect 47964 5042 47966 5094
rect 48018 5042 48020 5094
rect 47964 5030 48020 5042
rect 48188 5236 48244 5246
rect 48188 5094 48244 5180
rect 48188 5042 48190 5094
rect 48242 5042 48244 5094
rect 48300 5124 48356 5852
rect 48636 5842 48692 5852
rect 48300 5058 48356 5068
rect 48412 5348 48468 5358
rect 48412 5094 48468 5292
rect 48188 5030 48244 5042
rect 48412 5042 48414 5094
rect 48466 5042 48468 5094
rect 48412 5030 48468 5042
rect 47740 4510 47742 4562
rect 47794 4510 47796 4562
rect 47740 4498 47796 4510
rect 48524 5012 48580 5022
rect 48692 5012 48748 5022
rect 47516 3836 47796 3892
rect 47628 3668 47684 3678
rect 47628 3574 47684 3612
rect 47292 3556 47348 3566
rect 47180 3554 47348 3556
rect 47180 3502 47294 3554
rect 47346 3502 47348 3554
rect 47180 3500 47348 3502
rect 47292 3490 47348 3500
rect 46732 3378 46788 3388
rect 46620 3332 46676 3342
rect 46620 3238 46676 3276
rect 47740 800 47796 3836
rect 48300 3780 48356 3790
rect 48300 3686 48356 3724
rect 47964 3556 48020 3566
rect 48524 3556 48580 4956
rect 48636 5010 48748 5012
rect 48636 4958 48694 5010
rect 48746 4958 48748 5010
rect 48636 4946 48748 4958
rect 48636 4338 48692 4946
rect 48972 4562 49028 6636
rect 49084 5908 49140 9324
rect 49308 8258 49364 8270
rect 49308 8206 49310 8258
rect 49362 8206 49364 8258
rect 49084 5842 49140 5852
rect 49196 7924 49252 7934
rect 49196 6244 49252 7868
rect 49308 6692 49364 8206
rect 49308 6598 49364 6636
rect 49196 5236 49252 6188
rect 49196 5170 49252 5180
rect 49140 4900 49196 4910
rect 49140 4806 49196 4844
rect 48972 4510 48974 4562
rect 49026 4510 49028 4562
rect 48972 4498 49028 4510
rect 48636 4286 48638 4338
rect 48690 4286 48692 4338
rect 48636 4274 48692 4286
rect 48972 4228 49028 4238
rect 48972 3778 49028 4172
rect 48972 3726 48974 3778
rect 49026 3726 49028 3778
rect 48972 3714 49028 3726
rect 48636 3556 48692 3566
rect 48524 3554 48692 3556
rect 48524 3502 48638 3554
rect 48690 3502 48692 3554
rect 48524 3500 48692 3502
rect 47964 3462 48020 3500
rect 48636 3490 48692 3500
rect 49532 800 49588 9548
rect 1120 0 1232 800
rect 2912 0 3024 800
rect 4704 0 4816 800
rect 6496 0 6608 800
rect 8288 0 8400 800
rect 10080 0 10192 800
rect 11872 0 11984 800
rect 13664 0 13776 800
rect 15456 0 15568 800
rect 17248 0 17360 800
rect 19040 0 19152 800
rect 20832 0 20944 800
rect 22624 0 22736 800
rect 24416 0 24528 800
rect 26208 0 26320 800
rect 28000 0 28112 800
rect 29792 0 29904 800
rect 31584 0 31696 800
rect 33376 0 33488 800
rect 35168 0 35280 800
rect 36960 0 37072 800
rect 38752 0 38864 800
rect 40544 0 40656 800
rect 42336 0 42448 800
rect 44128 0 44240 800
rect 45920 0 46032 800
rect 47712 0 47824 800
rect 49504 0 49616 800
<< via2 >>
rect 5740 48300 5796 48356
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 5628 41244 5684 41300
rect 5404 40460 5460 40516
rect 6300 48300 6356 48356
rect 11116 45948 11172 46004
rect 11452 45836 11508 45892
rect 12012 45890 12068 45892
rect 12012 45838 12014 45890
rect 12014 45838 12066 45890
rect 12066 45838 12068 45890
rect 12012 45836 12068 45838
rect 11340 45724 11396 45780
rect 11676 45724 11732 45780
rect 9100 44546 9156 44548
rect 9100 44494 9102 44546
rect 9102 44494 9154 44546
rect 9154 44494 9156 44546
rect 9100 44492 9156 44494
rect 7868 44044 7924 44100
rect 8764 44268 8820 44324
rect 7532 43708 7588 43764
rect 7196 43260 7252 43316
rect 7439 43036 7495 43092
rect 6412 41970 6468 41972
rect 6412 41918 6414 41970
rect 6414 41918 6466 41970
rect 6466 41918 6468 41970
rect 6412 41916 6468 41918
rect 6916 41970 6972 41972
rect 6916 41918 6918 41970
rect 6918 41918 6970 41970
rect 6970 41918 6972 41970
rect 6916 41916 6972 41918
rect 6636 41804 6692 41860
rect 7756 41933 7758 41972
rect 7758 41933 7810 41972
rect 7810 41933 7812 41972
rect 7756 41916 7812 41933
rect 10220 44492 10276 44548
rect 9548 44268 9604 44324
rect 9884 44322 9940 44324
rect 9884 44270 9886 44322
rect 9886 44270 9938 44322
rect 9938 44270 9940 44322
rect 9884 44268 9940 44270
rect 9436 44156 9492 44212
rect 11340 44156 11396 44212
rect 11116 44044 11172 44100
rect 8876 43260 8932 43316
rect 9548 42140 9604 42196
rect 7420 41692 7476 41748
rect 6300 41298 6356 41300
rect 6300 41246 6302 41298
rect 6302 41246 6354 41298
rect 6354 41246 6356 41298
rect 6300 41244 6356 41246
rect 5964 40460 6020 40516
rect 6188 40460 6244 40516
rect 5852 40236 5908 40292
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 5964 39618 6020 39620
rect 5740 38892 5796 38948
rect 5964 39566 5966 39618
rect 5966 39566 6018 39618
rect 6018 39566 6020 39618
rect 5964 39564 6020 39566
rect 5516 38780 5572 38836
rect 3500 38722 3556 38724
rect 3500 38670 3502 38722
rect 3502 38670 3554 38722
rect 3554 38670 3556 38722
rect 3500 38668 3556 38670
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 6748 40572 6804 40628
rect 6636 40377 6638 40404
rect 6638 40377 6690 40404
rect 6690 40377 6692 40404
rect 6636 40348 6692 40377
rect 6412 39676 6468 39732
rect 6524 40236 6580 40292
rect 6188 38834 6244 38836
rect 6188 38782 6190 38834
rect 6190 38782 6242 38834
rect 6242 38782 6244 38834
rect 6188 38780 6244 38782
rect 6300 39452 6356 39508
rect 8204 41804 8260 41860
rect 8316 41916 8372 41972
rect 8316 41692 8372 41748
rect 8596 41746 8652 41748
rect 8596 41694 8598 41746
rect 8598 41694 8650 41746
rect 8650 41694 8652 41746
rect 8596 41692 8652 41694
rect 8204 41074 8260 41076
rect 8204 41022 8206 41074
rect 8206 41022 8258 41074
rect 8258 41022 8260 41074
rect 8204 41020 8260 41022
rect 7644 40572 7700 40628
rect 8316 40460 8372 40516
rect 8204 40348 8260 40404
rect 7308 39788 7364 39844
rect 6860 39676 6916 39732
rect 7756 39676 7812 39732
rect 6524 38946 6580 38948
rect 6524 38894 6526 38946
rect 6526 38894 6578 38946
rect 6578 38894 6580 38946
rect 6524 38892 6580 38894
rect 7644 38834 7700 38836
rect 7644 38782 7646 38834
rect 7646 38782 7698 38834
rect 7698 38782 7700 38834
rect 7644 38780 7700 38782
rect 8652 41020 8708 41076
rect 9996 43260 10052 43316
rect 9996 42194 10052 42196
rect 9996 42142 9998 42194
rect 9998 42142 10050 42194
rect 10050 42142 10052 42194
rect 9996 42140 10052 42142
rect 10332 42140 10388 42196
rect 9044 41074 9100 41076
rect 9044 41022 9046 41074
rect 9046 41022 9098 41074
rect 9098 41022 9100 41074
rect 9044 41020 9100 41022
rect 8876 40572 8932 40628
rect 9660 41916 9716 41972
rect 10892 43484 10948 43540
rect 10780 42476 10836 42532
rect 11452 43708 11508 43764
rect 12348 46396 12404 46452
rect 13356 45948 13412 46004
rect 13580 46508 13636 46564
rect 13748 46450 13804 46452
rect 13748 46398 13750 46450
rect 13750 46398 13802 46450
rect 13802 46398 13804 46450
rect 13748 46396 13804 46398
rect 13692 45948 13748 46004
rect 13468 45724 13524 45780
rect 12124 44156 12180 44212
rect 12012 43708 12068 43764
rect 11564 43372 11620 43428
rect 11228 42364 11284 42420
rect 11228 42140 11284 42196
rect 10724 41804 10780 41860
rect 10332 41692 10388 41748
rect 10108 41356 10164 41412
rect 9884 41186 9940 41188
rect 9884 41134 9886 41186
rect 9886 41134 9938 41186
rect 9938 41134 9940 41186
rect 9884 41132 9940 41134
rect 10220 40684 10276 40740
rect 8820 39676 8876 39732
rect 8316 39506 8372 39508
rect 8316 39454 8318 39506
rect 8318 39454 8370 39506
rect 8370 39454 8372 39506
rect 8316 39452 8372 39454
rect 8204 38162 8260 38164
rect 8204 38110 8206 38162
rect 8206 38110 8258 38162
rect 8258 38110 8260 38162
rect 8204 38108 8260 38110
rect 7868 36876 7924 36932
rect 6636 36482 6692 36484
rect 6636 36430 6638 36482
rect 6638 36430 6690 36482
rect 6690 36430 6692 36482
rect 6636 36428 6692 36430
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4844 34914 4900 34916
rect 4844 34862 4846 34914
rect 4846 34862 4898 34914
rect 4898 34862 4900 34914
rect 4844 34860 4900 34862
rect 5180 34860 5236 34916
rect 5516 34860 5572 34916
rect 8092 35868 8148 35924
rect 7868 35810 7924 35812
rect 7868 35758 7870 35810
rect 7870 35758 7922 35810
rect 7922 35758 7924 35810
rect 7868 35756 7924 35758
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 5852 34076 5908 34132
rect 5516 33628 5572 33684
rect 2044 31724 2100 31780
rect 1596 28588 1652 28644
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 6636 34636 6692 34692
rect 7420 34860 7476 34916
rect 6188 34412 6244 34468
rect 6300 34130 6356 34132
rect 6300 34078 6302 34130
rect 6302 34078 6354 34130
rect 6354 34078 6356 34130
rect 6300 34076 6356 34078
rect 6972 33628 7028 33684
rect 9660 40572 9716 40628
rect 9884 40572 9940 40628
rect 9212 39676 9268 39732
rect 9772 40348 9828 40404
rect 10612 41410 10668 41412
rect 10612 41358 10614 41410
rect 10614 41358 10666 41410
rect 10666 41358 10668 41410
rect 10612 41356 10668 41358
rect 10332 40572 10388 40628
rect 10220 40460 10276 40516
rect 10108 40290 10164 40292
rect 10108 40238 10110 40290
rect 10110 40238 10162 40290
rect 10162 40238 10164 40290
rect 10108 40236 10164 40238
rect 10892 41186 10948 41188
rect 10892 41134 10894 41186
rect 10894 41134 10946 41186
rect 10946 41134 10948 41186
rect 10892 41132 10948 41134
rect 11116 41132 11172 41188
rect 9548 39228 9604 39284
rect 8988 38892 9044 38948
rect 8596 38834 8652 38836
rect 8596 38782 8598 38834
rect 8598 38782 8650 38834
rect 8650 38782 8652 38834
rect 8596 38780 8652 38782
rect 8428 38556 8484 38612
rect 8876 38220 8932 38276
rect 8428 38108 8484 38164
rect 9660 38892 9716 38948
rect 10052 38892 10108 38948
rect 9492 38556 9548 38612
rect 9772 38668 9828 38724
rect 9324 38444 9380 38500
rect 11116 40684 11172 40740
rect 10668 40402 10724 40404
rect 10668 40350 10670 40402
rect 10670 40350 10722 40402
rect 10722 40350 10724 40402
rect 10668 40348 10724 40350
rect 10780 40236 10836 40292
rect 10892 39900 10948 39956
rect 11340 41132 11396 41188
rect 11452 42364 11508 42420
rect 13580 45164 13636 45220
rect 14700 45388 14756 45444
rect 16716 46562 16772 46564
rect 16716 46510 16718 46562
rect 16718 46510 16770 46562
rect 16770 46510 16772 46562
rect 16716 46508 16772 46510
rect 17444 46450 17500 46452
rect 17444 46398 17446 46450
rect 17446 46398 17498 46450
rect 17498 46398 17500 46450
rect 17444 46396 17500 46398
rect 12684 44156 12740 44212
rect 13020 43596 13076 43652
rect 12572 43484 12628 43540
rect 11676 42588 11732 42644
rect 12572 42924 12628 42980
rect 12236 42754 12292 42756
rect 12236 42702 12238 42754
rect 12238 42702 12290 42754
rect 12290 42702 12292 42754
rect 12236 42700 12292 42702
rect 12124 42588 12180 42644
rect 12908 42924 12964 42980
rect 12796 42700 12852 42756
rect 13020 42700 13076 42756
rect 12344 41956 12346 41972
rect 12346 41956 12398 41972
rect 12398 41956 12400 41972
rect 12344 41916 12400 41956
rect 13524 43596 13580 43652
rect 13692 43708 13748 43764
rect 13244 43484 13300 43540
rect 13804 43372 13860 43428
rect 14812 44380 14868 44436
rect 14364 43708 14420 43764
rect 14028 43538 14084 43540
rect 14028 43486 14030 43538
rect 14030 43486 14082 43538
rect 14082 43486 14084 43538
rect 14028 43484 14084 43486
rect 13412 43036 13468 43092
rect 12572 41804 12628 41860
rect 11676 41186 11732 41188
rect 11676 41134 11678 41186
rect 11678 41134 11730 41186
rect 11730 41134 11732 41186
rect 11676 41132 11732 41134
rect 11452 40572 11508 40628
rect 10444 39228 10500 39284
rect 11228 39564 11284 39620
rect 10444 39004 10500 39060
rect 11004 38834 11060 38836
rect 11004 38782 11006 38834
rect 11006 38782 11058 38834
rect 11058 38782 11060 38834
rect 11004 38780 11060 38782
rect 11228 39116 11284 39172
rect 11452 40290 11508 40292
rect 11452 40238 11454 40290
rect 11454 40238 11506 40290
rect 11506 40238 11508 40290
rect 11452 40236 11508 40238
rect 12552 41132 12608 41188
rect 11676 39788 11732 39844
rect 11452 39730 11508 39732
rect 11452 39678 11454 39730
rect 11454 39678 11506 39730
rect 11506 39678 11508 39730
rect 11452 39676 11508 39678
rect 9884 38220 9940 38276
rect 9996 38444 10052 38500
rect 9772 38108 9828 38164
rect 9548 38050 9604 38052
rect 9548 37998 9550 38050
rect 9550 37998 9602 38050
rect 9602 37998 9604 38050
rect 9548 37996 9604 37998
rect 9212 37660 9268 37716
rect 8428 36876 8484 36932
rect 8764 35922 8820 35924
rect 8764 35870 8766 35922
rect 8766 35870 8818 35922
rect 8818 35870 8820 35922
rect 8764 35868 8820 35870
rect 8316 34636 8372 34692
rect 8204 34130 8260 34132
rect 8204 34078 8206 34130
rect 8206 34078 8258 34130
rect 8258 34078 8260 34130
rect 8204 34076 8260 34078
rect 7420 33628 7476 33684
rect 7756 33852 7812 33908
rect 8764 33906 8820 33908
rect 8764 33854 8766 33906
rect 8766 33854 8818 33906
rect 8818 33854 8820 33906
rect 8764 33852 8820 33854
rect 9212 34636 9268 34692
rect 9100 33516 9156 33572
rect 8988 33292 9044 33348
rect 8764 32786 8820 32788
rect 8764 32734 8766 32786
rect 8766 32734 8818 32786
rect 8818 32734 8820 32786
rect 8764 32732 8820 32734
rect 3164 31778 3220 31780
rect 3164 31726 3166 31778
rect 3166 31726 3218 31778
rect 3218 31726 3220 31778
rect 3164 31724 3220 31726
rect 2380 31164 2436 31220
rect 4172 31164 4228 31220
rect 4060 30940 4116 30996
rect 2940 30268 2996 30324
rect 2828 30210 2884 30212
rect 2828 30158 2830 30210
rect 2830 30158 2882 30210
rect 2882 30158 2884 30210
rect 2828 30156 2884 30158
rect 4732 31052 4788 31108
rect 4284 30882 4340 30884
rect 4284 30830 4286 30882
rect 4286 30830 4338 30882
rect 4338 30830 4340 30882
rect 4284 30828 4340 30830
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4956 31164 5012 31220
rect 5124 30828 5180 30884
rect 4956 30322 5012 30324
rect 4956 30270 4958 30322
rect 4958 30270 5010 30322
rect 5010 30270 5012 30322
rect 4956 30268 5012 30270
rect 3948 30044 4004 30100
rect 3836 29596 3892 29652
rect 2940 28812 2996 28868
rect 2716 28476 2772 28532
rect 4732 29932 4788 29988
rect 5068 29820 5124 29876
rect 5404 31164 5460 31220
rect 5404 30994 5460 30996
rect 5404 30942 5406 30994
rect 5406 30942 5458 30994
rect 5458 30942 5460 30994
rect 5404 30940 5460 30942
rect 5684 31106 5740 31108
rect 5684 31054 5686 31106
rect 5686 31054 5738 31106
rect 5738 31054 5740 31106
rect 5684 31052 5740 31054
rect 5516 30828 5572 30884
rect 7084 31724 7140 31780
rect 5852 30940 5908 30996
rect 5292 30044 5348 30100
rect 5292 29708 5348 29764
rect 5740 30156 5796 30212
rect 6300 31164 6356 31220
rect 7532 32060 7588 32116
rect 9100 32060 9156 32116
rect 8540 31890 8596 31892
rect 8540 31838 8542 31890
rect 8542 31838 8594 31890
rect 8594 31838 8596 31890
rect 8540 31836 8596 31838
rect 7064 30994 7120 30996
rect 7064 30942 7066 30994
rect 7066 30942 7118 30994
rect 7118 30942 7120 30994
rect 7064 30940 7120 30942
rect 5628 29596 5684 29652
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4844 28700 4900 28756
rect 4060 28588 4116 28644
rect 3612 28476 3668 28532
rect 3836 27858 3892 27860
rect 3836 27806 3838 27858
rect 3838 27806 3890 27858
rect 3890 27806 3892 27858
rect 3836 27804 3892 27806
rect 4284 27804 4340 27860
rect 5964 28812 6020 28868
rect 5740 28754 5796 28756
rect 5740 28702 5742 28754
rect 5742 28702 5794 28754
rect 5794 28702 5796 28754
rect 5740 28700 5796 28702
rect 5292 28588 5348 28644
rect 5964 28252 6020 28308
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 6188 30268 6244 30324
rect 6300 30044 6356 30100
rect 6860 29820 6916 29876
rect 6972 30156 7028 30212
rect 6076 27692 6132 27748
rect 6188 28252 6244 28308
rect 4788 27020 4844 27076
rect 5628 27074 5684 27076
rect 5628 27022 5630 27074
rect 5630 27022 5682 27074
rect 5682 27022 5684 27074
rect 5628 27020 5684 27022
rect 2604 26796 2660 26852
rect 5404 26796 5460 26852
rect 1820 24668 1876 24724
rect 2268 24668 2324 24724
rect 5180 26290 5236 26292
rect 5180 26238 5182 26290
rect 5182 26238 5234 26290
rect 5234 26238 5236 26290
rect 5180 26236 5236 26238
rect 6636 29596 6692 29652
rect 6412 26572 6468 26628
rect 3164 26178 3220 26180
rect 3164 26126 3166 26178
rect 3166 26126 3218 26178
rect 3218 26126 3220 26178
rect 3164 26124 3220 26126
rect 3724 26124 3780 26180
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4508 25506 4564 25508
rect 4508 25454 4510 25506
rect 4510 25454 4562 25506
rect 4562 25454 4564 25506
rect 4508 25452 4564 25454
rect 5740 25340 5796 25396
rect 5404 25228 5460 25284
rect 4844 25004 4900 25060
rect 3500 24780 3556 24836
rect 3948 24834 4004 24836
rect 3948 24782 3950 24834
rect 3950 24782 4002 24834
rect 4002 24782 4004 24834
rect 3948 24780 4004 24782
rect 4564 24834 4620 24836
rect 4564 24782 4566 24834
rect 4566 24782 4618 24834
rect 4618 24782 4620 24834
rect 4564 24780 4620 24782
rect 2828 24722 2884 24724
rect 2828 24670 2830 24722
rect 2830 24670 2882 24722
rect 2882 24670 2884 24722
rect 2828 24668 2884 24670
rect 4956 24780 5012 24836
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 2492 23324 2548 23380
rect 2716 23154 2772 23156
rect 2716 23102 2718 23154
rect 2718 23102 2770 23154
rect 2770 23102 2772 23154
rect 2716 23100 2772 23102
rect 3612 23100 3668 23156
rect 2380 22204 2436 22260
rect 3444 22594 3500 22596
rect 3444 22542 3446 22594
rect 3446 22542 3498 22594
rect 3498 22542 3500 22594
rect 3444 22540 3500 22542
rect 3052 21756 3108 21812
rect 2604 20914 2660 20916
rect 2604 20862 2606 20914
rect 2606 20862 2658 20914
rect 2658 20862 2660 20914
rect 2604 20860 2660 20862
rect 2380 20802 2436 20804
rect 2380 20750 2382 20802
rect 2382 20750 2434 20802
rect 2434 20750 2436 20802
rect 2380 20748 2436 20750
rect 3276 21196 3332 21252
rect 3052 20972 3108 21028
rect 2716 20636 2772 20692
rect 3948 23436 4004 23492
rect 4284 23436 4340 23492
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 3836 22204 3892 22260
rect 4676 22258 4732 22260
rect 4676 22206 4678 22258
rect 4678 22206 4730 22258
rect 4730 22206 4732 22258
rect 4676 22204 4732 22206
rect 4172 22092 4228 22148
rect 3500 20748 3556 20804
rect 2380 19404 2436 19460
rect 3052 18508 3108 18564
rect 1596 18396 1652 18452
rect 2044 18450 2100 18452
rect 2044 18398 2046 18450
rect 2046 18398 2098 18450
rect 2098 18398 2100 18450
rect 2044 18396 2100 18398
rect 4284 21474 4340 21476
rect 4284 21422 4286 21474
rect 4286 21422 4338 21474
rect 4338 21422 4340 21474
rect 4284 21420 4340 21422
rect 5180 23436 5236 23492
rect 5068 22540 5124 22596
rect 5628 23436 5684 23492
rect 5348 23266 5404 23268
rect 5348 23214 5350 23266
rect 5350 23214 5402 23266
rect 5402 23214 5404 23266
rect 5348 23212 5404 23214
rect 5516 23212 5572 23268
rect 4956 22092 5012 22148
rect 5292 22204 5348 22260
rect 6188 26124 6244 26180
rect 5852 24780 5908 24836
rect 6076 25228 6132 25284
rect 4844 21420 4900 21476
rect 5180 21420 5236 21476
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4284 20972 4340 21028
rect 3724 20860 3780 20916
rect 4956 20636 5012 20692
rect 5852 22370 5908 22372
rect 5852 22318 5854 22370
rect 5854 22318 5906 22370
rect 5906 22318 5908 22370
rect 5852 22316 5908 22318
rect 6188 25004 6244 25060
rect 6412 25340 6468 25396
rect 7084 30044 7140 30100
rect 8316 30210 8372 30212
rect 8316 30158 8318 30210
rect 8318 30158 8370 30210
rect 8370 30158 8372 30210
rect 8316 30156 8372 30158
rect 7532 29932 7588 29988
rect 7196 29708 7252 29764
rect 9100 29820 9156 29876
rect 7868 29708 7924 29764
rect 9380 34690 9436 34692
rect 9380 34638 9382 34690
rect 9382 34638 9434 34690
rect 9434 34638 9436 34690
rect 9380 34636 9436 34638
rect 9604 34412 9660 34468
rect 10108 38108 10164 38164
rect 10612 38274 10668 38276
rect 10612 38222 10614 38274
rect 10614 38222 10666 38274
rect 10666 38222 10668 38274
rect 10612 38220 10668 38222
rect 11788 39340 11844 39396
rect 11788 39116 11844 39172
rect 10332 38050 10388 38052
rect 10332 37998 10334 38050
rect 10334 37998 10386 38050
rect 10386 37998 10388 38050
rect 10332 37996 10388 37998
rect 11676 37996 11732 38052
rect 12572 40572 12628 40628
rect 12012 39676 12068 39732
rect 12124 39004 12180 39060
rect 11900 37548 11956 37604
rect 12124 36988 12180 37044
rect 12796 40684 12852 40740
rect 13244 40684 13300 40740
rect 13468 42588 13524 42644
rect 13580 42700 13636 42756
rect 14588 43932 14644 43988
rect 14476 43596 14532 43652
rect 14476 43372 14532 43428
rect 15596 45164 15652 45220
rect 17612 45778 17668 45780
rect 17612 45726 17614 45778
rect 17614 45726 17666 45778
rect 17666 45726 17668 45778
rect 17612 45724 17668 45726
rect 17836 46508 17892 46564
rect 17724 45106 17780 45108
rect 17724 45054 17726 45106
rect 17726 45054 17778 45106
rect 17778 45054 17780 45106
rect 17724 45052 17780 45054
rect 18172 46396 18228 46452
rect 17948 45276 18004 45332
rect 18172 45388 18228 45444
rect 16828 44604 16884 44660
rect 15820 44434 15876 44436
rect 15820 44382 15822 44434
rect 15822 44382 15874 44434
rect 15874 44382 15876 44434
rect 15820 44380 15876 44382
rect 15372 44044 15428 44100
rect 16156 44044 16212 44100
rect 16268 44156 16324 44212
rect 15932 43932 15988 43988
rect 14924 43484 14980 43540
rect 16044 43484 16100 43540
rect 14476 42588 14532 42644
rect 16044 42700 16100 42756
rect 16156 43260 16212 43316
rect 15372 42588 15428 42644
rect 13692 41946 13694 41972
rect 13694 41946 13746 41972
rect 13746 41946 13748 41972
rect 13692 41916 13748 41946
rect 13916 41946 13918 41972
rect 13918 41946 13970 41972
rect 13970 41946 13972 41972
rect 13916 41916 13972 41946
rect 16268 42588 16324 42644
rect 16604 43596 16660 43652
rect 13468 41804 13524 41860
rect 13804 41153 13860 41188
rect 13804 41132 13806 41153
rect 13806 41132 13858 41153
rect 13858 41132 13860 41153
rect 15372 41916 15428 41972
rect 15708 41804 15764 41860
rect 16436 41970 16492 41972
rect 15596 41580 15652 41636
rect 16436 41918 16438 41970
rect 16438 41918 16490 41970
rect 16490 41918 16492 41970
rect 16436 41916 16492 41918
rect 15932 41356 15988 41412
rect 16156 41692 16212 41748
rect 12908 40402 12964 40404
rect 12908 40350 12910 40402
rect 12910 40350 12962 40402
rect 12962 40350 12964 40402
rect 12908 40348 12964 40350
rect 13020 40012 13076 40068
rect 12460 38892 12516 38948
rect 12348 38050 12404 38052
rect 12348 37998 12350 38050
rect 12350 37998 12402 38050
rect 12402 37998 12404 38050
rect 12348 37996 12404 37998
rect 12236 37436 12292 37492
rect 10780 36428 10836 36484
rect 10108 34914 10164 34916
rect 10108 34862 10110 34914
rect 10110 34862 10162 34914
rect 10162 34862 10164 34914
rect 10108 34860 10164 34862
rect 9996 34412 10052 34468
rect 9884 34076 9940 34132
rect 10556 35532 10612 35588
rect 10444 34412 10500 34468
rect 10164 33570 10220 33572
rect 10164 33518 10166 33570
rect 10166 33518 10218 33570
rect 10218 33518 10220 33570
rect 10164 33516 10220 33518
rect 10332 33516 10388 33572
rect 9996 33404 10052 33460
rect 9660 33346 9716 33348
rect 9660 33294 9662 33346
rect 9662 33294 9714 33346
rect 9714 33294 9716 33346
rect 9660 33292 9716 33294
rect 10444 33318 10500 33348
rect 10444 33292 10446 33318
rect 10446 33292 10498 33318
rect 10498 33292 10500 33318
rect 10332 32732 10388 32788
rect 7532 29260 7588 29316
rect 9212 29372 9268 29428
rect 9324 32508 9380 32564
rect 12460 37548 12516 37604
rect 12572 37324 12628 37380
rect 12572 36454 12628 36484
rect 12572 36428 12574 36454
rect 12574 36428 12626 36454
rect 12626 36428 12628 36454
rect 11116 35756 11172 35812
rect 10948 35586 11004 35588
rect 10948 35534 10950 35586
rect 10950 35534 11002 35586
rect 11002 35534 11004 35586
rect 10948 35532 11004 35534
rect 10892 34300 10948 34356
rect 11676 34636 11732 34692
rect 9996 32562 10052 32564
rect 9996 32510 9998 32562
rect 9998 32510 10050 32562
rect 10050 32510 10052 32562
rect 9996 32508 10052 32510
rect 11564 33516 11620 33572
rect 10668 33404 10724 33460
rect 9660 32172 9716 32228
rect 9772 32060 9828 32116
rect 8540 29260 8596 29316
rect 6972 28642 7028 28644
rect 6972 28590 6974 28642
rect 6974 28590 7026 28642
rect 7026 28590 7028 28642
rect 6972 28588 7028 28590
rect 6748 27858 6804 27860
rect 6748 27806 6750 27858
rect 6750 27806 6802 27858
rect 6802 27806 6804 27858
rect 6748 27804 6804 27806
rect 7252 28252 7308 28308
rect 9212 28700 9268 28756
rect 7980 28588 8036 28644
rect 7084 27858 7140 27860
rect 7084 27806 7086 27858
rect 7086 27806 7138 27858
rect 7138 27806 7140 27858
rect 8988 27916 9044 27972
rect 7084 27804 7140 27806
rect 10108 31778 10164 31780
rect 10108 31726 10110 31778
rect 10110 31726 10162 31778
rect 10162 31726 10164 31778
rect 10108 31724 10164 31726
rect 9548 29820 9604 29876
rect 9660 29484 9716 29540
rect 9996 29260 10052 29316
rect 11004 33180 11060 33236
rect 10892 32732 10948 32788
rect 14476 40402 14532 40404
rect 14476 40350 14478 40402
rect 14478 40350 14530 40402
rect 14530 40350 14532 40402
rect 14476 40348 14532 40350
rect 14252 40236 14308 40292
rect 14812 40684 14868 40740
rect 15372 40348 15428 40404
rect 15820 41020 15876 41076
rect 16716 43538 16772 43540
rect 16716 43486 16718 43538
rect 16718 43486 16770 43538
rect 16770 43486 16772 43538
rect 16716 43484 16772 43486
rect 16604 41580 16660 41636
rect 16492 41186 16548 41188
rect 16492 41134 16494 41186
rect 16494 41134 16546 41186
rect 16546 41134 16548 41186
rect 16492 41132 16548 41134
rect 17444 44604 17500 44660
rect 17948 45052 18004 45108
rect 16940 44268 16996 44324
rect 17052 43484 17108 43540
rect 18396 45724 18452 45780
rect 17612 43708 17668 43764
rect 17276 43538 17332 43540
rect 17276 43486 17278 43538
rect 17278 43486 17330 43538
rect 17330 43486 17332 43538
rect 17276 43484 17332 43486
rect 16044 40572 16100 40628
rect 16156 40796 16212 40852
rect 15036 39676 15092 39732
rect 16492 39900 16548 39956
rect 14812 39564 14868 39620
rect 14924 39452 14980 39508
rect 13580 38780 13636 38836
rect 15762 39618 15818 39620
rect 15762 39566 15764 39618
rect 15764 39566 15816 39618
rect 15816 39566 15818 39618
rect 15762 39564 15818 39566
rect 15484 39452 15540 39508
rect 17108 41186 17164 41188
rect 17108 41134 17110 41186
rect 17110 41134 17162 41186
rect 17162 41134 17164 41186
rect 17108 41132 17164 41134
rect 17276 43260 17332 43316
rect 17500 42476 17556 42532
rect 18396 45276 18452 45332
rect 18060 44294 18116 44324
rect 18060 44268 18062 44294
rect 18062 44268 18114 44294
rect 18114 44268 18116 44294
rect 18396 44268 18452 44324
rect 18284 44044 18340 44100
rect 17780 43314 17836 43316
rect 17780 43262 17782 43314
rect 17782 43262 17834 43314
rect 17834 43262 17836 43314
rect 17780 43260 17836 43262
rect 17948 42754 18004 42756
rect 17948 42702 17950 42754
rect 17950 42702 18002 42754
rect 18002 42702 18004 42754
rect 17948 42700 18004 42702
rect 18060 42588 18116 42644
rect 17500 41804 17556 41860
rect 17388 41580 17444 41636
rect 17500 41410 17556 41412
rect 17500 41358 17502 41410
rect 17502 41358 17554 41410
rect 17554 41358 17556 41410
rect 17500 41356 17556 41358
rect 18396 43708 18452 43764
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 18676 43820 18732 43876
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 20188 45276 20244 45332
rect 21084 47516 21140 47572
rect 20524 44380 20580 44436
rect 19964 44294 20020 44324
rect 19964 44268 19966 44294
rect 19966 44268 20018 44294
rect 20018 44268 20020 44294
rect 19628 44044 19684 44100
rect 18396 43036 18452 43092
rect 18228 41746 18284 41748
rect 18228 41694 18230 41746
rect 18230 41694 18282 41746
rect 18282 41694 18284 41746
rect 18228 41692 18284 41694
rect 18116 40962 18172 40964
rect 18116 40910 18118 40962
rect 18118 40910 18170 40962
rect 18170 40910 18172 40962
rect 18116 40908 18172 40910
rect 17276 40796 17332 40852
rect 17724 40402 17780 40404
rect 17724 40350 17726 40402
rect 17726 40350 17778 40402
rect 17778 40350 17780 40402
rect 17724 40348 17780 40350
rect 16716 39676 16772 39732
rect 15708 39340 15764 39396
rect 15372 38892 15428 38948
rect 14644 38780 14700 38836
rect 14812 38332 14868 38388
rect 15484 38834 15540 38836
rect 15484 38782 15486 38834
rect 15486 38782 15538 38834
rect 15538 38782 15540 38834
rect 15484 38780 15540 38782
rect 15876 38892 15932 38948
rect 18172 39004 18228 39060
rect 16828 38892 16884 38948
rect 15596 38668 15652 38724
rect 16548 38668 16604 38724
rect 15260 38108 15316 38164
rect 15820 38332 15876 38388
rect 12908 37436 12964 37492
rect 15820 37212 15876 37268
rect 15932 38108 15988 38164
rect 12236 34748 12292 34804
rect 12236 34354 12292 34356
rect 12236 34302 12238 34354
rect 12238 34302 12290 34354
rect 12290 34302 12292 34354
rect 12236 34300 12292 34302
rect 11900 33180 11956 33236
rect 12460 33180 12516 33236
rect 12684 35308 12740 35364
rect 12908 35308 12964 35364
rect 12796 34802 12852 34804
rect 12796 34750 12798 34802
rect 12798 34750 12850 34802
rect 12850 34750 12852 34802
rect 12796 34748 12852 34750
rect 12684 34636 12740 34692
rect 12908 34636 12964 34692
rect 13356 34412 13412 34468
rect 13020 34130 13076 34132
rect 13020 34078 13022 34130
rect 13022 34078 13074 34130
rect 13074 34078 13076 34130
rect 13020 34076 13076 34078
rect 12684 33404 12740 33460
rect 12908 33740 12964 33796
rect 12796 33331 12852 33348
rect 12796 33292 12798 33331
rect 12798 33292 12850 33331
rect 12850 33292 12852 33331
rect 11676 32732 11732 32788
rect 10668 32172 10724 32228
rect 10332 32060 10388 32116
rect 10612 31724 10668 31780
rect 11247 31778 11303 31780
rect 11247 31726 11249 31778
rect 11249 31726 11301 31778
rect 11301 31726 11303 31778
rect 11247 31724 11303 31726
rect 10668 30268 10724 30324
rect 10444 29538 10500 29540
rect 10444 29486 10446 29538
rect 10446 29486 10498 29538
rect 10498 29486 10500 29538
rect 10444 29484 10500 29486
rect 9996 28700 10052 28756
rect 10220 28812 10276 28868
rect 10220 28588 10276 28644
rect 9324 27804 9380 27860
rect 6972 26572 7028 26628
rect 6860 26178 6916 26180
rect 6860 26126 6862 26178
rect 6862 26126 6914 26178
rect 6914 26126 6916 26178
rect 6860 26124 6916 26126
rect 6636 25340 6692 25396
rect 8316 26796 8372 26852
rect 9884 27916 9940 27972
rect 9660 26908 9716 26964
rect 10108 27132 10164 27188
rect 9996 26290 10052 26292
rect 9996 26238 9998 26290
rect 9998 26238 10050 26290
rect 10050 26238 10052 26290
rect 9996 26236 10052 26238
rect 10276 26796 10332 26852
rect 10444 26460 10500 26516
rect 7196 25228 7252 25284
rect 7980 25506 8036 25508
rect 7980 25454 7982 25506
rect 7982 25454 8034 25506
rect 8034 25454 8036 25506
rect 7980 25452 8036 25454
rect 6524 25004 6580 25060
rect 6300 24892 6356 24948
rect 7308 24892 7364 24948
rect 8316 25506 8372 25508
rect 8316 25454 8318 25506
rect 8318 25454 8370 25506
rect 8370 25454 8372 25506
rect 8316 25452 8372 25454
rect 12124 31500 12180 31556
rect 11676 31388 11732 31444
rect 11004 30210 11060 30212
rect 11004 30158 11006 30210
rect 11006 30158 11058 30210
rect 11058 30158 11060 30210
rect 11004 30156 11060 30158
rect 12796 31778 12852 31780
rect 12796 31726 12798 31778
rect 12798 31726 12850 31778
rect 12850 31726 12852 31778
rect 12796 31724 12852 31726
rect 12516 31666 12572 31668
rect 12516 31614 12518 31666
rect 12518 31614 12570 31666
rect 12570 31614 12572 31666
rect 12516 31612 12572 31614
rect 12348 31388 12404 31444
rect 12516 31106 12572 31108
rect 12516 31054 12518 31106
rect 12518 31054 12570 31106
rect 12570 31054 12572 31106
rect 12516 31052 12572 31054
rect 12684 30828 12740 30884
rect 11676 30268 11732 30324
rect 12236 30210 12292 30212
rect 12236 30158 12238 30210
rect 12238 30158 12290 30210
rect 12290 30158 12292 30210
rect 12236 30156 12292 30158
rect 11452 29932 11508 29988
rect 12796 29820 12852 29876
rect 11564 29036 11620 29092
rect 11396 28866 11452 28868
rect 11396 28814 11398 28866
rect 11398 28814 11450 28866
rect 11450 28814 11452 28866
rect 11396 28812 11452 28814
rect 11340 27356 11396 27412
rect 10892 27020 10948 27076
rect 11116 26572 11172 26628
rect 11228 26460 11284 26516
rect 11228 26178 11284 26180
rect 11228 26126 11230 26178
rect 11230 26126 11282 26178
rect 11282 26126 11284 26178
rect 11228 26124 11284 26126
rect 6636 23212 6692 23268
rect 9100 24722 9156 24724
rect 9100 24670 9102 24722
rect 9102 24670 9154 24722
rect 9154 24670 9156 24722
rect 9100 24668 9156 24670
rect 10164 24722 10220 24724
rect 10164 24670 10166 24722
rect 10166 24670 10218 24722
rect 10218 24670 10220 24722
rect 10164 24668 10220 24670
rect 10668 25116 10724 25172
rect 10892 25004 10948 25060
rect 11004 24780 11060 24836
rect 11116 23772 11172 23828
rect 6860 23129 6862 23156
rect 6862 23129 6914 23156
rect 6914 23129 6916 23156
rect 6860 23100 6916 23129
rect 5628 21084 5684 21140
rect 4956 20076 5012 20132
rect 3612 19964 3668 20020
rect 4732 20018 4788 20020
rect 4732 19966 4734 20018
rect 4734 19966 4786 20018
rect 4786 19966 4788 20018
rect 4732 19964 4788 19966
rect 3836 18844 3892 18900
rect 3500 18284 3556 18340
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4732 19292 4788 19348
rect 4284 18508 4340 18564
rect 4060 18396 4116 18452
rect 4508 18284 4564 18340
rect 4396 18172 4452 18228
rect 3948 17052 4004 17108
rect 3388 16268 3444 16324
rect 2828 16098 2884 16100
rect 2828 16046 2830 16098
rect 2830 16046 2882 16098
rect 2882 16046 2884 16098
rect 2828 16044 2884 16046
rect 3164 15932 3220 15988
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 5404 20018 5460 20020
rect 5404 19966 5406 20018
rect 5406 19966 5458 20018
rect 5458 19966 5460 20018
rect 5404 19964 5460 19966
rect 6468 20972 6524 21028
rect 5908 20188 5964 20244
rect 5740 19964 5796 20020
rect 6188 20188 6244 20244
rect 5292 19404 5348 19460
rect 5628 19346 5684 19348
rect 5628 19294 5630 19346
rect 5630 19294 5682 19346
rect 5682 19294 5684 19346
rect 5628 19292 5684 19294
rect 5068 18844 5124 18900
rect 4844 17948 4900 18004
rect 4284 17666 4340 17668
rect 4284 17614 4286 17666
rect 4286 17614 4338 17666
rect 4338 17614 4340 17666
rect 4284 17612 4340 17614
rect 4284 17052 4340 17108
rect 4172 16828 4228 16884
rect 5460 18226 5516 18228
rect 5460 18174 5462 18226
rect 5462 18174 5514 18226
rect 5514 18174 5516 18226
rect 5460 18172 5516 18174
rect 5740 18172 5796 18228
rect 6636 20300 6692 20356
rect 5180 17836 5236 17892
rect 5516 17836 5572 17892
rect 5404 17500 5460 17556
rect 5180 17388 5236 17444
rect 5068 16857 5070 16884
rect 5070 16857 5122 16884
rect 5122 16857 5124 16884
rect 5068 16828 5124 16857
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4732 16268 4788 16324
rect 3500 15708 3556 15764
rect 4284 15932 4340 15988
rect 2828 15314 2884 15316
rect 2828 15262 2830 15314
rect 2830 15262 2882 15314
rect 2882 15262 2884 15314
rect 2828 15260 2884 15262
rect 4620 15932 4676 15988
rect 4620 15708 4676 15764
rect 4620 15260 4676 15316
rect 5404 16268 5460 16324
rect 5292 16044 5348 16100
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 5180 14364 5236 14420
rect 6412 20076 6468 20132
rect 6076 18284 6132 18340
rect 5964 17724 6020 17780
rect 6300 18060 6356 18116
rect 5740 17612 5796 17668
rect 5908 17554 5964 17556
rect 5908 17502 5910 17554
rect 5910 17502 5962 17554
rect 5962 17502 5964 17554
rect 5908 17500 5964 17502
rect 9660 23378 9716 23380
rect 9660 23326 9662 23378
rect 9662 23326 9714 23378
rect 9714 23326 9716 23378
rect 9660 23324 9716 23326
rect 10836 23154 10892 23156
rect 10836 23102 10838 23154
rect 10838 23102 10890 23154
rect 10890 23102 10892 23154
rect 10836 23100 10892 23102
rect 10892 22876 10948 22932
rect 7868 22316 7924 22372
rect 8876 22370 8932 22372
rect 8876 22318 8878 22370
rect 8878 22318 8930 22370
rect 8930 22318 8932 22370
rect 8876 22316 8932 22318
rect 7084 21084 7140 21140
rect 6860 20188 6916 20244
rect 6972 20972 7028 21028
rect 7700 21026 7756 21028
rect 7700 20974 7702 21026
rect 7702 20974 7754 21026
rect 7754 20974 7756 21026
rect 7700 20972 7756 20974
rect 7868 20802 7924 20804
rect 7868 20750 7870 20802
rect 7870 20750 7922 20802
rect 7922 20750 7924 20802
rect 7868 20748 7924 20750
rect 8092 20748 8148 20804
rect 6524 18396 6580 18452
rect 6636 17948 6692 18004
rect 7084 18172 7140 18228
rect 6972 17836 7028 17892
rect 6524 17724 6580 17780
rect 5852 17052 5908 17108
rect 5964 16940 6020 16996
rect 6132 16828 6188 16884
rect 6636 17052 6692 17108
rect 6972 17276 7028 17332
rect 7308 20188 7364 20244
rect 7756 20004 7758 20020
rect 7758 20004 7810 20020
rect 7810 20004 7812 20020
rect 7756 19964 7812 20004
rect 8540 20748 8596 20804
rect 9324 20802 9380 20804
rect 9324 20750 9326 20802
rect 9326 20750 9378 20802
rect 9378 20750 9380 20802
rect 9324 20748 9380 20750
rect 8820 20242 8876 20244
rect 8820 20190 8822 20242
rect 8822 20190 8874 20242
rect 8874 20190 8876 20242
rect 8820 20188 8876 20190
rect 7644 18172 7700 18228
rect 8316 17724 8372 17780
rect 6748 16770 6804 16772
rect 6748 16718 6750 16770
rect 6750 16718 6802 16770
rect 6802 16718 6804 16770
rect 6748 16716 6804 16718
rect 6300 15932 6356 15988
rect 8988 17778 9044 17780
rect 8988 17726 8990 17778
rect 8990 17726 9042 17778
rect 9042 17726 9044 17778
rect 8988 17724 9044 17726
rect 8876 17612 8932 17668
rect 7420 16940 7476 16996
rect 8540 17052 8596 17108
rect 8204 16716 8260 16772
rect 6412 15202 6468 15204
rect 6412 15150 6414 15202
rect 6414 15150 6466 15202
rect 6466 15150 6468 15202
rect 6412 15148 6468 15150
rect 5964 14812 6020 14868
rect 7084 16604 7140 16660
rect 6972 15314 7028 15316
rect 6972 15262 6974 15314
rect 6974 15262 7026 15314
rect 7026 15262 7028 15314
rect 6972 15260 7028 15262
rect 6860 15148 6916 15204
rect 9100 17388 9156 17444
rect 10220 22092 10276 22148
rect 12684 29148 12740 29204
rect 12348 28812 12404 28868
rect 11676 28642 11732 28644
rect 11676 28590 11678 28642
rect 11678 28590 11730 28642
rect 11730 28590 11732 28642
rect 11676 28588 11732 28590
rect 12236 28627 12292 28644
rect 12236 28588 12238 28627
rect 12238 28588 12290 28627
rect 12290 28588 12292 28627
rect 11900 28476 11956 28532
rect 11676 27468 11732 27524
rect 12460 28476 12516 28532
rect 13020 32508 13076 32564
rect 13244 32284 13300 32340
rect 14252 35420 14308 35476
rect 15372 36428 15428 36484
rect 15148 35308 15204 35364
rect 14924 35196 14980 35252
rect 16044 38050 16100 38052
rect 16044 37998 16046 38050
rect 16046 37998 16098 38050
rect 16098 37998 16100 38050
rect 16044 37996 16100 37998
rect 16940 38556 16996 38612
rect 17500 38108 17556 38164
rect 17388 38015 17444 38052
rect 17388 37996 17390 38015
rect 17390 37996 17442 38015
rect 17442 37996 17444 38015
rect 17948 38556 18004 38612
rect 17948 38220 18004 38276
rect 18956 43036 19012 43092
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 20076 42140 20132 42196
rect 18620 41970 18676 41972
rect 18620 41918 18622 41970
rect 18622 41918 18674 41970
rect 18674 41918 18676 41970
rect 18620 41916 18676 41918
rect 18788 41356 18844 41412
rect 22428 47570 22484 47572
rect 22428 47518 22430 47570
rect 22430 47518 22482 47570
rect 22482 47518 22484 47570
rect 22428 47516 22484 47518
rect 22764 47458 22820 47460
rect 22764 47406 22766 47458
rect 22766 47406 22818 47458
rect 22818 47406 22820 47458
rect 22764 47404 22820 47406
rect 21196 45052 21252 45108
rect 21308 45276 21364 45332
rect 23268 47234 23324 47236
rect 23268 47182 23270 47234
rect 23270 47182 23322 47234
rect 23322 47182 23324 47234
rect 23268 47180 23324 47182
rect 24892 47458 24948 47460
rect 24892 47406 24894 47458
rect 24894 47406 24946 47458
rect 24946 47406 24948 47458
rect 24892 47404 24948 47406
rect 23884 47180 23940 47236
rect 20748 44604 20804 44660
rect 20748 44380 20804 44436
rect 21532 44380 21588 44436
rect 22764 45276 22820 45332
rect 21084 44268 21140 44324
rect 20636 44044 20692 44100
rect 20636 43708 20692 43764
rect 20748 43372 20804 43428
rect 20636 42700 20692 42756
rect 20636 42140 20692 42196
rect 21028 43426 21084 43428
rect 21028 43374 21030 43426
rect 21030 43374 21082 43426
rect 21082 43374 21084 43426
rect 21028 43372 21084 43374
rect 21196 42754 21252 42756
rect 21196 42702 21198 42754
rect 21198 42702 21250 42754
rect 21250 42702 21252 42754
rect 21196 42700 21252 42702
rect 22764 44716 22820 44772
rect 21644 44044 21700 44100
rect 21532 43538 21588 43540
rect 21532 43486 21534 43538
rect 21534 43486 21586 43538
rect 21586 43486 21588 43538
rect 21532 43484 21588 43486
rect 21364 42530 21420 42532
rect 21364 42478 21366 42530
rect 21366 42478 21418 42530
rect 21418 42478 21420 42530
rect 21364 42476 21420 42478
rect 19068 40796 19124 40852
rect 19292 39788 19348 39844
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19964 40348 20020 40404
rect 19404 39618 19460 39620
rect 19404 39566 19406 39618
rect 19406 39566 19458 39618
rect 19458 39566 19460 39618
rect 19404 39564 19460 39566
rect 20524 41132 20580 41188
rect 20356 40962 20412 40964
rect 20356 40910 20358 40962
rect 20358 40910 20410 40962
rect 20410 40910 20412 40962
rect 20356 40908 20412 40910
rect 20748 40514 20804 40516
rect 20748 40462 20750 40514
rect 20750 40462 20802 40514
rect 20802 40462 20804 40514
rect 20748 40460 20804 40462
rect 18508 39394 18564 39396
rect 18508 39342 18510 39394
rect 18510 39342 18562 39394
rect 18562 39342 18564 39394
rect 18508 39340 18564 39342
rect 19068 39506 19124 39508
rect 19068 39454 19070 39506
rect 19070 39454 19122 39506
rect 19122 39454 19124 39506
rect 19068 39452 19124 39454
rect 20188 39452 20244 39508
rect 20300 39564 20356 39620
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 18620 38108 18676 38164
rect 19964 38668 20020 38724
rect 20524 39452 20580 39508
rect 20412 39340 20468 39396
rect 20860 39340 20916 39396
rect 21084 39452 21140 39508
rect 21196 41244 21252 41300
rect 21420 41132 21476 41188
rect 20972 39228 21028 39284
rect 21308 39228 21364 39284
rect 20972 39004 21028 39060
rect 20300 38668 20356 38724
rect 20860 38722 20916 38724
rect 20860 38670 20862 38722
rect 20862 38670 20914 38722
rect 20914 38670 20916 38722
rect 20860 38668 20916 38670
rect 18844 38108 18900 38164
rect 17500 37378 17556 37380
rect 17500 37326 17502 37378
rect 17502 37326 17554 37378
rect 17554 37326 17556 37378
rect 17500 37324 17556 37326
rect 17743 37324 17799 37380
rect 18396 38050 18452 38052
rect 18396 37998 18398 38050
rect 18398 37998 18450 38050
rect 18450 37998 18452 38050
rect 18396 37996 18452 37998
rect 18620 37436 18676 37492
rect 17948 37324 18004 37380
rect 17836 36988 17892 37044
rect 16716 36454 16772 36484
rect 16380 35532 16436 35588
rect 16716 36428 16718 36454
rect 16718 36428 16770 36454
rect 16770 36428 16772 36454
rect 16492 35868 16548 35924
rect 15932 35420 15988 35476
rect 17220 35756 17276 35812
rect 16492 35308 16548 35364
rect 16884 35308 16940 35364
rect 17500 35308 17556 35364
rect 15372 35196 15428 35252
rect 15260 34636 15316 34692
rect 13468 34076 13524 34132
rect 13804 33740 13860 33796
rect 13580 33346 13636 33348
rect 13580 33294 13582 33346
rect 13582 33294 13634 33346
rect 13634 33294 13636 33346
rect 13580 33292 13636 33294
rect 13580 33068 13636 33124
rect 14700 33068 14756 33124
rect 13804 32284 13860 32340
rect 14252 32620 14308 32676
rect 13132 31724 13188 31780
rect 13020 31612 13076 31668
rect 15148 33346 15204 33348
rect 15148 33294 15150 33346
rect 15150 33294 15202 33346
rect 15202 33294 15204 33346
rect 15148 33292 15204 33294
rect 16156 34636 16212 34692
rect 16492 34636 16548 34692
rect 15484 33068 15540 33124
rect 15708 32956 15764 33012
rect 15820 34076 15876 34132
rect 15036 32620 15092 32676
rect 14364 32537 14366 32564
rect 14366 32537 14418 32564
rect 14418 32537 14420 32564
rect 14364 32508 14420 32537
rect 15820 32508 15876 32564
rect 16380 33852 16436 33908
rect 16380 33180 16436 33236
rect 16268 32562 16324 32564
rect 16268 32510 16270 32562
rect 16270 32510 16322 32562
rect 16322 32510 16324 32562
rect 16268 32508 16324 32510
rect 13916 31612 13972 31668
rect 14476 31836 14532 31892
rect 13356 31388 13412 31444
rect 13020 30716 13076 30772
rect 11900 27356 11956 27412
rect 12460 27356 12516 27412
rect 11788 27074 11844 27076
rect 11788 27022 11790 27074
rect 11790 27022 11842 27074
rect 11842 27022 11844 27074
rect 11788 27020 11844 27022
rect 12852 27298 12908 27300
rect 12852 27246 12854 27298
rect 12854 27246 12906 27298
rect 12906 27246 12908 27298
rect 12852 27244 12908 27246
rect 12572 27074 12628 27076
rect 12572 27022 12574 27074
rect 12574 27022 12626 27074
rect 12626 27022 12628 27074
rect 12572 27020 12628 27022
rect 11956 26908 12012 26964
rect 11452 26460 11508 26516
rect 11508 26236 11564 26292
rect 11340 24668 11396 24724
rect 11788 26572 11844 26628
rect 12012 25116 12068 25172
rect 11676 24780 11732 24836
rect 12012 24892 12068 24948
rect 12348 25228 12404 25284
rect 12236 25116 12292 25172
rect 11676 23996 11732 24052
rect 12460 25004 12516 25060
rect 13356 30977 13358 30996
rect 13358 30977 13410 30996
rect 13410 30977 13412 30996
rect 13356 30940 13412 30977
rect 14028 31164 14084 31220
rect 15596 31612 15652 31668
rect 13524 30940 13580 30996
rect 13692 30828 13748 30884
rect 13244 30380 13300 30436
rect 13916 30716 13972 30772
rect 14588 30380 14644 30436
rect 13356 29148 13412 29204
rect 13244 28588 13300 28644
rect 13692 28642 13748 28644
rect 13692 28590 13694 28642
rect 13694 28590 13746 28642
rect 13746 28590 13748 28642
rect 13692 28588 13748 28590
rect 13468 27132 13524 27188
rect 13300 27020 13356 27076
rect 13804 27046 13860 27076
rect 13804 27020 13806 27046
rect 13806 27020 13858 27046
rect 13858 27020 13860 27046
rect 13580 26908 13636 26964
rect 13692 26460 13748 26516
rect 14924 31164 14980 31220
rect 14812 30994 14868 30996
rect 14812 30942 14814 30994
rect 14814 30942 14866 30994
rect 14866 30942 14868 30994
rect 14812 30940 14868 30942
rect 14084 30044 14140 30100
rect 14476 28588 14532 28644
rect 14364 27916 14420 27972
rect 14028 27858 14084 27860
rect 14028 27806 14030 27858
rect 14030 27806 14082 27858
rect 14082 27806 14084 27858
rect 14028 27804 14084 27806
rect 14028 27356 14084 27412
rect 15820 31164 15876 31220
rect 16044 31052 16100 31108
rect 15484 30492 15540 30548
rect 15148 30380 15204 30436
rect 15260 30044 15316 30100
rect 15372 29932 15428 29988
rect 15820 30044 15876 30100
rect 15708 29932 15764 29988
rect 15932 29426 15988 29428
rect 15932 29374 15934 29426
rect 15934 29374 15986 29426
rect 15986 29374 15988 29426
rect 15932 29372 15988 29374
rect 15260 29148 15316 29204
rect 16380 31948 16436 32004
rect 16772 34690 16828 34692
rect 16772 34638 16774 34690
rect 16774 34638 16826 34690
rect 16826 34638 16828 34690
rect 16772 34636 16828 34638
rect 16716 34188 16772 34244
rect 16940 34076 16996 34132
rect 17724 34860 17780 34916
rect 18620 37266 18676 37268
rect 18620 37214 18622 37266
rect 18622 37214 18674 37266
rect 18674 37214 18676 37266
rect 18620 37212 18676 37214
rect 19292 38050 19348 38052
rect 19292 37998 19294 38050
rect 19294 37998 19346 38050
rect 19346 37998 19348 38050
rect 19292 37996 19348 37998
rect 19124 37884 19180 37940
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20076 37436 20132 37492
rect 20300 37884 20356 37940
rect 18956 36988 19012 37044
rect 18396 35922 18452 35924
rect 18396 35870 18398 35922
rect 18398 35870 18450 35922
rect 18450 35870 18452 35922
rect 18396 35868 18452 35870
rect 17500 34242 17556 34244
rect 17500 34190 17502 34242
rect 17502 34190 17554 34242
rect 17554 34190 17556 34242
rect 17500 34188 17556 34190
rect 17743 34130 17799 34132
rect 17743 34078 17745 34130
rect 17745 34078 17797 34130
rect 17797 34078 17799 34130
rect 17743 34076 17799 34078
rect 17388 33740 17444 33796
rect 16492 32396 16548 32452
rect 16380 29484 16436 29540
rect 16716 31276 16772 31332
rect 16604 31218 16660 31220
rect 16604 31166 16606 31218
rect 16606 31166 16658 31218
rect 16658 31166 16660 31218
rect 16604 31164 16660 31166
rect 17724 33292 17780 33348
rect 17388 33068 17444 33124
rect 16828 30604 16884 30660
rect 16716 30492 16772 30548
rect 16940 30380 16996 30436
rect 16940 29820 16996 29876
rect 16492 29372 16548 29428
rect 16828 29372 16884 29428
rect 14812 28642 14868 28644
rect 14812 28590 14814 28642
rect 14814 28590 14866 28642
rect 14866 28590 14868 28642
rect 16268 28700 16324 28756
rect 14812 28588 14868 28590
rect 15932 28642 15988 28644
rect 15932 28590 15934 28642
rect 15934 28590 15986 28642
rect 15986 28590 15988 28642
rect 15932 28588 15988 28590
rect 14812 28140 14868 28196
rect 15036 28140 15092 28196
rect 15036 27916 15092 27972
rect 14700 27244 14756 27300
rect 15148 27356 15204 27412
rect 15596 27244 15652 27300
rect 15820 27244 15876 27300
rect 16044 27858 16100 27860
rect 16044 27806 16046 27858
rect 16046 27806 16098 27858
rect 16098 27806 16100 27858
rect 16044 27804 16100 27806
rect 16324 27356 16380 27412
rect 16268 26908 16324 26964
rect 16940 28866 16996 28868
rect 16940 28814 16942 28866
rect 16942 28814 16994 28866
rect 16994 28814 16996 28866
rect 16940 28812 16996 28814
rect 17164 32508 17220 32564
rect 17724 33068 17780 33124
rect 17836 33740 17892 33796
rect 18172 34802 18228 34804
rect 18172 34750 18174 34802
rect 18174 34750 18226 34802
rect 18226 34750 18228 34802
rect 18172 34748 18228 34750
rect 18060 34412 18116 34468
rect 20524 37660 20580 37716
rect 20748 38050 20804 38052
rect 20748 37998 20750 38050
rect 20750 37998 20802 38050
rect 20802 37998 20804 38050
rect 20748 37996 20804 37998
rect 20636 37212 20692 37268
rect 20972 37884 21028 37940
rect 19516 36428 19572 36484
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 18844 35756 18900 35812
rect 18732 35532 18788 35588
rect 20300 35698 20356 35700
rect 20300 35646 20302 35698
rect 20302 35646 20354 35698
rect 20354 35646 20356 35698
rect 20300 35644 20356 35646
rect 20076 35084 20132 35140
rect 18508 34188 18564 34244
rect 18620 34524 18676 34580
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 20804 36652 20860 36708
rect 20524 36092 20580 36148
rect 21868 43596 21924 43652
rect 21756 43484 21812 43540
rect 21644 42140 21700 42196
rect 22204 43596 22260 43652
rect 22092 43538 22148 43540
rect 22092 43486 22094 43538
rect 22094 43486 22146 43538
rect 22146 43486 22148 43538
rect 22092 43484 22148 43486
rect 23007 43596 23063 43652
rect 23436 44322 23492 44324
rect 23436 44270 23438 44322
rect 23438 44270 23490 44322
rect 23490 44270 23492 44322
rect 23436 44268 23492 44270
rect 24556 47180 24612 47236
rect 24668 47068 24724 47124
rect 25340 47068 25396 47124
rect 26628 47458 26684 47460
rect 26628 47406 26630 47458
rect 26630 47406 26682 47458
rect 26682 47406 26684 47458
rect 26628 47404 26684 47406
rect 23884 45052 23940 45108
rect 25228 45106 25284 45108
rect 25228 45054 25230 45106
rect 25230 45054 25282 45106
rect 25282 45054 25284 45106
rect 25228 45052 25284 45054
rect 23772 44380 23828 44436
rect 23660 44268 23716 44324
rect 24780 44434 24836 44436
rect 24780 44382 24782 44434
rect 24782 44382 24834 44434
rect 24834 44382 24836 44434
rect 24780 44380 24836 44382
rect 26348 45890 26404 45892
rect 26348 45838 26350 45890
rect 26350 45838 26402 45890
rect 26402 45838 26404 45890
rect 26348 45836 26404 45838
rect 27580 46674 27636 46676
rect 27580 46622 27582 46674
rect 27582 46622 27634 46674
rect 27634 46622 27636 46674
rect 27580 46620 27636 46622
rect 29240 47458 29296 47460
rect 29240 47406 29242 47458
rect 29242 47406 29294 47458
rect 29294 47406 29296 47458
rect 29240 47404 29296 47406
rect 30492 47404 30548 47460
rect 28364 46620 28420 46676
rect 29260 47180 29316 47236
rect 26684 45836 26740 45892
rect 27804 45890 27860 45892
rect 27804 45838 27806 45890
rect 27806 45838 27858 45890
rect 27858 45838 27860 45890
rect 27804 45836 27860 45838
rect 26684 45612 26740 45668
rect 25564 44380 25620 44436
rect 24220 43484 24276 43540
rect 22428 42140 22484 42196
rect 25228 44268 25284 44324
rect 22764 41970 22820 41972
rect 22764 41918 22766 41970
rect 22766 41918 22818 41970
rect 22818 41918 22820 41970
rect 22764 41916 22820 41918
rect 22540 41804 22596 41860
rect 21756 41244 21812 41300
rect 21868 41186 21924 41188
rect 21868 41134 21870 41186
rect 21870 41134 21922 41186
rect 21922 41134 21924 41186
rect 21868 41132 21924 41134
rect 21532 40908 21588 40964
rect 22316 40684 22372 40740
rect 22428 40572 22484 40628
rect 21980 40012 22036 40068
rect 21308 38050 21364 38052
rect 21308 37998 21310 38050
rect 21310 37998 21362 38050
rect 21362 37998 21364 38050
rect 21308 37996 21364 37998
rect 21420 37660 21476 37716
rect 21420 37266 21476 37268
rect 21420 37214 21422 37266
rect 21422 37214 21474 37266
rect 21474 37214 21476 37266
rect 21420 37212 21476 37214
rect 21644 37324 21700 37380
rect 20972 36428 21028 36484
rect 20804 35698 20860 35700
rect 20804 35646 20806 35698
rect 20806 35646 20858 35698
rect 20858 35646 20860 35698
rect 20804 35644 20860 35646
rect 21196 36092 21252 36148
rect 20972 35084 21028 35140
rect 19012 34130 19068 34132
rect 19012 34078 19014 34130
rect 19014 34078 19066 34130
rect 19066 34078 19068 34130
rect 19012 34076 19068 34078
rect 17948 33292 18004 33348
rect 18172 33628 18228 33684
rect 17388 31276 17444 31332
rect 17276 30604 17332 30660
rect 18508 33458 18564 33460
rect 18508 33406 18510 33458
rect 18510 33406 18562 33458
rect 18562 33406 18564 33458
rect 18508 33404 18564 33406
rect 19404 33516 19460 33572
rect 18284 31724 18340 31780
rect 18508 32562 18564 32564
rect 18508 32510 18510 32562
rect 18510 32510 18562 32562
rect 18562 32510 18564 32562
rect 18508 32508 18564 32510
rect 19236 33180 19292 33236
rect 20636 34130 20692 34132
rect 19740 33852 19796 33908
rect 20636 34078 20638 34130
rect 20638 34078 20690 34130
rect 20690 34078 20692 34130
rect 20636 34076 20692 34078
rect 20188 33404 20244 33460
rect 19740 33318 19796 33348
rect 19740 33292 19742 33318
rect 19742 33292 19794 33318
rect 19794 33292 19796 33318
rect 19964 33180 20020 33236
rect 20972 34018 21028 34020
rect 20972 33966 20974 34018
rect 20974 33966 21026 34018
rect 21026 33966 21028 34018
rect 20972 33964 21028 33966
rect 20860 33852 20916 33908
rect 19628 32956 19684 33012
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19404 32549 19406 32564
rect 19406 32549 19458 32564
rect 19458 32549 19460 32564
rect 19404 32508 19460 32549
rect 20300 33180 20356 33236
rect 19516 32284 19572 32340
rect 19180 32060 19236 32116
rect 20524 31948 20580 32004
rect 20188 31500 20244 31556
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 18620 31164 18676 31220
rect 17388 30492 17444 30548
rect 17836 30268 17892 30324
rect 17612 30210 17668 30212
rect 17612 30158 17614 30210
rect 17614 30158 17666 30210
rect 17666 30158 17668 30210
rect 17612 30156 17668 30158
rect 17052 27804 17108 27860
rect 17500 29820 17556 29876
rect 12852 25282 12908 25284
rect 12852 25230 12854 25282
rect 12854 25230 12906 25282
rect 12906 25230 12908 25282
rect 12852 25228 12908 25230
rect 12572 24892 12628 24948
rect 12236 23884 12292 23940
rect 12348 24332 12404 24388
rect 12460 23996 12516 24052
rect 11732 23826 11788 23828
rect 11732 23774 11734 23826
rect 11734 23774 11786 23826
rect 11786 23774 11788 23826
rect 11732 23772 11788 23774
rect 12572 23910 12628 23940
rect 12572 23884 12574 23910
rect 12574 23884 12626 23910
rect 12626 23884 12628 23910
rect 12796 23910 12852 23940
rect 12796 23884 12798 23910
rect 12798 23884 12850 23910
rect 12850 23884 12852 23910
rect 12908 23772 12964 23828
rect 11396 23266 11452 23268
rect 11396 23214 11398 23266
rect 11398 23214 11450 23266
rect 11450 23214 11452 23266
rect 11396 23212 11452 23214
rect 11732 22930 11788 22932
rect 11732 22878 11734 22930
rect 11734 22878 11786 22930
rect 11786 22878 11788 22930
rect 11732 22876 11788 22878
rect 11228 22316 11284 22372
rect 11564 22370 11620 22372
rect 11564 22318 11566 22370
rect 11566 22318 11618 22370
rect 11618 22318 11620 22370
rect 11564 22316 11620 22318
rect 11396 21810 11452 21812
rect 11396 21758 11398 21810
rect 11398 21758 11450 21810
rect 11450 21758 11452 21810
rect 11396 21756 11452 21758
rect 11900 22316 11956 22372
rect 12068 22258 12124 22260
rect 12068 22206 12070 22258
rect 12070 22206 12122 22258
rect 12122 22206 12124 22258
rect 12068 22204 12124 22206
rect 12460 22428 12516 22484
rect 12348 22342 12404 22372
rect 12348 22316 12350 22342
rect 12350 22316 12402 22342
rect 12402 22316 12404 22342
rect 12796 22342 12852 22372
rect 12236 22092 12292 22148
rect 12796 22316 12798 22342
rect 12798 22316 12850 22342
rect 12850 22316 12852 22342
rect 13356 25228 13412 25284
rect 13244 25004 13300 25060
rect 13244 23884 13300 23940
rect 13132 23772 13188 23828
rect 13804 25004 13860 25060
rect 15764 26460 15820 26516
rect 14364 26124 14420 26180
rect 16604 26460 16660 26516
rect 14140 25116 14196 25172
rect 13468 24332 13524 24388
rect 15260 25004 15316 25060
rect 14476 24780 14532 24836
rect 15596 24780 15652 24836
rect 14700 24722 14756 24724
rect 14700 24670 14702 24722
rect 14702 24670 14754 24722
rect 14754 24670 14756 24722
rect 14700 24668 14756 24670
rect 13916 24332 13972 24388
rect 13916 24108 13972 24164
rect 13580 24050 13636 24052
rect 13580 23998 13582 24050
rect 13582 23998 13634 24050
rect 13634 23998 13636 24050
rect 13580 23996 13636 23998
rect 13356 23436 13412 23492
rect 16660 26178 16716 26180
rect 16660 26126 16662 26178
rect 16662 26126 16714 26178
rect 16714 26126 16716 26178
rect 16660 26124 16716 26126
rect 17724 28588 17780 28644
rect 17052 25116 17108 25172
rect 17164 26460 17220 26516
rect 15988 24220 16044 24276
rect 13188 23378 13244 23380
rect 13188 23326 13190 23378
rect 13190 23326 13242 23378
rect 13242 23326 13244 23378
rect 13188 23324 13244 23326
rect 13916 23324 13972 23380
rect 14252 23436 14308 23492
rect 12572 22092 12628 22148
rect 12348 21980 12404 22036
rect 11844 21474 11900 21476
rect 11844 21422 11846 21474
rect 11846 21422 11898 21474
rect 11898 21422 11900 21474
rect 11844 21420 11900 21422
rect 12908 21756 12964 21812
rect 13020 23100 13076 23156
rect 12348 21420 12404 21476
rect 9660 20748 9716 20804
rect 11564 17778 11620 17780
rect 11564 17726 11566 17778
rect 11566 17726 11618 17778
rect 11618 17726 11620 17778
rect 11564 17724 11620 17726
rect 9548 17612 9604 17668
rect 9940 17666 9996 17668
rect 9940 17614 9942 17666
rect 9942 17614 9994 17666
rect 9994 17614 9996 17666
rect 9940 17612 9996 17614
rect 9324 17052 9380 17108
rect 11452 17651 11508 17668
rect 11452 17612 11454 17651
rect 11454 17612 11506 17651
rect 11506 17612 11508 17651
rect 12460 20748 12516 20804
rect 12572 20860 12628 20916
rect 12572 20188 12628 20244
rect 12684 20076 12740 20132
rect 14588 23212 14644 23268
rect 14252 22342 14308 22372
rect 14252 22316 14254 22342
rect 14254 22316 14306 22342
rect 14306 22316 14308 22342
rect 15988 23772 16044 23828
rect 14700 22876 14756 22932
rect 14588 22764 14644 22820
rect 15260 22652 15316 22708
rect 15484 23100 15540 23156
rect 14028 22092 14084 22148
rect 14364 21980 14420 22036
rect 13804 21868 13860 21924
rect 14588 21644 14644 21700
rect 14028 20860 14084 20916
rect 13356 20802 13412 20804
rect 13356 20750 13358 20802
rect 13358 20750 13410 20802
rect 13410 20750 13412 20802
rect 13356 20748 13412 20750
rect 13468 20076 13524 20132
rect 12460 19516 12516 19572
rect 13020 19794 13076 19796
rect 13020 19742 13022 19794
rect 13022 19742 13074 19794
rect 13074 19742 13076 19794
rect 13020 19740 13076 19742
rect 13916 19516 13972 19572
rect 11900 19180 11956 19236
rect 13356 19234 13412 19236
rect 13356 19182 13358 19234
rect 13358 19182 13410 19234
rect 13410 19182 13412 19234
rect 13356 19180 13412 19182
rect 13748 19068 13804 19124
rect 13524 19010 13580 19012
rect 13524 18958 13526 19010
rect 13526 18958 13578 19010
rect 13578 18958 13580 19010
rect 13524 18956 13580 18958
rect 11919 17948 11975 18004
rect 12796 18060 12852 18116
rect 12236 17724 12292 17780
rect 11900 17388 11956 17444
rect 12572 17500 12628 17556
rect 11228 17052 11284 17108
rect 8708 16994 8764 16996
rect 8708 16942 8710 16994
rect 8710 16942 8762 16994
rect 8762 16942 8764 16994
rect 8708 16940 8764 16942
rect 9436 16940 9492 16996
rect 6524 14812 6580 14868
rect 6076 14700 6132 14756
rect 5516 14364 5572 14420
rect 2548 13132 2604 13188
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4396 13132 4452 13188
rect 3724 12962 3780 12964
rect 3724 12910 3726 12962
rect 3726 12910 3778 12962
rect 3778 12910 3780 12962
rect 3724 12908 3780 12910
rect 2716 12348 2772 12404
rect 1596 12236 1652 12292
rect 2716 11394 2772 11396
rect 2716 11342 2718 11394
rect 2718 11342 2770 11394
rect 2770 11342 2772 11394
rect 2716 11340 2772 11342
rect 3388 11228 3444 11284
rect 3164 10780 3220 10836
rect 3948 11340 4004 11396
rect 4060 11228 4116 11284
rect 3724 9996 3780 10052
rect 2716 9826 2772 9828
rect 2716 9774 2718 9826
rect 2718 9774 2770 9826
rect 2770 9774 2772 9826
rect 2716 9772 2772 9774
rect 3612 9772 3668 9828
rect 2380 8316 2436 8372
rect 3388 8652 3444 8708
rect 4060 10556 4116 10612
rect 4284 12178 4340 12180
rect 4284 12126 4286 12178
rect 4286 12126 4338 12178
rect 4338 12126 4340 12178
rect 4284 12124 4340 12126
rect 4844 12012 4900 12068
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 6412 14700 6468 14756
rect 6300 14515 6356 14532
rect 6300 14476 6302 14515
rect 6302 14476 6354 14515
rect 6354 14476 6356 14515
rect 6972 14502 7028 14532
rect 6972 14476 6974 14502
rect 6974 14476 7026 14502
rect 7026 14476 7028 14502
rect 7084 14812 7140 14868
rect 7196 14700 7252 14756
rect 5292 13746 5348 13748
rect 5292 13694 5294 13746
rect 5294 13694 5346 13746
rect 5346 13694 5348 13746
rect 6748 14364 6804 14420
rect 6412 13746 6468 13748
rect 5292 13692 5348 13694
rect 6412 13694 6414 13746
rect 6414 13694 6466 13746
rect 6466 13694 6468 13746
rect 6412 13692 6468 13694
rect 5740 12908 5796 12964
rect 6076 13132 6132 13188
rect 5068 12124 5124 12180
rect 5180 12236 5236 12292
rect 4956 11900 5012 11956
rect 5180 11788 5236 11844
rect 5628 12124 5684 12180
rect 4284 10780 4340 10836
rect 4788 10610 4844 10612
rect 4788 10558 4790 10610
rect 4790 10558 4842 10610
rect 4842 10558 4844 10610
rect 4788 10556 4844 10558
rect 5404 10780 5460 10836
rect 5292 10668 5348 10724
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 3724 8652 3780 8708
rect 3612 8428 3668 8484
rect 4732 9884 4788 9940
rect 5628 10668 5684 10724
rect 5572 9996 5628 10052
rect 5964 10780 6020 10836
rect 5852 10610 5908 10612
rect 5852 10558 5854 10610
rect 5854 10558 5906 10610
rect 5906 10558 5908 10610
rect 5852 10556 5908 10558
rect 6300 12796 6356 12852
rect 6636 12796 6692 12852
rect 6412 12402 6468 12404
rect 6412 12350 6414 12402
rect 6414 12350 6466 12402
rect 6466 12350 6468 12402
rect 6412 12348 6468 12350
rect 6300 11394 6356 11396
rect 6300 11342 6302 11394
rect 6302 11342 6354 11394
rect 6354 11342 6356 11394
rect 6300 11340 6356 11342
rect 8036 15314 8092 15316
rect 8036 15262 8038 15314
rect 8038 15262 8090 15314
rect 8090 15262 8092 15314
rect 8036 15260 8092 15262
rect 9772 16658 9828 16660
rect 9772 16606 9774 16658
rect 9774 16606 9826 16658
rect 9826 16606 9828 16658
rect 9772 16604 9828 16606
rect 7420 14642 7476 14644
rect 7420 14590 7422 14642
rect 7422 14590 7474 14642
rect 7474 14590 7476 14642
rect 7420 14588 7476 14590
rect 8540 14642 8596 14644
rect 8540 14590 8542 14642
rect 8542 14590 8594 14642
rect 8594 14590 8596 14642
rect 8540 14588 8596 14590
rect 7756 14530 7812 14532
rect 7756 14478 7758 14530
rect 7758 14478 7810 14530
rect 7810 14478 7812 14530
rect 7756 14476 7812 14478
rect 6972 12962 7028 12964
rect 6972 12910 6974 12962
rect 6974 12910 7026 12962
rect 7026 12910 7028 12962
rect 6972 12908 7028 12910
rect 6748 11676 6804 11732
rect 6188 10668 6244 10724
rect 6300 10332 6356 10388
rect 5818 9212 5874 9268
rect 4900 8988 4956 9044
rect 5628 8988 5684 9044
rect 6692 10386 6748 10388
rect 6692 10334 6694 10386
rect 6694 10334 6746 10386
rect 6746 10334 6748 10386
rect 6692 10332 6748 10334
rect 7868 13746 7924 13748
rect 7868 13694 7870 13746
rect 7870 13694 7922 13746
rect 7922 13694 7924 13746
rect 7868 13692 7924 13694
rect 7812 13468 7868 13524
rect 9548 14812 9604 14868
rect 9772 15260 9828 15316
rect 9100 13746 9156 13748
rect 9100 13694 9102 13746
rect 9102 13694 9154 13746
rect 9154 13694 9156 13746
rect 9100 13692 9156 13694
rect 7532 12908 7588 12964
rect 8092 12796 8148 12852
rect 7532 12178 7588 12180
rect 7532 12126 7534 12178
rect 7534 12126 7586 12178
rect 7586 12126 7588 12178
rect 7532 12124 7588 12126
rect 7420 11900 7476 11956
rect 6412 9884 6468 9940
rect 6412 9660 6468 9716
rect 4284 8652 4340 8708
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4732 8428 4788 8484
rect 1596 7644 1652 7700
rect 2268 7644 2324 7700
rect 2828 6690 2884 6692
rect 2828 6638 2830 6690
rect 2830 6638 2882 6690
rect 2882 6638 2884 6690
rect 2828 6636 2884 6638
rect 3724 7644 3780 7700
rect 4956 8370 5012 8372
rect 4956 8318 4958 8370
rect 4958 8318 5010 8370
rect 5010 8318 5012 8370
rect 4956 8316 5012 8318
rect 6076 9042 6132 9044
rect 6076 8990 6078 9042
rect 6078 8990 6130 9042
rect 6130 8990 6132 9042
rect 6076 8988 6132 8990
rect 4004 7980 4060 8036
rect 4284 7980 4340 8036
rect 5852 7698 5908 7700
rect 5852 7646 5854 7698
rect 5854 7646 5906 7698
rect 5906 7646 5908 7698
rect 5852 7644 5908 7646
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4284 6860 4340 6916
rect 4956 6748 5012 6804
rect 3836 6524 3892 6580
rect 3612 6412 3668 6468
rect 5628 6412 5684 6468
rect 5740 6636 5796 6692
rect 5740 6188 5796 6244
rect 5628 6076 5684 6132
rect 4956 5906 5012 5908
rect 4956 5854 4958 5906
rect 4958 5854 5010 5906
rect 5010 5854 5012 5906
rect 4956 5852 5012 5854
rect 4620 5740 4676 5796
rect 3052 5628 3108 5684
rect 4396 5682 4452 5684
rect 4396 5630 4398 5682
rect 4398 5630 4450 5682
rect 4450 5630 4452 5682
rect 4396 5628 4452 5630
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4956 5234 5012 5236
rect 4956 5182 4958 5234
rect 4958 5182 5010 5234
rect 5010 5182 5012 5234
rect 4956 5180 5012 5182
rect 6076 6636 6132 6692
rect 5964 6524 6020 6580
rect 6300 6748 6356 6804
rect 6300 6300 6356 6356
rect 6580 9266 6636 9268
rect 6580 9214 6582 9266
rect 6582 9214 6634 9266
rect 6634 9214 6636 9266
rect 6580 9212 6636 9214
rect 7532 11394 7588 11396
rect 7532 11342 7534 11394
rect 7534 11342 7586 11394
rect 7586 11342 7588 11394
rect 7532 11340 7588 11342
rect 8316 12124 8372 12180
rect 8428 12348 8484 12404
rect 7924 12066 7980 12068
rect 7924 12014 7926 12066
rect 7926 12014 7978 12066
rect 7978 12014 7980 12066
rect 7924 12012 7980 12014
rect 8652 12012 8708 12068
rect 8540 11788 8596 11844
rect 7868 11676 7924 11732
rect 8204 11282 8260 11284
rect 8204 11230 8206 11282
rect 8206 11230 8258 11282
rect 8258 11230 8260 11282
rect 8204 11228 8260 11230
rect 7868 11116 7924 11172
rect 8092 10834 8148 10836
rect 8092 10782 8094 10834
rect 8094 10782 8146 10834
rect 8146 10782 8148 10834
rect 8092 10780 8148 10782
rect 8428 10610 8484 10612
rect 8428 10558 8430 10610
rect 8430 10558 8482 10610
rect 8482 10558 8484 10610
rect 8428 10556 8484 10558
rect 8402 9793 8458 9828
rect 7084 9266 7140 9268
rect 7084 9214 7086 9266
rect 7086 9214 7138 9266
rect 7138 9214 7140 9266
rect 7084 9212 7140 9214
rect 7420 9042 7476 9044
rect 7420 8990 7422 9042
rect 7422 8990 7474 9042
rect 7474 8990 7476 9042
rect 7420 8988 7476 8990
rect 8402 9772 8404 9793
rect 8404 9772 8456 9793
rect 8456 9772 8458 9793
rect 8092 9660 8148 9716
rect 7868 8988 7924 9044
rect 7756 8204 7812 8260
rect 7420 7644 7476 7700
rect 8204 7532 8260 7588
rect 7756 6972 7812 7028
rect 7084 6860 7140 6916
rect 6916 6636 6972 6692
rect 8092 7460 8094 7476
rect 8094 7460 8146 7476
rect 8146 7460 8148 7476
rect 8092 7420 8148 7460
rect 8092 6972 8148 7028
rect 6412 6188 6468 6244
rect 6860 6300 6916 6356
rect 6580 6076 6636 6132
rect 6076 5740 6132 5796
rect 5740 5180 5796 5236
rect 7868 6636 7924 6692
rect 7532 6300 7588 6356
rect 6972 5906 7028 5908
rect 6972 5854 6974 5906
rect 6974 5854 7026 5906
rect 7026 5854 7028 5906
rect 6972 5852 7028 5854
rect 8988 13244 9044 13300
rect 8876 12796 8932 12852
rect 9660 13692 9716 13748
rect 9884 14588 9940 14644
rect 10444 16604 10500 16660
rect 10892 16268 10948 16324
rect 11004 16716 11060 16772
rect 11676 16322 11732 16324
rect 11676 16270 11678 16322
rect 11678 16270 11730 16322
rect 11730 16270 11732 16322
rect 11676 16268 11732 16270
rect 11004 15820 11060 15876
rect 11004 15289 11006 15316
rect 11006 15289 11058 15316
rect 11058 15289 11060 15316
rect 11004 15260 11060 15289
rect 13356 18450 13412 18452
rect 13356 18398 13358 18450
rect 13358 18398 13410 18450
rect 13410 18398 13412 18450
rect 13356 18396 13412 18398
rect 14476 20748 14532 20804
rect 14194 19740 14250 19796
rect 15148 21868 15204 21924
rect 16604 23884 16660 23940
rect 16716 24444 16772 24500
rect 16996 24162 17052 24164
rect 16996 24110 16998 24162
rect 16998 24110 17050 24162
rect 17050 24110 17052 24162
rect 16996 24108 17052 24110
rect 17388 27244 17444 27300
rect 17836 28028 17892 28084
rect 18956 31052 19012 31108
rect 19124 31052 19180 31108
rect 18620 30828 18676 30884
rect 18844 30828 18900 30884
rect 19404 30994 19460 30996
rect 19404 30942 19406 30994
rect 19406 30942 19458 30994
rect 19458 30942 19460 30994
rect 19404 30940 19460 30942
rect 19628 30994 19684 30996
rect 19628 30942 19630 30994
rect 19630 30942 19682 30994
rect 19682 30942 19684 30994
rect 19628 30940 19684 30942
rect 20188 30940 20244 30996
rect 20860 31948 20916 32004
rect 20748 31612 20804 31668
rect 20412 31052 20468 31108
rect 18172 30156 18228 30212
rect 18396 30156 18452 30212
rect 20636 30828 20692 30884
rect 19068 30492 19124 30548
rect 19348 30380 19404 30436
rect 18284 30044 18340 30100
rect 18060 28924 18116 28980
rect 18060 28642 18116 28644
rect 18060 28590 18062 28642
rect 18062 28590 18114 28642
rect 18114 28590 18116 28642
rect 18060 28588 18116 28590
rect 18620 29932 18676 29988
rect 19908 30210 19964 30212
rect 19908 30158 19910 30210
rect 19910 30158 19962 30210
rect 19962 30158 19964 30210
rect 19908 30156 19964 30158
rect 18844 29820 18900 29876
rect 19292 29932 19348 29988
rect 18396 28924 18452 28980
rect 18508 28812 18564 28868
rect 18284 28028 18340 28084
rect 18060 27858 18116 27860
rect 18060 27806 18062 27858
rect 18062 27806 18114 27858
rect 18114 27806 18116 27858
rect 18060 27804 18116 27806
rect 18060 27580 18116 27636
rect 17612 27244 17668 27300
rect 17500 27132 17556 27188
rect 17388 26908 17444 26964
rect 17836 27244 17892 27300
rect 17500 26460 17556 26516
rect 17612 26684 17668 26740
rect 16380 23826 16436 23828
rect 16380 23774 16382 23826
rect 16382 23774 16434 23826
rect 16434 23774 16436 23826
rect 16380 23772 16436 23774
rect 16156 23100 16212 23156
rect 15596 22316 15652 22372
rect 16044 22092 16100 22148
rect 16268 21644 16324 21700
rect 14924 20748 14980 20804
rect 15932 20774 15988 20804
rect 15932 20748 15934 20774
rect 15934 20748 15986 20774
rect 15986 20748 15988 20774
rect 15328 20300 15384 20356
rect 16828 20300 16884 20356
rect 14700 20188 14756 20244
rect 16716 20018 16772 20020
rect 16716 19966 16718 20018
rect 16718 19966 16770 20018
rect 16770 19966 16772 20018
rect 16716 19964 16772 19966
rect 17276 23212 17332 23268
rect 17724 26012 17780 26068
rect 18340 27244 18396 27300
rect 20412 30492 20468 30548
rect 20076 29932 20132 29988
rect 19404 29820 19460 29876
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19628 29372 19684 29428
rect 19964 29426 20020 29428
rect 19964 29374 19966 29426
rect 19966 29374 20018 29426
rect 20018 29374 20020 29426
rect 19964 29372 20020 29374
rect 20524 30268 20580 30324
rect 20300 28700 20356 28756
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 18732 27804 18788 27860
rect 18956 27356 19012 27412
rect 20412 28028 20468 28084
rect 19628 27916 19684 27972
rect 21308 35084 21364 35140
rect 21644 35196 21700 35252
rect 21420 34748 21476 34804
rect 21420 34076 21476 34132
rect 22652 40908 22708 40964
rect 23212 41804 23268 41860
rect 23940 41746 23996 41748
rect 23940 41694 23942 41746
rect 23942 41694 23994 41746
rect 23994 41694 23996 41746
rect 23940 41692 23996 41694
rect 23548 41244 23604 41300
rect 23212 41020 23268 41076
rect 23324 41132 23380 41188
rect 25116 43596 25172 43652
rect 24948 42588 25004 42644
rect 24332 41916 24388 41972
rect 24556 41692 24612 41748
rect 24220 41020 24276 41076
rect 24108 40962 24164 40964
rect 24108 40910 24110 40962
rect 24110 40910 24162 40962
rect 24162 40910 24164 40962
rect 24108 40908 24164 40910
rect 23884 40572 23940 40628
rect 24332 40460 24388 40516
rect 23436 40402 23492 40404
rect 23436 40350 23438 40402
rect 23438 40350 23490 40402
rect 23490 40350 23492 40402
rect 23436 40348 23492 40350
rect 23100 39004 23156 39060
rect 22316 38668 22372 38724
rect 22316 38444 22372 38500
rect 22204 38220 22260 38276
rect 21980 37884 22036 37940
rect 22092 37996 22148 38052
rect 22316 38050 22372 38052
rect 22316 37998 22318 38050
rect 22318 37998 22370 38050
rect 22370 37998 22372 38050
rect 22316 37996 22372 37998
rect 22204 37212 22260 37268
rect 23436 39452 23492 39508
rect 23324 38780 23380 38836
rect 24444 40348 24500 40404
rect 24556 40684 24612 40740
rect 24668 40460 24724 40516
rect 24948 40348 25004 40404
rect 23772 38722 23828 38724
rect 23772 38670 23774 38722
rect 23774 38670 23826 38722
rect 23826 38670 23828 38722
rect 23772 38668 23828 38670
rect 23324 38220 23380 38276
rect 22652 36652 22708 36708
rect 22876 35644 22932 35700
rect 22876 35308 22932 35364
rect 23212 35308 23268 35364
rect 22204 35196 22260 35252
rect 21980 35084 22036 35140
rect 21756 34636 21812 34692
rect 21532 33516 21588 33572
rect 21644 33852 21700 33908
rect 23436 35308 23492 35364
rect 22652 33516 22708 33572
rect 21756 33122 21812 33124
rect 21756 33070 21758 33122
rect 21758 33070 21810 33122
rect 21810 33070 21812 33122
rect 21756 33068 21812 33070
rect 21532 32060 21588 32116
rect 21420 31890 21476 31892
rect 21420 31838 21422 31890
rect 21422 31838 21474 31890
rect 21474 31838 21476 31890
rect 21420 31836 21476 31838
rect 21308 31724 21364 31780
rect 21196 31164 21252 31220
rect 20860 31052 20916 31108
rect 21140 30994 21196 30996
rect 21140 30942 21142 30994
rect 21142 30942 21194 30994
rect 21194 30942 21196 30994
rect 21140 30940 21196 30942
rect 21196 30156 21252 30212
rect 21084 29484 21140 29540
rect 21812 31500 21868 31556
rect 22092 31612 22148 31668
rect 22540 33068 22596 33124
rect 22316 31948 22372 32004
rect 22652 32060 22708 32116
rect 22484 31724 22540 31780
rect 22876 33516 22932 33572
rect 23212 33311 23268 33348
rect 23212 33292 23214 33311
rect 23214 33292 23266 33311
rect 23266 33292 23268 33311
rect 25452 42978 25508 42980
rect 25452 42926 25454 42978
rect 25454 42926 25506 42978
rect 25506 42926 25508 42978
rect 25452 42924 25508 42926
rect 25788 42754 25844 42756
rect 25788 42702 25790 42754
rect 25790 42702 25842 42754
rect 25842 42702 25844 42754
rect 25788 42700 25844 42702
rect 26236 45052 26292 45108
rect 26012 42924 26068 42980
rect 25228 41970 25284 41972
rect 25228 41918 25230 41970
rect 25230 41918 25282 41970
rect 25282 41918 25284 41970
rect 25228 41916 25284 41918
rect 25900 41916 25956 41972
rect 25396 41746 25452 41748
rect 25396 41694 25398 41746
rect 25398 41694 25450 41746
rect 25450 41694 25452 41746
rect 25396 41692 25452 41694
rect 27356 45666 27412 45668
rect 27356 45614 27358 45666
rect 27358 45614 27410 45666
rect 27410 45614 27412 45666
rect 27356 45612 27412 45614
rect 27692 44044 27748 44100
rect 28252 44940 28308 44996
rect 28028 44716 28084 44772
rect 28252 44294 28308 44324
rect 28252 44268 28254 44294
rect 28254 44268 28306 44294
rect 28306 44268 28308 44294
rect 27916 44044 27972 44100
rect 28028 43932 28084 43988
rect 27468 43260 27524 43316
rect 27412 42754 27468 42756
rect 27412 42702 27414 42754
rect 27414 42702 27466 42754
rect 27466 42702 27468 42754
rect 27412 42700 27468 42702
rect 27692 42726 27748 42756
rect 27692 42700 27694 42726
rect 27694 42700 27746 42726
rect 27746 42700 27748 42726
rect 27916 43148 27972 43204
rect 26460 41970 26516 41972
rect 26460 41918 26462 41970
rect 26462 41918 26514 41970
rect 26514 41918 26516 41970
rect 26460 41916 26516 41918
rect 26236 41468 26292 41524
rect 25900 40908 25956 40964
rect 25564 40572 25620 40628
rect 25452 40402 25508 40404
rect 25452 40350 25454 40402
rect 25454 40350 25506 40402
rect 25506 40350 25508 40402
rect 25452 40348 25508 40350
rect 25116 39116 25172 39172
rect 23996 38444 24052 38500
rect 24444 38332 24500 38388
rect 23996 37772 24052 37828
rect 24220 37772 24276 37828
rect 23940 36988 23996 37044
rect 23660 36482 23716 36484
rect 23660 36430 23662 36482
rect 23662 36430 23714 36482
rect 23714 36430 23716 36482
rect 24444 36988 24500 37044
rect 24668 37884 24724 37940
rect 24668 36876 24724 36932
rect 25116 38834 25172 38836
rect 25116 38782 25118 38834
rect 25118 38782 25170 38834
rect 25170 38782 25172 38834
rect 25116 38780 25172 38782
rect 25788 38834 25844 38836
rect 25788 38782 25790 38834
rect 25790 38782 25842 38834
rect 25842 38782 25844 38834
rect 25788 38780 25844 38782
rect 25676 38668 25732 38724
rect 27916 41692 27972 41748
rect 27916 41158 27972 41188
rect 27916 41132 27918 41158
rect 27918 41132 27970 41158
rect 27970 41132 27972 41158
rect 26460 40908 26516 40964
rect 26124 40572 26180 40628
rect 26628 40348 26684 40404
rect 27636 40796 27692 40852
rect 30212 47234 30268 47236
rect 30212 47182 30214 47234
rect 30214 47182 30266 47234
rect 30266 47182 30268 47234
rect 30212 47180 30268 47182
rect 28588 44716 28644 44772
rect 28588 43484 28644 43540
rect 29036 44322 29092 44324
rect 29036 44270 29038 44322
rect 29038 44270 29090 44322
rect 29090 44270 29092 44322
rect 29036 44268 29092 44270
rect 29036 44044 29092 44100
rect 28140 43372 28196 43428
rect 28812 43372 28868 43428
rect 28252 43260 28308 43316
rect 28700 43148 28756 43204
rect 28476 41804 28532 41860
rect 28252 41356 28308 41412
rect 28140 41020 28196 41076
rect 28028 40572 28084 40628
rect 28252 40572 28308 40628
rect 28140 40514 28196 40516
rect 28140 40462 28142 40514
rect 28142 40462 28194 40514
rect 28194 40462 28196 40514
rect 28140 40460 28196 40462
rect 27692 40348 27748 40404
rect 26124 39058 26180 39060
rect 26124 39006 26126 39058
rect 26126 39006 26178 39058
rect 26178 39006 26180 39058
rect 26124 39004 26180 39006
rect 26796 40012 26852 40068
rect 26572 38668 26628 38724
rect 25004 38444 25060 38500
rect 26012 38332 26068 38388
rect 25004 37436 25060 37492
rect 25732 37660 25788 37716
rect 25732 37490 25788 37492
rect 25732 37438 25734 37490
rect 25734 37438 25786 37490
rect 25786 37438 25788 37490
rect 25732 37436 25788 37438
rect 26684 37548 26740 37604
rect 27692 39900 27748 39956
rect 27580 39788 27636 39844
rect 28476 40684 28532 40740
rect 28700 40684 28756 40740
rect 28476 39788 28532 39844
rect 28420 39618 28476 39620
rect 28420 39566 28422 39618
rect 28422 39566 28474 39618
rect 28474 39566 28476 39618
rect 28420 39564 28476 39566
rect 27580 38722 27636 38724
rect 27580 38670 27582 38722
rect 27582 38670 27634 38722
rect 27634 38670 27636 38722
rect 27580 38668 27636 38670
rect 27132 37548 27188 37604
rect 28364 39228 28420 39284
rect 23660 36428 23716 36430
rect 23772 36092 23828 36148
rect 23660 35420 23716 35476
rect 23884 33628 23940 33684
rect 23772 33516 23828 33572
rect 23772 33180 23828 33236
rect 23100 32732 23156 32788
rect 23660 32732 23716 32788
rect 23212 32060 23268 32116
rect 22932 32002 22988 32004
rect 22932 31950 22934 32002
rect 22934 31950 22986 32002
rect 22986 31950 22988 32002
rect 22932 31948 22988 31950
rect 22876 31724 22932 31780
rect 22316 30268 22372 30324
rect 22428 30994 22484 30996
rect 22428 30942 22430 30994
rect 22430 30942 22482 30994
rect 22482 30942 22484 30994
rect 22428 30940 22484 30942
rect 22540 30492 22596 30548
rect 22764 31052 22820 31108
rect 23436 31750 23492 31780
rect 23436 31724 23438 31750
rect 23438 31724 23490 31750
rect 23490 31724 23492 31750
rect 22988 30828 23044 30884
rect 26124 35980 26180 36036
rect 25116 35868 25172 35924
rect 25788 35922 25844 35924
rect 25788 35870 25790 35922
rect 25790 35870 25842 35922
rect 25842 35870 25844 35922
rect 25788 35868 25844 35870
rect 25396 35698 25452 35700
rect 25396 35646 25398 35698
rect 25398 35646 25450 35698
rect 25450 35646 25452 35698
rect 25396 35644 25452 35646
rect 24612 35420 24668 35476
rect 25564 35532 25620 35588
rect 24220 35308 24276 35364
rect 24444 34076 24500 34132
rect 24108 33292 24164 33348
rect 24780 33628 24836 33684
rect 26516 35420 26572 35476
rect 25564 34636 25620 34692
rect 25004 33628 25060 33684
rect 26460 34524 26516 34580
rect 26572 34300 26628 34356
rect 26516 34130 26572 34132
rect 26516 34078 26518 34130
rect 26518 34078 26570 34130
rect 26570 34078 26572 34130
rect 26516 34076 26572 34078
rect 25788 33292 25844 33348
rect 24556 32732 24612 32788
rect 26460 33346 26516 33348
rect 26460 33294 26462 33346
rect 26462 33294 26514 33346
rect 26514 33294 26516 33346
rect 26460 33292 26516 33294
rect 25116 33068 25172 33124
rect 24444 32060 24500 32116
rect 23884 31724 23940 31780
rect 20972 29314 21028 29316
rect 20972 29262 20974 29314
rect 20974 29262 21026 29314
rect 21026 29262 21028 29314
rect 20972 29260 21028 29262
rect 21308 28924 21364 28980
rect 21420 29372 21476 29428
rect 21420 28700 21476 28756
rect 21532 28812 21588 28868
rect 20524 27916 20580 27972
rect 19964 27858 20020 27860
rect 19964 27806 19966 27858
rect 19966 27806 20018 27858
rect 20018 27806 20020 27858
rect 19964 27804 20020 27806
rect 21868 29932 21924 29988
rect 21868 29036 21924 29092
rect 22540 29372 22596 29428
rect 22876 29426 22932 29428
rect 22876 29374 22878 29426
rect 22878 29374 22930 29426
rect 22930 29374 22932 29426
rect 22876 29372 22932 29374
rect 23268 30492 23324 30548
rect 23548 29596 23604 29652
rect 24444 31612 24500 31668
rect 25340 32786 25396 32788
rect 25340 32734 25342 32786
rect 25342 32734 25394 32786
rect 25394 32734 25396 32786
rect 25340 32732 25396 32734
rect 25452 31750 25508 31780
rect 25452 31724 25454 31750
rect 25454 31724 25506 31750
rect 25506 31724 25508 31750
rect 25676 31836 25732 31892
rect 25564 31612 25620 31668
rect 24780 31164 24836 31220
rect 24556 30994 24612 30996
rect 24556 30942 24558 30994
rect 24558 30942 24610 30994
rect 24610 30942 24612 30994
rect 24556 30940 24612 30942
rect 24668 30828 24724 30884
rect 24444 29650 24500 29652
rect 24444 29598 24446 29650
rect 24446 29598 24498 29650
rect 24498 29598 24500 29650
rect 24444 29596 24500 29598
rect 23100 29260 23156 29316
rect 22316 29036 22372 29092
rect 22428 28642 22484 28644
rect 22428 28590 22430 28642
rect 22430 28590 22482 28642
rect 22482 28590 22484 28642
rect 22428 28588 22484 28590
rect 19516 27356 19572 27412
rect 20860 27833 20862 27860
rect 20862 27833 20914 27860
rect 20914 27833 20916 27860
rect 20860 27804 20916 27833
rect 21644 27839 21646 27860
rect 21646 27839 21698 27860
rect 21698 27839 21700 27860
rect 21644 27804 21700 27839
rect 19180 26796 19236 26852
rect 18284 26066 18340 26068
rect 18284 26014 18286 26066
rect 18286 26014 18338 26066
rect 18338 26014 18340 26066
rect 18284 26012 18340 26014
rect 17500 24444 17556 24500
rect 17612 25116 17668 25172
rect 17724 24220 17780 24276
rect 17612 23996 17668 24052
rect 17388 23826 17444 23828
rect 17388 23774 17390 23826
rect 17390 23774 17442 23826
rect 17442 23774 17444 23826
rect 17388 23772 17444 23774
rect 17556 23772 17612 23828
rect 17612 23212 17668 23268
rect 17052 21420 17108 21476
rect 17948 23938 18004 23940
rect 17948 23886 17950 23938
rect 17950 23886 18002 23938
rect 18002 23886 18004 23938
rect 17948 23884 18004 23886
rect 17724 22988 17780 23044
rect 16940 19964 16996 20020
rect 17276 21868 17332 21924
rect 17500 21644 17556 21700
rect 17612 21756 17668 21812
rect 17444 20860 17500 20916
rect 17948 20300 18004 20356
rect 18564 24498 18620 24500
rect 18564 24446 18566 24498
rect 18566 24446 18618 24498
rect 18618 24446 18620 24498
rect 18564 24444 18620 24446
rect 18284 24108 18340 24164
rect 18844 24444 18900 24500
rect 18284 23772 18340 23828
rect 18340 23212 18396 23268
rect 18060 20748 18116 20804
rect 17612 20076 17668 20132
rect 18172 22988 18228 23044
rect 17612 19906 17668 19908
rect 17612 19854 17614 19906
rect 17614 19854 17666 19906
rect 17666 19854 17668 19906
rect 17612 19852 17668 19854
rect 13916 18844 13972 18900
rect 13916 18508 13972 18564
rect 16716 19628 16772 19684
rect 14588 19346 14644 19348
rect 14588 19294 14590 19346
rect 14590 19294 14642 19346
rect 14642 19294 14644 19346
rect 14588 19292 14644 19294
rect 15092 19234 15148 19236
rect 15092 19182 15094 19234
rect 15094 19182 15146 19234
rect 15146 19182 15148 19234
rect 15092 19180 15148 19182
rect 15596 18956 15652 19012
rect 15820 18620 15876 18676
rect 15036 18396 15092 18452
rect 13580 17948 13636 18004
rect 12796 17052 12852 17108
rect 13860 17666 13916 17668
rect 13860 17614 13862 17666
rect 13862 17614 13914 17666
rect 13914 17614 13916 17666
rect 13860 17612 13916 17614
rect 13468 16044 13524 16100
rect 13692 16828 13748 16884
rect 14812 17724 14868 17780
rect 15540 18060 15596 18116
rect 15932 18060 15988 18116
rect 16436 19292 16492 19348
rect 16268 19234 16324 19236
rect 16268 19182 16270 19234
rect 16270 19182 16322 19234
rect 16322 19182 16324 19234
rect 16268 19180 16324 19182
rect 21532 26796 21588 26852
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19180 25564 19236 25620
rect 19628 25618 19684 25620
rect 19628 25566 19630 25618
rect 19630 25566 19682 25618
rect 19682 25566 19684 25618
rect 19628 25564 19684 25566
rect 19852 25676 19908 25732
rect 20188 25900 20244 25956
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 18956 23884 19012 23940
rect 18732 23548 18788 23604
rect 18788 23378 18844 23380
rect 18788 23326 18790 23378
rect 18790 23326 18842 23378
rect 18842 23326 18844 23378
rect 18788 23324 18844 23326
rect 18620 21308 18676 21364
rect 18508 21196 18564 21252
rect 19292 23548 19348 23604
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 22428 27842 22430 27860
rect 22430 27842 22482 27860
rect 22482 27842 22484 27860
rect 22428 27804 22484 27842
rect 23380 29202 23436 29204
rect 23380 29150 23382 29202
rect 23382 29150 23434 29202
rect 23434 29150 23436 29202
rect 23380 29148 23436 29150
rect 21980 27468 22036 27524
rect 20300 25730 20356 25732
rect 20300 25678 20302 25730
rect 20302 25678 20354 25730
rect 20354 25678 20356 25730
rect 20300 25676 20356 25678
rect 22316 26684 22372 26740
rect 22744 27468 22800 27524
rect 22764 26348 22820 26404
rect 22764 25564 22820 25620
rect 20412 24668 20468 24724
rect 20412 23884 20468 23940
rect 19908 23154 19964 23156
rect 19908 23102 19910 23154
rect 19910 23102 19962 23154
rect 19962 23102 19964 23154
rect 19908 23100 19964 23102
rect 18844 21756 18900 21812
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 21756 24722 21812 24724
rect 21756 24670 21758 24722
rect 21758 24670 21810 24722
rect 21810 24670 21812 24722
rect 21756 24668 21812 24670
rect 23324 28924 23380 28980
rect 23436 27858 23492 27860
rect 23436 27806 23438 27858
rect 23438 27806 23490 27858
rect 23490 27806 23492 27858
rect 23436 27804 23492 27806
rect 23100 27132 23156 27188
rect 23436 25618 23492 25620
rect 23436 25566 23438 25618
rect 23438 25566 23490 25618
rect 23490 25566 23492 25618
rect 23436 25564 23492 25566
rect 23100 24892 23156 24948
rect 23884 24892 23940 24948
rect 23772 24556 23828 24612
rect 22671 23996 22727 24052
rect 21420 23714 21476 23716
rect 21420 23662 21422 23714
rect 21422 23662 21474 23714
rect 21474 23662 21476 23714
rect 21420 23660 21476 23662
rect 21084 23324 21140 23380
rect 20916 23212 20972 23268
rect 20636 22988 20692 23044
rect 21084 22988 21140 23044
rect 22428 23938 22484 23940
rect 22428 23886 22430 23938
rect 22430 23886 22482 23938
rect 22482 23886 22484 23938
rect 22428 23884 22484 23886
rect 20860 22370 20916 22372
rect 20860 22318 20862 22370
rect 20862 22318 20914 22370
rect 20914 22318 20916 22370
rect 20860 22316 20916 22318
rect 20524 22146 20580 22148
rect 20524 22094 20526 22146
rect 20526 22094 20578 22146
rect 20578 22094 20580 22146
rect 20524 22092 20580 22094
rect 19272 20972 19328 21028
rect 18396 20300 18452 20356
rect 18508 20748 18564 20804
rect 20188 21196 20244 21252
rect 20356 21196 20412 21252
rect 20188 20972 20244 21028
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 21644 22316 21700 22372
rect 21868 21980 21924 22036
rect 22484 22652 22540 22708
rect 22484 21756 22540 21812
rect 24444 29036 24500 29092
rect 24220 28588 24276 28644
rect 24220 27186 24276 27188
rect 24220 27134 24222 27186
rect 24222 27134 24274 27186
rect 24274 27134 24276 27186
rect 24220 27132 24276 27134
rect 24276 26178 24332 26180
rect 24276 26126 24278 26178
rect 24278 26126 24330 26178
rect 24330 26126 24332 26178
rect 24276 26124 24332 26126
rect 24780 30716 24836 30772
rect 25284 30770 25340 30772
rect 25284 30718 25286 30770
rect 25286 30718 25338 30770
rect 25338 30718 25340 30770
rect 25284 30716 25340 30718
rect 25340 29426 25396 29428
rect 25340 29374 25342 29426
rect 25342 29374 25394 29426
rect 25394 29374 25396 29426
rect 25340 29372 25396 29374
rect 26888 36988 26944 37044
rect 27748 36988 27804 37044
rect 28924 43148 28980 43204
rect 30044 45890 30100 45892
rect 30044 45838 30046 45890
rect 30046 45838 30098 45890
rect 30098 45838 30100 45890
rect 30044 45836 30100 45838
rect 30380 46674 30436 46676
rect 30380 46622 30382 46674
rect 30382 46622 30434 46674
rect 30434 46622 30436 46674
rect 30380 46620 30436 46622
rect 31164 46956 31220 47012
rect 30268 45836 30324 45892
rect 30884 46450 30940 46452
rect 30884 46398 30886 46450
rect 30886 46398 30938 46450
rect 30938 46398 30940 46450
rect 30884 46396 30940 46398
rect 30828 46002 30884 46004
rect 30828 45950 30830 46002
rect 30830 45950 30882 46002
rect 30882 45950 30884 46002
rect 30828 45948 30884 45950
rect 31500 46396 31556 46452
rect 39284 48076 39340 48132
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 38836 47628 38892 47684
rect 32620 47570 32676 47572
rect 32620 47518 32622 47570
rect 32622 47518 32674 47570
rect 32674 47518 32676 47570
rect 32620 47516 32676 47518
rect 33852 47516 33908 47572
rect 32172 47180 32228 47236
rect 32508 47068 32564 47124
rect 32956 46674 33012 46676
rect 32956 46622 32958 46674
rect 32958 46622 33010 46674
rect 33010 46622 33012 46674
rect 32956 46620 33012 46622
rect 31724 45612 31780 45668
rect 30604 45106 30660 45108
rect 30604 45054 30606 45106
rect 30606 45054 30658 45106
rect 30658 45054 30660 45106
rect 30604 45052 30660 45054
rect 31052 45093 31054 45108
rect 31054 45093 31106 45108
rect 31106 45093 31108 45108
rect 31052 45052 31108 45093
rect 29260 44716 29316 44772
rect 29372 44604 29428 44660
rect 32060 45612 32116 45668
rect 32228 45106 32284 45108
rect 32228 45054 32230 45106
rect 32230 45054 32282 45106
rect 32282 45054 32284 45106
rect 32228 45052 32284 45054
rect 29540 44322 29596 44324
rect 29540 44270 29542 44322
rect 29542 44270 29594 44322
rect 29594 44270 29596 44322
rect 29540 44268 29596 44270
rect 29148 43932 29204 43988
rect 29148 43372 29204 43428
rect 29372 43484 29428 43540
rect 29260 42754 29316 42756
rect 29260 42702 29262 42754
rect 29262 42702 29314 42754
rect 29314 42702 29316 42754
rect 29260 42700 29316 42702
rect 29148 42252 29204 42308
rect 28980 41858 29036 41860
rect 28980 41806 28982 41858
rect 28982 41806 29034 41858
rect 29034 41806 29036 41858
rect 28980 41804 29036 41806
rect 29036 41186 29092 41188
rect 29036 41134 29038 41186
rect 29038 41134 29090 41186
rect 29090 41134 29092 41186
rect 29036 41132 29092 41134
rect 28980 40572 29036 40628
rect 28812 39004 28868 39060
rect 28364 38556 28420 38612
rect 28476 38332 28532 38388
rect 28588 38108 28644 38164
rect 28924 38220 28980 38276
rect 28028 36454 28084 36484
rect 28028 36428 28030 36454
rect 28030 36428 28082 36454
rect 28082 36428 28084 36454
rect 27356 36316 27412 36372
rect 27524 35980 27580 36036
rect 28028 36204 28084 36260
rect 27132 35674 27134 35700
rect 27134 35674 27186 35700
rect 27186 35674 27188 35700
rect 27692 35756 27748 35812
rect 27132 35644 27188 35674
rect 27580 35420 27636 35476
rect 27020 34636 27076 34692
rect 26852 33234 26908 33236
rect 26852 33182 26854 33234
rect 26854 33182 26906 33234
rect 26906 33182 26908 33234
rect 26852 33180 26908 33182
rect 27244 34354 27300 34356
rect 27244 34302 27246 34354
rect 27246 34302 27298 34354
rect 27298 34302 27300 34354
rect 27244 34300 27300 34302
rect 27692 34188 27748 34244
rect 26012 31948 26068 32004
rect 25788 31164 25844 31220
rect 26124 31276 26180 31332
rect 25788 30970 25790 30996
rect 25790 30970 25842 30996
rect 25842 30970 25844 30996
rect 25788 30940 25844 30970
rect 25676 29372 25732 29428
rect 26012 30210 26068 30212
rect 26012 30158 26014 30210
rect 26014 30158 26066 30210
rect 26066 30158 26068 30210
rect 26012 30156 26068 30158
rect 26124 29596 26180 29652
rect 25732 28754 25788 28756
rect 25732 28702 25734 28754
rect 25734 28702 25786 28754
rect 25786 28702 25788 28754
rect 25732 28700 25788 28702
rect 25396 27746 25452 27748
rect 25396 27694 25398 27746
rect 25398 27694 25450 27746
rect 25450 27694 25452 27746
rect 25396 27692 25452 27694
rect 25676 27692 25732 27748
rect 25452 26796 25508 26852
rect 25340 26572 25396 26628
rect 24724 26290 24780 26292
rect 24724 26238 24726 26290
rect 24726 26238 24778 26290
rect 24778 26238 24780 26290
rect 24724 26236 24780 26238
rect 25228 26273 25230 26292
rect 25230 26273 25282 26292
rect 25282 26273 25284 26292
rect 25228 26236 25284 26273
rect 24220 24780 24276 24836
rect 24444 24610 24500 24612
rect 24444 24558 24446 24610
rect 24446 24558 24498 24610
rect 24498 24558 24500 24610
rect 24444 24556 24500 24558
rect 24220 23938 24276 23940
rect 24220 23886 24222 23938
rect 24222 23886 24274 23938
rect 24274 23886 24276 23938
rect 24220 23884 24276 23886
rect 24444 23938 24500 23940
rect 24444 23886 24446 23938
rect 24446 23886 24498 23938
rect 24498 23886 24500 23938
rect 24444 23884 24500 23886
rect 23212 21868 23268 21924
rect 22652 21756 22708 21812
rect 21756 21532 21812 21588
rect 22428 21196 22484 21252
rect 22092 21084 22148 21140
rect 22652 21196 22708 21252
rect 22876 21586 22932 21588
rect 22876 21534 22878 21586
rect 22878 21534 22930 21586
rect 22930 21534 22932 21586
rect 22876 21532 22932 21534
rect 22204 20636 22260 20692
rect 16604 19122 16660 19124
rect 16604 19070 16606 19122
rect 16606 19070 16658 19122
rect 16658 19070 16660 19122
rect 16604 19068 16660 19070
rect 18732 19852 18788 19908
rect 16156 17836 16212 17892
rect 16492 18844 16548 18900
rect 15820 17778 15876 17780
rect 15820 17726 15822 17778
rect 15822 17726 15874 17778
rect 15874 17726 15876 17778
rect 15820 17724 15876 17726
rect 14812 17500 14868 17556
rect 17500 18508 17556 18564
rect 16716 18060 16772 18116
rect 17276 18060 17332 18116
rect 19852 20076 19908 20132
rect 18956 19852 19012 19908
rect 19628 19794 19684 19796
rect 19628 19742 19630 19794
rect 19630 19742 19682 19794
rect 19682 19742 19684 19794
rect 19628 19740 19684 19742
rect 20412 19964 20468 20020
rect 20188 19852 20244 19908
rect 20076 19740 20132 19796
rect 18396 18284 18452 18340
rect 18060 17836 18116 17892
rect 18396 17836 18452 17892
rect 16716 17666 16772 17668
rect 16716 17614 16718 17666
rect 16718 17614 16770 17666
rect 16770 17614 16772 17666
rect 16716 17612 16772 17614
rect 17948 17666 18004 17668
rect 17948 17614 17950 17666
rect 17950 17614 18002 17666
rect 18002 17614 18004 17666
rect 17948 17612 18004 17614
rect 18956 18426 18958 18452
rect 18958 18426 19010 18452
rect 19010 18426 19012 18452
rect 18956 18396 19012 18426
rect 19348 17836 19404 17892
rect 18844 17612 18900 17668
rect 16996 17554 17052 17556
rect 16996 17502 16998 17554
rect 16998 17502 17050 17554
rect 17050 17502 17052 17554
rect 16996 17500 17052 17502
rect 16156 17388 16212 17444
rect 16604 17388 16660 17444
rect 14028 16828 14084 16884
rect 15036 16940 15092 16996
rect 13636 15874 13692 15876
rect 13636 15822 13638 15874
rect 13638 15822 13690 15874
rect 13690 15822 13692 15874
rect 13636 15820 13692 15822
rect 9996 15036 10052 15092
rect 11228 15036 11284 15092
rect 10444 14642 10500 14644
rect 10444 14590 10446 14642
rect 10446 14590 10498 14642
rect 10498 14590 10500 14642
rect 10444 14588 10500 14590
rect 9996 14476 10052 14532
rect 10220 14476 10276 14532
rect 13916 16098 13972 16100
rect 13916 16046 13918 16098
rect 13918 16046 13970 16098
rect 13970 16046 13972 16098
rect 13916 16044 13972 16046
rect 16380 16940 16436 16996
rect 16044 16882 16100 16884
rect 16044 16830 16046 16882
rect 16046 16830 16098 16882
rect 16098 16830 16100 16882
rect 17612 17442 17668 17444
rect 17612 17390 17614 17442
rect 17614 17390 17666 17442
rect 17666 17390 17668 17442
rect 17612 17388 17668 17390
rect 16044 16828 16100 16830
rect 16660 16604 16716 16660
rect 15932 15820 15988 15876
rect 14588 15202 14644 15204
rect 14588 15150 14590 15202
rect 14590 15150 14642 15202
rect 14642 15150 14644 15202
rect 14588 15148 14644 15150
rect 11900 15036 11956 15092
rect 13468 15036 13524 15092
rect 12124 14588 12180 14644
rect 10220 13468 10276 13524
rect 9884 13244 9940 13300
rect 10220 12236 10276 12292
rect 10444 12178 10500 12180
rect 10444 12126 10446 12178
rect 10446 12126 10498 12178
rect 10498 12126 10500 12178
rect 10444 12124 10500 12126
rect 13132 14588 13188 14644
rect 12460 14530 12516 14532
rect 12460 14478 12462 14530
rect 12462 14478 12514 14530
rect 12514 14478 12516 14530
rect 12460 14476 12516 14478
rect 13020 14476 13076 14532
rect 11004 12012 11060 12068
rect 9716 11900 9772 11956
rect 9548 11788 9604 11844
rect 9212 11228 9268 11284
rect 8876 11116 8932 11172
rect 10444 11228 10500 11284
rect 9324 10780 9380 10836
rect 9660 10556 9716 10612
rect 11228 11116 11284 11172
rect 11676 12124 11732 12180
rect 11564 11116 11620 11172
rect 11900 11564 11956 11620
rect 11228 10722 11284 10724
rect 11228 10670 11230 10722
rect 11230 10670 11282 10722
rect 11282 10670 11284 10722
rect 11228 10668 11284 10670
rect 12460 12348 12516 12404
rect 13804 14476 13860 14532
rect 14252 13020 14308 13076
rect 13188 12348 13244 12404
rect 11900 11394 11956 11396
rect 11900 11342 11902 11394
rect 11902 11342 11954 11394
rect 11954 11342 11956 11394
rect 11900 11340 11956 11342
rect 12348 11452 12404 11508
rect 13188 11340 13244 11396
rect 11788 10668 11844 10724
rect 11900 11116 11956 11172
rect 10108 9884 10164 9940
rect 10780 9826 10836 9828
rect 10780 9774 10782 9826
rect 10782 9774 10834 9826
rect 10834 9774 10836 9826
rect 10780 9772 10836 9774
rect 8652 8818 8708 8820
rect 8652 8766 8654 8818
rect 8654 8766 8706 8818
rect 8706 8766 8708 8818
rect 8652 8764 8708 8766
rect 10444 8764 10500 8820
rect 8652 7586 8708 7588
rect 8652 7534 8654 7586
rect 8654 7534 8706 7586
rect 8706 7534 8708 7586
rect 8652 7532 8708 7534
rect 7980 6300 8036 6356
rect 8428 6636 8484 6692
rect 7140 5740 7196 5796
rect 7308 5740 7364 5796
rect 7532 5740 7588 5796
rect 7700 5682 7756 5684
rect 7700 5630 7702 5682
rect 7702 5630 7754 5682
rect 7754 5630 7756 5682
rect 7700 5628 7756 5630
rect 8092 5906 8148 5908
rect 8092 5854 8094 5906
rect 8094 5854 8146 5906
rect 8146 5854 8148 5906
rect 8428 6300 8484 6356
rect 8540 6076 8596 6132
rect 8428 6018 8484 6020
rect 8428 5966 8430 6018
rect 8430 5966 8482 6018
rect 8482 5966 8484 6018
rect 8428 5964 8484 5966
rect 10108 8146 10164 8148
rect 10108 8094 10110 8146
rect 10110 8094 10162 8146
rect 10162 8094 10164 8146
rect 10108 8092 10164 8094
rect 9884 7644 9940 7700
rect 9660 7474 9716 7476
rect 9660 7422 9662 7474
rect 9662 7422 9714 7474
rect 9714 7422 9716 7474
rect 9660 7420 9716 7422
rect 9772 6802 9828 6804
rect 9772 6750 9774 6802
rect 9774 6750 9826 6802
rect 9826 6750 9828 6802
rect 9772 6748 9828 6750
rect 9548 6300 9604 6356
rect 9436 6076 9492 6132
rect 8988 5964 9044 6020
rect 8092 5852 8148 5854
rect 7868 5292 7924 5348
rect 8428 5628 8484 5684
rect 7980 5234 8036 5236
rect 7980 5182 7982 5234
rect 7982 5182 8034 5234
rect 8034 5182 8036 5234
rect 7980 5180 8036 5182
rect 7868 5107 7924 5124
rect 7868 5068 7870 5107
rect 7870 5068 7922 5107
rect 7922 5068 7924 5107
rect 6972 4338 7028 4340
rect 6972 4286 6974 4338
rect 6974 4286 7026 4338
rect 7026 4286 7028 4338
rect 6972 4284 7028 4286
rect 9436 5852 9492 5908
rect 8876 5292 8932 5348
rect 8540 5068 8596 5124
rect 8652 5180 8708 5236
rect 9212 5292 9268 5348
rect 9772 5852 9828 5908
rect 10444 7532 10500 7588
rect 10108 7362 10164 7364
rect 10108 7310 10110 7362
rect 10110 7310 10162 7362
rect 10162 7310 10164 7362
rect 10108 7308 10164 7310
rect 10668 8204 10724 8260
rect 10892 8092 10948 8148
rect 11228 7644 11284 7700
rect 10556 6860 10612 6916
rect 10780 6748 10836 6804
rect 9996 6300 10052 6356
rect 10220 5964 10276 6020
rect 9996 5292 10052 5348
rect 10332 5906 10388 5908
rect 10332 5854 10334 5906
rect 10334 5854 10386 5906
rect 10386 5854 10388 5906
rect 10332 5852 10388 5854
rect 12572 11228 12628 11284
rect 13524 11282 13580 11284
rect 13524 11230 13526 11282
rect 13526 11230 13578 11282
rect 13578 11230 13580 11282
rect 13524 11228 13580 11230
rect 12572 10780 12628 10836
rect 12236 10220 12292 10276
rect 12348 9938 12404 9940
rect 12348 9886 12350 9938
rect 12350 9886 12402 9938
rect 12402 9886 12404 9938
rect 12348 9884 12404 9886
rect 11564 8988 11620 9044
rect 12796 9042 12852 9044
rect 12796 8990 12798 9042
rect 12798 8990 12850 9042
rect 12850 8990 12852 9042
rect 12796 8988 12852 8990
rect 14476 12236 14532 12292
rect 14812 12066 14868 12068
rect 14812 12014 14814 12066
rect 14814 12014 14866 12066
rect 14866 12014 14868 12066
rect 14812 12012 14868 12014
rect 13916 11564 13972 11620
rect 13804 11394 13860 11396
rect 13804 11342 13806 11394
rect 13806 11342 13858 11394
rect 13858 11342 13860 11394
rect 13804 11340 13860 11342
rect 14588 11564 14644 11620
rect 14252 11506 14308 11508
rect 14252 11454 14254 11506
rect 14254 11454 14306 11506
rect 14306 11454 14308 11506
rect 14252 11452 14308 11454
rect 14364 11379 14420 11396
rect 14364 11340 14366 11379
rect 14366 11340 14418 11379
rect 14418 11340 14420 11379
rect 17164 16098 17220 16100
rect 17164 16046 17166 16098
rect 17166 16046 17218 16098
rect 17218 16046 17220 16098
rect 17164 16044 17220 16046
rect 17948 16828 18004 16884
rect 18172 16604 18228 16660
rect 18396 16380 18452 16436
rect 18844 16604 18900 16660
rect 16492 14476 16548 14532
rect 17276 14530 17332 14532
rect 16156 14418 16212 14420
rect 16156 14366 16158 14418
rect 16158 14366 16210 14418
rect 16210 14366 16212 14418
rect 16156 14364 16212 14366
rect 16716 14364 16772 14420
rect 16324 13522 16380 13524
rect 16324 13470 16326 13522
rect 16326 13470 16378 13522
rect 16378 13470 16380 13522
rect 16324 13468 16380 13470
rect 17276 14478 17278 14530
rect 17278 14478 17330 14530
rect 17330 14478 17332 14530
rect 17276 14476 17332 14478
rect 17500 14476 17556 14532
rect 16940 14364 16996 14420
rect 17612 13916 17668 13972
rect 16828 13804 16884 13860
rect 18060 15202 18116 15204
rect 18060 15150 18062 15202
rect 18062 15150 18114 15202
rect 18114 15150 18116 15202
rect 18060 15148 18116 15150
rect 18620 15148 18676 15204
rect 18396 14530 18452 14532
rect 18396 14478 18398 14530
rect 18398 14478 18450 14530
rect 18450 14478 18452 14530
rect 18396 14476 18452 14478
rect 19516 16828 19572 16884
rect 19068 16380 19124 16436
rect 19516 16156 19572 16212
rect 19218 15300 19220 15316
rect 19220 15300 19272 15316
rect 19272 15300 19274 15316
rect 19218 15260 19274 15300
rect 18956 14588 19012 14644
rect 18116 14418 18172 14420
rect 18116 14366 18118 14418
rect 18118 14366 18170 14418
rect 18170 14366 18172 14418
rect 18116 14364 18172 14366
rect 17836 13804 17892 13860
rect 17948 13746 18004 13748
rect 17948 13694 17950 13746
rect 17950 13694 18002 13746
rect 18002 13694 18004 13746
rect 17948 13692 18004 13694
rect 17836 13468 17892 13524
rect 19292 15036 19348 15092
rect 19068 14502 19124 14532
rect 19068 14476 19070 14502
rect 19070 14476 19122 14502
rect 19122 14476 19124 14502
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 22428 20300 22484 20356
rect 21028 20018 21084 20020
rect 21028 19966 21030 20018
rect 21030 19966 21082 20018
rect 21082 19966 21084 20018
rect 21028 19964 21084 19966
rect 21868 20018 21924 20020
rect 21868 19966 21870 20018
rect 21870 19966 21922 20018
rect 21922 19966 21924 20018
rect 21868 19964 21924 19966
rect 21476 19906 21532 19908
rect 21476 19854 21478 19906
rect 21478 19854 21530 19906
rect 21530 19854 21532 19906
rect 21476 19852 21532 19854
rect 20860 19234 20916 19236
rect 20860 19182 20862 19234
rect 20862 19182 20914 19234
rect 20914 19182 20916 19234
rect 20860 19180 20916 19182
rect 21196 19234 21252 19236
rect 21196 19182 21198 19234
rect 21198 19182 21250 19234
rect 21250 19182 21252 19234
rect 21196 19180 21252 19182
rect 20524 18508 20580 18564
rect 20916 18732 20972 18788
rect 20748 18450 20804 18452
rect 20748 18398 20750 18450
rect 20750 18398 20802 18450
rect 20802 18398 20804 18450
rect 20748 18396 20804 18398
rect 23100 21420 23156 21476
rect 23100 20860 23156 20916
rect 23436 20748 23492 20804
rect 22540 19852 22596 19908
rect 22876 19964 22932 20020
rect 23212 19068 23268 19124
rect 21980 18732 22036 18788
rect 21868 18396 21924 18452
rect 22272 18508 22328 18564
rect 21532 18284 21588 18340
rect 22540 18284 22596 18340
rect 21420 17724 21476 17780
rect 20860 17500 20916 17556
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20132 16156 20188 16212
rect 19964 16077 20020 16100
rect 19964 16044 19966 16077
rect 19966 16044 20018 16077
rect 20018 16044 20020 16077
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20020 15538 20076 15540
rect 20020 15486 20022 15538
rect 20022 15486 20074 15538
rect 20074 15486 20076 15538
rect 20020 15484 20076 15486
rect 19516 15148 19572 15204
rect 19404 14588 19460 14644
rect 19068 13970 19124 13972
rect 19068 13918 19070 13970
rect 19070 13918 19122 13970
rect 19122 13918 19124 13970
rect 19068 13916 19124 13918
rect 20300 15484 20356 15540
rect 20524 15260 20580 15316
rect 20636 14588 20692 14644
rect 20188 14252 20244 14308
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19516 13804 19572 13860
rect 18956 13692 19012 13748
rect 18116 13356 18172 13412
rect 18060 13074 18116 13076
rect 18060 13022 18062 13074
rect 18062 13022 18114 13074
rect 18114 13022 18116 13074
rect 18060 13020 18116 13022
rect 18620 13468 18676 13524
rect 19740 13746 19796 13748
rect 19740 13694 19742 13746
rect 19742 13694 19794 13746
rect 19794 13694 19796 13746
rect 19740 13692 19796 13694
rect 20188 13692 20244 13748
rect 20524 13804 20580 13860
rect 20300 13580 20356 13636
rect 19404 13468 19460 13524
rect 19628 13468 19684 13524
rect 18788 13356 18844 13412
rect 18620 12962 18676 12964
rect 18620 12910 18622 12962
rect 18622 12910 18674 12962
rect 18674 12910 18676 12962
rect 18620 12908 18676 12910
rect 18060 12290 18116 12292
rect 18060 12238 18062 12290
rect 18062 12238 18114 12290
rect 18114 12238 18116 12290
rect 18060 12236 18116 12238
rect 18228 12236 18284 12292
rect 17836 12178 17892 12180
rect 17836 12126 17838 12178
rect 17838 12126 17890 12178
rect 17890 12126 17892 12178
rect 18508 12178 18564 12180
rect 17836 12124 17892 12126
rect 14812 10498 14868 10500
rect 14812 10446 14814 10498
rect 14814 10446 14866 10498
rect 14866 10446 14868 10498
rect 14812 10444 14868 10446
rect 16324 11506 16380 11508
rect 16324 11454 16326 11506
rect 16326 11454 16378 11506
rect 16378 11454 16380 11506
rect 16324 11452 16380 11454
rect 16940 11452 16996 11508
rect 18508 12126 18510 12178
rect 18510 12126 18562 12178
rect 18562 12126 18564 12178
rect 18508 12124 18564 12126
rect 19068 12908 19124 12964
rect 18116 11788 18172 11844
rect 18284 11564 18340 11620
rect 16660 11170 16716 11172
rect 16660 11118 16662 11170
rect 16662 11118 16714 11170
rect 16714 11118 16716 11170
rect 16660 11116 16716 11118
rect 17612 11116 17668 11172
rect 17276 10780 17332 10836
rect 17556 10668 17612 10724
rect 14812 9660 14868 9716
rect 17724 10498 17780 10500
rect 17724 10446 17726 10498
rect 17726 10446 17778 10498
rect 17778 10446 17780 10498
rect 17724 10444 17780 10446
rect 16716 9772 16772 9828
rect 17724 9826 17780 9828
rect 17724 9774 17726 9826
rect 17726 9774 17778 9826
rect 17778 9774 17780 9826
rect 17724 9772 17780 9774
rect 15148 9212 15204 9268
rect 17052 9548 17108 9604
rect 12348 8258 12404 8260
rect 12348 8206 12350 8258
rect 12350 8206 12402 8258
rect 12402 8206 12404 8258
rect 12348 8204 12404 8206
rect 11844 7586 11900 7588
rect 11844 7534 11846 7586
rect 11846 7534 11898 7586
rect 11898 7534 11900 7586
rect 11844 7532 11900 7534
rect 12292 7586 12348 7588
rect 12292 7534 12294 7586
rect 12294 7534 12346 7586
rect 12346 7534 12348 7586
rect 12292 7532 12348 7534
rect 13448 7532 13504 7588
rect 11116 7308 11172 7364
rect 12236 6802 12292 6804
rect 12236 6750 12238 6802
rect 12238 6750 12290 6802
rect 12290 6750 12292 6802
rect 12236 6748 12292 6750
rect 13692 6748 13748 6804
rect 11452 6412 11508 6468
rect 14812 8540 14868 8596
rect 17948 10610 18004 10612
rect 17948 10558 17950 10610
rect 17950 10558 18002 10610
rect 18002 10558 18004 10610
rect 17948 10556 18004 10558
rect 19964 12962 20020 12964
rect 19964 12910 19966 12962
rect 19966 12910 20018 12962
rect 20018 12910 20020 12962
rect 19964 12908 20020 12910
rect 20860 15484 20916 15540
rect 21980 17554 22036 17556
rect 21980 17502 21982 17554
rect 21982 17502 22034 17554
rect 22034 17502 22036 17554
rect 21980 17500 22036 17502
rect 21756 17052 21812 17108
rect 22092 16828 22148 16884
rect 22204 16098 22260 16100
rect 22204 16046 22206 16098
rect 22206 16046 22258 16098
rect 22258 16046 22260 16098
rect 22204 16044 22260 16046
rect 21980 15260 22036 15316
rect 22428 15484 22484 15540
rect 22428 15260 22484 15316
rect 21084 14476 21140 14532
rect 21644 14252 21700 14308
rect 21084 14028 21140 14084
rect 22540 14252 22596 14308
rect 21756 13692 21812 13748
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19180 12236 19236 12292
rect 19740 12066 19796 12068
rect 19740 12014 19742 12066
rect 19742 12014 19794 12066
rect 19794 12014 19796 12066
rect 19740 12012 19796 12014
rect 19014 11394 19070 11396
rect 19014 11342 19016 11394
rect 19016 11342 19068 11394
rect 19068 11342 19070 11394
rect 19014 11340 19070 11342
rect 18620 10668 18676 10724
rect 19292 11676 19348 11732
rect 18060 10444 18116 10500
rect 18060 9548 18116 9604
rect 16716 8930 16772 8932
rect 16716 8878 16718 8930
rect 16718 8878 16770 8930
rect 16770 8878 16772 8930
rect 16716 8876 16772 8878
rect 16156 8230 16212 8260
rect 16156 8204 16158 8230
rect 16158 8204 16210 8230
rect 16210 8204 16212 8230
rect 16044 8092 16100 8148
rect 14140 6802 14196 6804
rect 14140 6750 14142 6802
rect 14142 6750 14194 6802
rect 14194 6750 14196 6802
rect 14140 6748 14196 6750
rect 16044 6412 16100 6468
rect 16716 6636 16772 6692
rect 16604 6300 16660 6356
rect 17164 6524 17220 6580
rect 18060 8988 18116 9044
rect 18284 10108 18340 10164
rect 18732 10610 18788 10612
rect 18732 10558 18734 10610
rect 18734 10558 18786 10610
rect 18786 10558 18788 10610
rect 18732 10556 18788 10558
rect 19002 10780 19058 10836
rect 19180 10556 19236 10612
rect 18732 9100 18788 9156
rect 18956 10108 19012 10164
rect 22428 13468 22484 13524
rect 23212 18508 23268 18564
rect 24780 23154 24836 23156
rect 24780 23102 24782 23154
rect 24782 23102 24834 23154
rect 24834 23102 24836 23154
rect 24780 23100 24836 23102
rect 23884 22316 23940 22372
rect 23660 21868 23716 21924
rect 23996 21756 24052 21812
rect 24108 21026 24164 21028
rect 24108 20974 24110 21026
rect 24110 20974 24162 21026
rect 24162 20974 24164 21026
rect 24108 20972 24164 20974
rect 23772 20860 23828 20916
rect 23548 20636 23604 20692
rect 26236 28812 26292 28868
rect 26012 28476 26068 28532
rect 26124 28588 26180 28644
rect 26236 28476 26292 28532
rect 26012 26908 26068 26964
rect 25900 26572 25956 26628
rect 25788 26348 25844 26404
rect 26572 32396 26628 32452
rect 26628 31276 26684 31332
rect 26460 30940 26516 30996
rect 26628 30268 26684 30324
rect 26684 30044 26740 30100
rect 27580 31778 27636 31780
rect 27580 31726 27582 31778
rect 27582 31726 27634 31778
rect 27634 31726 27636 31778
rect 27580 31724 27636 31726
rect 27916 32450 27972 32452
rect 27916 32398 27918 32450
rect 27918 32398 27970 32450
rect 27970 32398 27972 32450
rect 27916 32396 27972 32398
rect 27860 32172 27916 32228
rect 28140 35756 28196 35812
rect 28364 36316 28420 36372
rect 28364 35420 28420 35476
rect 29036 37212 29092 37268
rect 28476 35644 28532 35700
rect 27356 30940 27412 30996
rect 27748 30882 27804 30884
rect 27748 30830 27750 30882
rect 27750 30830 27802 30882
rect 27802 30830 27804 30882
rect 27748 30828 27804 30830
rect 28364 31778 28420 31780
rect 28364 31726 28366 31778
rect 28366 31726 28418 31778
rect 28418 31726 28420 31778
rect 28364 31724 28420 31726
rect 28140 30156 28196 30212
rect 27524 29426 27580 29428
rect 27524 29374 27526 29426
rect 27526 29374 27578 29426
rect 27578 29374 27580 29426
rect 27524 29372 27580 29374
rect 26460 29148 26516 29204
rect 26460 28812 26516 28868
rect 26908 28924 26964 28980
rect 26796 28700 26852 28756
rect 26684 28476 26740 28532
rect 26796 28364 26852 28420
rect 26684 28252 26740 28308
rect 25900 25004 25956 25060
rect 25228 23996 25284 24052
rect 25452 24892 25508 24948
rect 25116 21868 25172 21924
rect 24780 21084 24836 21140
rect 24444 20802 24500 20804
rect 24444 20750 24446 20802
rect 24446 20750 24498 20802
rect 24498 20750 24500 20802
rect 24444 20748 24500 20750
rect 25228 23660 25284 23716
rect 26124 25506 26180 25508
rect 26124 25454 26126 25506
rect 26126 25454 26178 25506
rect 26178 25454 26180 25506
rect 26124 25452 26180 25454
rect 26348 25506 26404 25508
rect 26348 25454 26350 25506
rect 26350 25454 26402 25506
rect 26402 25454 26404 25506
rect 26348 25452 26404 25454
rect 26572 25004 26628 25060
rect 27804 29820 27860 29876
rect 27916 29260 27972 29316
rect 27132 28642 27188 28644
rect 27132 28590 27134 28642
rect 27134 28590 27186 28642
rect 27186 28590 27188 28642
rect 27132 28588 27188 28590
rect 27636 28642 27692 28644
rect 27636 28590 27638 28642
rect 27638 28590 27690 28642
rect 27690 28590 27692 28642
rect 27636 28588 27692 28590
rect 28140 28924 28196 28980
rect 28364 29260 28420 29316
rect 28252 28812 28308 28868
rect 28924 35420 28980 35476
rect 28812 34412 28868 34468
rect 28700 33292 28756 33348
rect 29260 41020 29316 41076
rect 29260 40684 29316 40740
rect 29820 43538 29876 43540
rect 29820 43486 29822 43538
rect 29822 43486 29874 43538
rect 29874 43486 29876 43538
rect 29820 43484 29876 43486
rect 29540 43036 29596 43092
rect 30268 44268 30324 44324
rect 30492 44322 30548 44324
rect 30492 44270 30494 44322
rect 30494 44270 30546 44322
rect 30546 44270 30548 44322
rect 30492 44268 30548 44270
rect 32228 44716 32284 44772
rect 32396 44604 32452 44660
rect 32956 45836 33012 45892
rect 32732 45612 32788 45668
rect 33516 45862 33572 45892
rect 33516 45836 33518 45862
rect 33518 45836 33570 45862
rect 33570 45836 33572 45862
rect 33740 45836 33796 45892
rect 35196 47430 35252 47460
rect 35196 47404 35198 47430
rect 35198 47404 35250 47430
rect 35250 47404 35252 47430
rect 33964 47292 34020 47348
rect 35420 47068 35476 47124
rect 49308 48860 49364 48916
rect 44604 48076 44660 48132
rect 47292 48076 47348 48132
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 34860 45724 34916 45780
rect 31724 44294 31780 44324
rect 31724 44268 31726 44294
rect 31726 44268 31778 44294
rect 31778 44268 31780 44294
rect 32844 44604 32900 44660
rect 32732 44322 32788 44324
rect 32732 44270 32734 44322
rect 32734 44270 32786 44322
rect 32786 44270 32788 44322
rect 32732 44268 32788 44270
rect 30548 43426 30604 43428
rect 30548 43374 30550 43426
rect 30550 43374 30602 43426
rect 30602 43374 30604 43426
rect 30548 43372 30604 43374
rect 30716 42812 30772 42868
rect 30940 43596 30996 43652
rect 29820 42588 29876 42644
rect 30716 42588 30772 42644
rect 29540 41298 29596 41300
rect 29540 41246 29542 41298
rect 29542 41246 29594 41298
rect 29594 41246 29596 41298
rect 29540 41244 29596 41246
rect 30268 41946 30270 41972
rect 30270 41946 30322 41972
rect 30322 41946 30324 41972
rect 30268 41916 30324 41946
rect 30828 41916 30884 41972
rect 30716 41692 30772 41748
rect 30156 41244 30212 41300
rect 29372 40348 29428 40404
rect 29820 40572 29876 40628
rect 29932 40796 29988 40852
rect 29708 40402 29764 40404
rect 29708 40350 29710 40402
rect 29710 40350 29762 40402
rect 29762 40350 29764 40402
rect 30044 40460 30100 40516
rect 30324 41074 30380 41076
rect 30324 41022 30326 41074
rect 30326 41022 30378 41074
rect 30378 41022 30380 41074
rect 30324 41020 30380 41022
rect 29708 40348 29764 40350
rect 29876 39618 29932 39620
rect 29876 39566 29878 39618
rect 29878 39566 29930 39618
rect 29930 39566 29932 39618
rect 29876 39564 29932 39566
rect 30044 39618 30100 39620
rect 30044 39566 30046 39618
rect 30046 39566 30098 39618
rect 30098 39566 30100 39618
rect 30044 39564 30100 39566
rect 30268 40572 30324 40628
rect 30492 40124 30548 40180
rect 29932 39058 29988 39060
rect 29932 39006 29934 39058
rect 29934 39006 29986 39058
rect 29986 39006 29988 39058
rect 29932 39004 29988 39006
rect 29260 38892 29316 38948
rect 30604 39564 30660 39620
rect 31500 43596 31556 43652
rect 31836 43708 31892 43764
rect 31052 43036 31108 43092
rect 31164 42924 31220 42980
rect 31388 42812 31444 42868
rect 31052 41970 31108 41972
rect 31052 41918 31054 41970
rect 31054 41918 31106 41970
rect 31106 41918 31108 41970
rect 31052 41916 31108 41918
rect 31052 41580 31108 41636
rect 30828 40796 30884 40852
rect 30940 40572 30996 40628
rect 31052 41020 31108 41076
rect 31836 42924 31892 42980
rect 32172 43538 32228 43540
rect 32172 43486 32174 43538
rect 32174 43486 32226 43538
rect 32226 43486 32228 43538
rect 32172 43484 32228 43486
rect 32060 43148 32116 43204
rect 33516 44156 33572 44212
rect 32956 43596 33012 43652
rect 33404 43650 33460 43652
rect 33404 43598 33406 43650
rect 33406 43598 33458 43650
rect 33458 43598 33460 43650
rect 33404 43596 33460 43598
rect 32620 42924 32676 42980
rect 33236 43372 33292 43428
rect 33068 43148 33124 43204
rect 33516 43036 33572 43092
rect 32788 42812 32844 42868
rect 32956 42754 33012 42756
rect 31724 41692 31780 41748
rect 31836 42476 31892 42532
rect 32004 41580 32060 41636
rect 32956 42702 32958 42754
rect 32958 42702 33010 42754
rect 33010 42702 33012 42754
rect 32956 42700 33012 42702
rect 32508 42476 32564 42532
rect 32620 41580 32676 41636
rect 33180 42924 33236 42980
rect 32060 40796 32116 40852
rect 31612 40124 31668 40180
rect 29596 38220 29652 38276
rect 30268 38444 30324 38500
rect 29260 38108 29316 38164
rect 29596 38022 29652 38052
rect 29596 37996 29598 38022
rect 29598 37996 29650 38022
rect 29650 37996 29652 38022
rect 29372 37884 29428 37940
rect 29820 37772 29876 37828
rect 29260 37266 29316 37268
rect 29260 37214 29262 37266
rect 29262 37214 29314 37266
rect 29314 37214 29316 37266
rect 29260 37212 29316 37214
rect 29820 37212 29876 37268
rect 29596 36428 29652 36484
rect 29316 36370 29372 36372
rect 29316 36318 29318 36370
rect 29318 36318 29370 36370
rect 29370 36318 29372 36370
rect 29316 36316 29372 36318
rect 29260 35532 29316 35588
rect 29372 35420 29428 35476
rect 29372 34748 29428 34804
rect 29148 34300 29204 34356
rect 29036 33292 29092 33348
rect 29260 32620 29316 32676
rect 28588 30828 28644 30884
rect 30380 37772 30436 37828
rect 30604 38050 30660 38052
rect 30604 37998 30606 38050
rect 30606 37998 30658 38050
rect 30658 37998 30660 38050
rect 30604 37996 30660 37998
rect 30828 38444 30884 38500
rect 31612 39116 31668 39172
rect 31724 39004 31780 39060
rect 31948 38892 32004 38948
rect 32172 38810 32174 38836
rect 32174 38810 32226 38836
rect 32226 38810 32228 38836
rect 32172 38780 32228 38810
rect 31780 38444 31836 38500
rect 31612 38332 31668 38388
rect 31332 37884 31388 37940
rect 32172 38220 32228 38276
rect 30380 36876 30436 36932
rect 30492 36540 30548 36596
rect 30828 37266 30884 37268
rect 30828 37214 30830 37266
rect 30830 37214 30882 37266
rect 30882 37214 30884 37266
rect 30828 37212 30884 37214
rect 30380 35980 30436 36036
rect 31220 35980 31276 36036
rect 30660 35586 30716 35588
rect 30660 35534 30662 35586
rect 30662 35534 30714 35586
rect 30714 35534 30716 35586
rect 30660 35532 30716 35534
rect 29596 34300 29652 34356
rect 29820 34300 29876 34356
rect 30044 34412 30100 34468
rect 29708 33346 29764 33348
rect 29708 33294 29710 33346
rect 29710 33294 29762 33346
rect 29762 33294 29764 33346
rect 29708 33292 29764 33294
rect 29820 32284 29876 32340
rect 29484 31276 29540 31332
rect 28700 30210 28756 30212
rect 28700 30158 28702 30210
rect 28702 30158 28754 30210
rect 28754 30158 28756 30210
rect 28700 30156 28756 30158
rect 28924 29820 28980 29876
rect 29036 30994 29092 30996
rect 29036 30942 29038 30994
rect 29038 30942 29090 30994
rect 29090 30942 29092 30994
rect 29036 30940 29092 30942
rect 30268 34354 30324 34356
rect 30268 34302 30270 34354
rect 30270 34302 30322 34354
rect 30322 34302 30324 34354
rect 30268 34300 30324 34302
rect 31892 37378 31948 37380
rect 31892 37326 31894 37378
rect 31894 37326 31946 37378
rect 31946 37326 31948 37378
rect 31892 37324 31948 37326
rect 32060 36988 32116 37044
rect 31724 36594 31780 36596
rect 31724 36542 31726 36594
rect 31726 36542 31778 36594
rect 31778 36542 31780 36594
rect 31724 36540 31780 36542
rect 31612 36092 31668 36148
rect 32060 35980 32116 36036
rect 31948 34972 32004 35028
rect 31500 34748 31556 34804
rect 31724 34802 31780 34804
rect 31724 34750 31726 34802
rect 31726 34750 31778 34802
rect 31778 34750 31780 34802
rect 31724 34748 31780 34750
rect 31668 34412 31724 34468
rect 31612 32732 31668 32788
rect 31052 32620 31108 32676
rect 30380 32060 30436 32116
rect 30380 31500 30436 31556
rect 30380 31218 30436 31220
rect 30380 31166 30382 31218
rect 30382 31166 30434 31218
rect 30434 31166 30436 31218
rect 30380 31164 30436 31166
rect 31948 32338 32004 32340
rect 31948 32286 31950 32338
rect 31950 32286 32002 32338
rect 32002 32286 32004 32338
rect 31948 32284 32004 32286
rect 32172 32284 32228 32340
rect 32566 39228 32622 39284
rect 32508 37996 32564 38052
rect 33796 42812 33852 42868
rect 34076 42754 34132 42756
rect 34076 42702 34078 42754
rect 34078 42702 34130 42754
rect 34130 42702 34132 42754
rect 34076 42700 34132 42702
rect 34392 44716 34448 44772
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 34392 44322 34448 44324
rect 34392 44270 34394 44322
rect 34394 44270 34446 44322
rect 34446 44270 34448 44322
rect 34392 44268 34448 44270
rect 35196 44284 35252 44324
rect 35196 44268 35198 44284
rect 35198 44268 35250 44284
rect 35250 44268 35252 44284
rect 34748 44156 34804 44212
rect 35532 44156 35588 44212
rect 36316 47180 36372 47236
rect 36932 47234 36988 47236
rect 36932 47182 36934 47234
rect 36934 47182 36986 47234
rect 36986 47182 36988 47234
rect 36932 47180 36988 47182
rect 36652 46562 36708 46564
rect 36652 46510 36654 46562
rect 36654 46510 36706 46562
rect 36706 46510 36708 46562
rect 36652 46508 36708 46510
rect 36316 45836 36372 45892
rect 36092 45724 36148 45780
rect 36484 45276 36540 45332
rect 36316 45164 36372 45220
rect 36876 45890 36932 45892
rect 36876 45838 36878 45890
rect 36878 45838 36930 45890
rect 36930 45838 36932 45890
rect 36876 45836 36932 45838
rect 38276 47458 38332 47460
rect 38276 47406 38278 47458
rect 38278 47406 38330 47458
rect 38330 47406 38332 47458
rect 38276 47404 38332 47406
rect 41916 47292 41972 47348
rect 40572 47068 40628 47124
rect 36204 44940 36260 44996
rect 36876 45276 36932 45332
rect 36540 44828 36596 44884
rect 34748 43372 34804 43428
rect 34468 42812 34524 42868
rect 34524 42588 34580 42644
rect 34972 43260 35028 43316
rect 35644 43484 35700 43540
rect 35532 43260 35588 43316
rect 35756 43372 35812 43428
rect 36428 43708 36484 43764
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 34748 42364 34804 42420
rect 35028 42588 35084 42644
rect 35420 42812 35476 42868
rect 35644 42812 35700 42868
rect 35308 42476 35364 42532
rect 34972 42364 35028 42420
rect 33292 41186 33348 41188
rect 33292 41134 33294 41186
rect 33294 41134 33346 41186
rect 33346 41134 33348 41186
rect 33292 41132 33348 41134
rect 33628 41132 33684 41188
rect 33068 40572 33124 40628
rect 32956 38220 33012 38276
rect 33068 40236 33124 40292
rect 32956 38050 33012 38052
rect 32956 37998 32958 38050
rect 32958 37998 33010 38050
rect 33010 37998 33012 38050
rect 32956 37996 33012 37998
rect 32396 37378 32452 37380
rect 32396 37326 32398 37378
rect 32398 37326 32450 37378
rect 32450 37326 32452 37378
rect 32396 37324 32452 37326
rect 32620 36988 32676 37044
rect 32284 36652 32340 36708
rect 34076 41244 34132 41300
rect 33292 40236 33348 40292
rect 33348 39116 33404 39172
rect 33180 39004 33236 39060
rect 34468 40626 34524 40628
rect 34468 40574 34470 40626
rect 34470 40574 34522 40626
rect 34522 40574 34524 40626
rect 34468 40572 34524 40574
rect 34860 40402 34916 40404
rect 34860 40350 34862 40402
rect 34862 40350 34914 40402
rect 34914 40350 34916 40402
rect 34860 40348 34916 40350
rect 34076 40012 34132 40068
rect 35252 42252 35308 42308
rect 35252 41858 35308 41860
rect 35252 41806 35254 41858
rect 35254 41806 35306 41858
rect 35306 41806 35308 41858
rect 35252 41804 35308 41806
rect 36092 42588 36148 42644
rect 36092 42364 36148 42420
rect 35980 42028 36036 42084
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35196 41298 35252 41300
rect 35196 41246 35198 41298
rect 35198 41246 35250 41298
rect 35250 41246 35252 41298
rect 35196 41244 35252 41246
rect 35196 40684 35252 40740
rect 35308 40236 35364 40292
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35420 39788 35476 39844
rect 34972 39603 35028 39620
rect 34972 39564 34974 39603
rect 34974 39564 35026 39603
rect 35026 39564 35028 39603
rect 35420 39618 35476 39620
rect 35420 39566 35422 39618
rect 35422 39566 35474 39618
rect 35474 39566 35476 39618
rect 35420 39564 35476 39566
rect 33796 39228 33852 39284
rect 33516 38892 33572 38948
rect 33180 38834 33236 38836
rect 33180 38782 33182 38834
rect 33182 38782 33234 38834
rect 33234 38782 33236 38834
rect 33180 38780 33236 38782
rect 33292 38668 33348 38724
rect 33740 38556 33796 38612
rect 33964 38444 34020 38500
rect 34860 38780 34916 38836
rect 35084 38722 35140 38724
rect 35084 38670 35086 38722
rect 35086 38670 35138 38722
rect 35138 38670 35140 38722
rect 35084 38668 35140 38670
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 33908 37826 33964 37828
rect 33908 37774 33910 37826
rect 33910 37774 33962 37826
rect 33962 37774 33964 37826
rect 33908 37772 33964 37774
rect 33292 37266 33348 37268
rect 33292 37214 33294 37266
rect 33294 37214 33346 37266
rect 33346 37214 33348 37266
rect 33292 37212 33348 37214
rect 33292 36876 33348 36932
rect 32508 35868 32564 35924
rect 32396 34972 32452 35028
rect 32452 34188 32508 34244
rect 33180 36482 33236 36484
rect 33180 36430 33182 36482
rect 33182 36430 33234 36482
rect 33234 36430 33236 36482
rect 33180 36428 33236 36430
rect 32732 35644 32788 35700
rect 33180 35698 33236 35700
rect 33180 35646 33182 35698
rect 33182 35646 33234 35698
rect 33234 35646 33236 35698
rect 33180 35644 33236 35646
rect 33852 36764 33908 36820
rect 33628 36092 33684 36148
rect 33404 35644 33460 35700
rect 32956 34972 33012 35028
rect 33516 34972 33572 35028
rect 33516 34748 33572 34804
rect 33404 34636 33460 34692
rect 33740 34972 33796 35028
rect 33852 34748 33908 34804
rect 34468 37548 34524 37604
rect 34168 37324 34224 37380
rect 35644 41804 35700 41860
rect 35868 41804 35924 41860
rect 35644 41580 35700 41636
rect 36204 41916 36260 41972
rect 36652 42364 36708 42420
rect 36540 42028 36596 42084
rect 36428 41468 36484 41524
rect 38332 45276 38388 45332
rect 38220 45164 38276 45220
rect 37044 45106 37100 45108
rect 37044 45054 37046 45106
rect 37046 45054 37098 45106
rect 37098 45054 37100 45106
rect 37044 45052 37100 45054
rect 37996 44828 38052 44884
rect 37772 44716 37828 44772
rect 37324 44156 37380 44212
rect 36988 42812 37044 42868
rect 37100 43708 37156 43764
rect 37212 43260 37268 43316
rect 38556 45106 38612 45108
rect 38556 45054 38558 45106
rect 38558 45054 38610 45106
rect 38610 45054 38612 45106
rect 38556 45052 38612 45054
rect 38668 44828 38724 44884
rect 38220 43708 38276 43764
rect 36876 41692 36932 41748
rect 37548 42924 37604 42980
rect 38556 43484 38612 43540
rect 39508 44828 39564 44884
rect 39340 44716 39396 44772
rect 40012 46674 40068 46676
rect 40012 46622 40014 46674
rect 40014 46622 40066 46674
rect 40066 46622 40068 46674
rect 40012 46620 40068 46622
rect 40460 45724 40516 45780
rect 39956 45330 40012 45332
rect 39956 45278 39958 45330
rect 39958 45278 40010 45330
rect 40010 45278 40012 45330
rect 39956 45276 40012 45278
rect 39676 44604 39732 44660
rect 40236 45052 40292 45108
rect 39340 43820 39396 43876
rect 40460 44434 40516 44436
rect 40460 44382 40462 44434
rect 40462 44382 40514 44434
rect 40514 44382 40516 44434
rect 40460 44380 40516 44382
rect 38108 42754 38164 42756
rect 38108 42702 38110 42754
rect 38110 42702 38162 42754
rect 38162 42702 38164 42754
rect 38108 42700 38164 42702
rect 37324 42364 37380 42420
rect 37436 41970 37492 41972
rect 37436 41918 37438 41970
rect 37438 41918 37490 41970
rect 37490 41918 37492 41970
rect 37436 41916 37492 41918
rect 36988 41580 37044 41636
rect 38220 41580 38276 41636
rect 36428 40572 36484 40628
rect 35980 40236 36036 40292
rect 35644 38892 35700 38948
rect 35308 37100 35364 37156
rect 35196 36988 35252 37044
rect 36540 40124 36596 40180
rect 36540 39564 36596 39620
rect 35980 38834 36036 38836
rect 35980 38782 35982 38834
rect 35982 38782 36034 38834
rect 36034 38782 36036 38834
rect 35980 38780 36036 38782
rect 36092 38668 36148 38724
rect 35756 38556 35812 38612
rect 35532 37548 35588 37604
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35532 36092 35588 36148
rect 36316 38610 36372 38612
rect 36316 38558 36318 38610
rect 36318 38558 36370 38610
rect 36370 38558 36372 38610
rect 36316 38556 36372 38558
rect 36372 38050 36428 38052
rect 36372 37998 36374 38050
rect 36374 37998 36426 38050
rect 36426 37998 36428 38050
rect 36372 37996 36428 37998
rect 36092 37324 36148 37380
rect 36148 37154 36204 37156
rect 36148 37102 36150 37154
rect 36150 37102 36202 37154
rect 36202 37102 36204 37154
rect 36148 37100 36204 37102
rect 35644 36428 35700 36484
rect 35420 35922 35476 35924
rect 35420 35870 35422 35922
rect 35422 35870 35474 35922
rect 35474 35870 35476 35922
rect 35420 35868 35476 35870
rect 36204 36092 36260 36148
rect 34076 35026 34132 35028
rect 34076 34974 34078 35026
rect 34078 34974 34130 35026
rect 34130 34974 34132 35026
rect 34076 34972 34132 34974
rect 34076 34748 34132 34804
rect 33852 34300 33908 34356
rect 34412 35308 34468 35364
rect 34300 34636 34356 34692
rect 33740 33964 33796 34020
rect 32564 32674 32620 32676
rect 32564 32622 32566 32674
rect 32566 32622 32618 32674
rect 32618 32622 32620 32674
rect 32564 32620 32620 32622
rect 32396 32284 32452 32340
rect 30044 30828 30100 30884
rect 28588 29596 28644 29652
rect 28476 29148 28532 29204
rect 28476 28924 28532 28980
rect 28140 28700 28196 28756
rect 28812 28588 28868 28644
rect 27916 28028 27972 28084
rect 28924 28364 28980 28420
rect 29372 28924 29428 28980
rect 29036 28140 29092 28196
rect 27916 27580 27972 27636
rect 27804 27244 27860 27300
rect 27356 27074 27412 27076
rect 27356 27022 27358 27074
rect 27358 27022 27410 27074
rect 27410 27022 27412 27074
rect 27356 27020 27412 27022
rect 28084 27074 28140 27076
rect 28084 27022 28086 27074
rect 28086 27022 28138 27074
rect 28138 27022 28140 27074
rect 28084 27020 28140 27022
rect 27020 26908 27076 26964
rect 27020 26124 27076 26180
rect 27580 25452 27636 25508
rect 27804 26236 27860 26292
rect 27916 26124 27972 26180
rect 26796 25116 26852 25172
rect 26684 24892 26740 24948
rect 25452 21868 25508 21924
rect 25228 20972 25284 21028
rect 25340 20860 25396 20916
rect 24780 20748 24836 20804
rect 24052 20130 24108 20132
rect 24052 20078 24054 20130
rect 24054 20078 24106 20130
rect 24106 20078 24108 20130
rect 24052 20076 24108 20078
rect 23492 19852 23548 19908
rect 24444 19794 24500 19796
rect 24444 19742 24446 19794
rect 24446 19742 24498 19794
rect 24498 19742 24500 19794
rect 24444 19740 24500 19742
rect 24892 20076 24948 20132
rect 23884 19122 23940 19124
rect 23884 19070 23886 19122
rect 23886 19070 23938 19122
rect 23938 19070 23940 19122
rect 23884 19068 23940 19070
rect 23436 18396 23492 18452
rect 23100 17666 23156 17668
rect 23100 17614 23102 17666
rect 23102 17614 23154 17666
rect 23154 17614 23156 17666
rect 23100 17612 23156 17614
rect 24220 18450 24276 18452
rect 24220 18398 24222 18450
rect 24222 18398 24274 18450
rect 24274 18398 24276 18450
rect 24220 18396 24276 18398
rect 24052 17836 24108 17892
rect 23772 17666 23828 17668
rect 23772 17614 23774 17666
rect 23774 17614 23826 17666
rect 23826 17614 23828 17666
rect 23772 17612 23828 17614
rect 24332 17612 24388 17668
rect 23100 17052 23156 17108
rect 22764 16716 22820 16772
rect 23660 17554 23716 17556
rect 23660 17502 23662 17554
rect 23662 17502 23714 17554
rect 23714 17502 23716 17554
rect 23660 17500 23716 17502
rect 23660 17276 23716 17332
rect 23548 17052 23604 17108
rect 23436 16994 23492 16996
rect 23436 16942 23438 16994
rect 23438 16942 23490 16994
rect 23490 16942 23492 16994
rect 23436 16940 23492 16942
rect 23324 16716 23380 16772
rect 22988 16098 23044 16100
rect 22988 16046 22990 16098
rect 22990 16046 23042 16098
rect 23042 16046 23044 16098
rect 22988 16044 23044 16046
rect 22988 15484 23044 15540
rect 22764 15372 22820 15428
rect 23324 16044 23380 16100
rect 24108 17052 24164 17108
rect 27244 25116 27300 25172
rect 27132 24556 27188 24612
rect 25900 24220 25956 24276
rect 25732 24050 25788 24052
rect 25732 23998 25734 24050
rect 25734 23998 25786 24050
rect 25786 23998 25788 24050
rect 25732 23996 25788 23998
rect 26684 24108 26740 24164
rect 26572 23910 26628 23940
rect 25732 23154 25788 23156
rect 25732 23102 25734 23154
rect 25734 23102 25786 23154
rect 25786 23102 25788 23154
rect 25732 23100 25788 23102
rect 26012 23130 26014 23156
rect 26014 23130 26066 23156
rect 26066 23130 26068 23156
rect 26012 23100 26068 23130
rect 26572 23884 26574 23910
rect 26574 23884 26626 23910
rect 26626 23884 26628 23910
rect 26348 23436 26404 23492
rect 27244 24108 27300 24164
rect 27356 23938 27412 23940
rect 27356 23886 27358 23938
rect 27358 23886 27410 23938
rect 27410 23886 27412 23938
rect 27356 23884 27412 23886
rect 26460 23212 26516 23268
rect 27020 23154 27076 23156
rect 27020 23102 27022 23154
rect 27022 23102 27074 23154
rect 27074 23102 27076 23154
rect 27020 23100 27076 23102
rect 26796 22988 26852 23044
rect 26572 22204 26628 22260
rect 25676 21586 25732 21588
rect 25676 21534 25678 21586
rect 25678 21534 25730 21586
rect 25730 21534 25732 21586
rect 25676 21532 25732 21534
rect 26964 21586 27020 21588
rect 26964 21534 26966 21586
rect 26966 21534 27018 21586
rect 27018 21534 27020 21586
rect 26964 21532 27020 21534
rect 25228 19993 25230 20020
rect 25230 19993 25282 20020
rect 25282 19993 25284 20020
rect 25228 19964 25284 19993
rect 24892 19234 24948 19236
rect 24892 19182 24894 19234
rect 24894 19182 24946 19234
rect 24946 19182 24948 19234
rect 24892 19180 24948 19182
rect 24556 18338 24612 18340
rect 24556 18286 24558 18338
rect 24558 18286 24610 18338
rect 24610 18286 24612 18338
rect 24556 18284 24612 18286
rect 24892 18284 24948 18340
rect 24780 17500 24836 17556
rect 24612 17276 24668 17332
rect 24220 16268 24276 16324
rect 24220 16098 24276 16100
rect 24220 16046 24222 16098
rect 24222 16046 24274 16098
rect 24274 16046 24276 16098
rect 24220 16044 24276 16046
rect 23212 15314 23268 15316
rect 23212 15262 23214 15314
rect 23214 15262 23266 15314
rect 23266 15262 23268 15314
rect 23212 15260 23268 15262
rect 22652 13132 22708 13188
rect 21924 12348 21980 12404
rect 20412 11676 20468 11732
rect 19740 11618 19796 11620
rect 19740 11566 19742 11618
rect 19742 11566 19794 11618
rect 19794 11566 19796 11618
rect 19740 11564 19796 11566
rect 20748 11564 20804 11620
rect 20412 11394 20468 11396
rect 20412 11342 20414 11394
rect 20414 11342 20466 11394
rect 20466 11342 20468 11394
rect 20412 11340 20468 11342
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 20338 10780 20394 10836
rect 20524 10668 20580 10724
rect 21420 11788 21476 11844
rect 23212 14364 23268 14420
rect 22988 13468 23044 13524
rect 23100 14028 23156 14084
rect 23436 14252 23492 14308
rect 23212 13356 23268 13412
rect 22876 12348 22932 12404
rect 23884 15596 23940 15652
rect 23660 15148 23716 15204
rect 23884 15314 23940 15316
rect 23884 15262 23886 15314
rect 23886 15262 23938 15314
rect 23938 15262 23940 15314
rect 23884 15260 23940 15262
rect 24724 15986 24780 15988
rect 24724 15934 24726 15986
rect 24726 15934 24778 15986
rect 24778 15934 24780 15986
rect 24724 15932 24780 15934
rect 25228 17724 25284 17780
rect 25564 19740 25620 19796
rect 25340 17388 25396 17444
rect 25452 17666 25508 17668
rect 25452 17614 25454 17666
rect 25454 17614 25506 17666
rect 25506 17614 25508 17666
rect 25452 17612 25508 17614
rect 26348 18508 26404 18564
rect 27804 22876 27860 22932
rect 28364 26796 28420 26852
rect 28588 27132 28644 27188
rect 29036 27074 29092 27076
rect 29036 27022 29038 27074
rect 29038 27022 29090 27074
rect 29090 27022 29092 27074
rect 29036 27020 29092 27022
rect 29708 28812 29764 28868
rect 29484 28642 29540 28644
rect 29484 28590 29486 28642
rect 29486 28590 29538 28642
rect 29538 28590 29540 28642
rect 29484 28588 29540 28590
rect 29372 28140 29428 28196
rect 29372 26962 29428 26964
rect 29372 26910 29374 26962
rect 29374 26910 29426 26962
rect 29426 26910 29428 26962
rect 29372 26908 29428 26910
rect 28140 23996 28196 24052
rect 28252 23938 28308 23940
rect 28252 23886 28254 23938
rect 28254 23886 28306 23938
rect 28306 23886 28308 23938
rect 28252 23884 28308 23886
rect 28140 23436 28196 23492
rect 27916 22540 27972 22596
rect 27804 22428 27860 22484
rect 27916 22342 27972 22372
rect 27916 22316 27918 22342
rect 27918 22316 27970 22342
rect 27970 22316 27972 22342
rect 27636 22258 27692 22260
rect 27636 22206 27638 22258
rect 27638 22206 27690 22258
rect 27690 22206 27692 22258
rect 27636 22204 27692 22206
rect 27468 21756 27524 21812
rect 28532 24444 28588 24500
rect 29036 25506 29092 25508
rect 29036 25454 29038 25506
rect 29038 25454 29090 25506
rect 29090 25454 29092 25506
rect 29036 25452 29092 25454
rect 28924 25340 28980 25396
rect 28588 23436 28644 23492
rect 28140 21756 28196 21812
rect 28476 22540 28532 22596
rect 27468 20076 27524 20132
rect 28700 23154 28756 23156
rect 28700 23102 28702 23154
rect 28702 23102 28754 23154
rect 28754 23102 28756 23154
rect 28700 23100 28756 23102
rect 28588 22092 28644 22148
rect 30044 28140 30100 28196
rect 29708 27244 29764 27300
rect 29484 25116 29540 25172
rect 30324 29036 30380 29092
rect 30380 27916 30436 27972
rect 31724 29932 31780 29988
rect 30604 29820 30660 29876
rect 31836 29820 31892 29876
rect 32172 31890 32228 31892
rect 32172 31838 32174 31890
rect 32174 31838 32226 31890
rect 32226 31838 32228 31890
rect 32172 31836 32228 31838
rect 33124 32732 33180 32788
rect 33628 32732 33684 32788
rect 33068 31948 33124 32004
rect 32396 31388 32452 31444
rect 32396 31164 32452 31220
rect 32284 30970 32286 30996
rect 32286 30970 32338 30996
rect 32338 30970 32340 30996
rect 32284 30940 32340 30970
rect 32508 30940 32564 30996
rect 33404 31388 33460 31444
rect 31948 29708 32004 29764
rect 30940 28700 30996 28756
rect 31164 28140 31220 28196
rect 31388 27916 31444 27972
rect 31276 27804 31332 27860
rect 30828 27692 30884 27748
rect 31836 28812 31892 28868
rect 32620 28364 32676 28420
rect 33628 32538 33630 32564
rect 33630 32538 33682 32564
rect 33682 32538 33684 32564
rect 33628 32508 33684 32538
rect 33852 33852 33908 33908
rect 34916 35308 34972 35364
rect 34412 33964 34468 34020
rect 34132 33906 34188 33908
rect 34132 33854 34134 33906
rect 34134 33854 34186 33906
rect 34186 33854 34188 33906
rect 34132 33852 34188 33854
rect 33964 33068 34020 33124
rect 33852 32732 33908 32788
rect 34860 32844 34916 32900
rect 34412 32732 34468 32788
rect 34188 32508 34244 32564
rect 34636 32538 34638 32564
rect 34638 32538 34690 32564
rect 34690 32538 34692 32564
rect 34636 32508 34692 32538
rect 34300 32284 34356 32340
rect 34300 32060 34356 32116
rect 34076 31836 34132 31892
rect 33516 30940 33572 30996
rect 33628 31052 33684 31108
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35532 34972 35588 35028
rect 35196 33852 35252 33908
rect 35644 33964 35700 34020
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35644 33180 35700 33236
rect 35756 33516 35812 33572
rect 35756 32844 35812 32900
rect 35532 32732 35588 32788
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35532 31948 35588 32004
rect 34188 31388 34244 31444
rect 34748 31052 34804 31108
rect 33404 30268 33460 30324
rect 33292 30210 33348 30212
rect 33292 30158 33294 30210
rect 33294 30158 33346 30210
rect 33346 30158 33348 30210
rect 33292 30156 33348 30158
rect 32732 29708 32788 29764
rect 32844 28700 32900 28756
rect 32508 28140 32564 28196
rect 31612 27692 31668 27748
rect 30772 27298 30828 27300
rect 30772 27246 30774 27298
rect 30774 27246 30826 27298
rect 30826 27246 30828 27298
rect 30772 27244 30828 27246
rect 31836 27074 31892 27076
rect 31836 27022 31838 27074
rect 31838 27022 31890 27074
rect 31890 27022 31892 27074
rect 31836 27020 31892 27022
rect 32060 27858 32116 27860
rect 32060 27806 32062 27858
rect 32062 27806 32114 27858
rect 32114 27806 32116 27858
rect 32060 27804 32116 27806
rect 32340 27186 32396 27188
rect 32340 27134 32342 27186
rect 32342 27134 32394 27186
rect 32394 27134 32396 27186
rect 32340 27132 32396 27134
rect 32620 27074 32676 27076
rect 32620 27022 32622 27074
rect 32622 27022 32674 27074
rect 32674 27022 32676 27074
rect 32620 27020 32676 27022
rect 31052 26348 31108 26404
rect 31388 26572 31444 26628
rect 32284 26402 32340 26404
rect 32284 26350 32286 26402
rect 32286 26350 32338 26402
rect 32338 26350 32340 26402
rect 32284 26348 32340 26350
rect 31724 26276 31726 26292
rect 31726 26276 31778 26292
rect 31778 26276 31780 26292
rect 31724 26236 31780 26276
rect 30604 25788 30660 25844
rect 30044 25340 30100 25396
rect 30940 25340 30996 25396
rect 31164 25788 31220 25844
rect 30716 25228 30772 25284
rect 30044 25116 30100 25172
rect 29708 24444 29764 24500
rect 29932 24892 29988 24948
rect 29596 23436 29652 23492
rect 29708 23100 29764 23156
rect 29820 23324 29876 23380
rect 29316 22482 29372 22484
rect 29316 22430 29318 22482
rect 29318 22430 29370 22482
rect 29370 22430 29372 22482
rect 29316 22428 29372 22430
rect 31052 25228 31108 25284
rect 30940 24780 30996 24836
rect 30044 23212 30100 23268
rect 30380 23436 30436 23492
rect 29932 22428 29988 22484
rect 29484 22370 29540 22372
rect 29484 22318 29486 22370
rect 29486 22318 29538 22370
rect 29538 22318 29540 22370
rect 29484 22316 29540 22318
rect 29708 21756 29764 21812
rect 29484 21196 29540 21252
rect 28700 20802 28756 20804
rect 28700 20750 28702 20802
rect 28702 20750 28754 20802
rect 28754 20750 28756 20802
rect 28700 20748 28756 20750
rect 28252 20076 28308 20132
rect 27580 19516 27636 19572
rect 27356 19404 27412 19460
rect 27132 18396 27188 18452
rect 28140 19404 28196 19460
rect 28812 20076 28868 20132
rect 28364 19516 28420 19572
rect 29204 20802 29260 20804
rect 29204 20750 29206 20802
rect 29206 20750 29258 20802
rect 29258 20750 29260 20802
rect 29204 20748 29260 20750
rect 29988 21756 30044 21812
rect 30156 22092 30212 22148
rect 30268 21868 30324 21924
rect 29820 21308 29876 21364
rect 29596 20524 29652 20580
rect 29148 20300 29204 20356
rect 29484 20130 29540 20132
rect 29484 20078 29486 20130
rect 29486 20078 29538 20130
rect 29538 20078 29540 20130
rect 29484 20076 29540 20078
rect 29260 19852 29316 19908
rect 28924 19628 28980 19684
rect 28588 19292 28644 19348
rect 28252 19180 28308 19236
rect 30044 20300 30100 20356
rect 30268 20188 30324 20244
rect 30548 22540 30604 22596
rect 30548 22146 30604 22148
rect 30548 22094 30550 22146
rect 30550 22094 30602 22146
rect 30602 22094 30604 22146
rect 30548 22092 30604 22094
rect 30604 21868 30660 21924
rect 30492 21308 30548 21364
rect 30884 22930 30940 22932
rect 30884 22878 30886 22930
rect 30886 22878 30938 22930
rect 30938 22878 30940 22930
rect 30884 22876 30940 22878
rect 30716 21532 30772 21588
rect 30940 21756 30996 21812
rect 31164 24780 31220 24836
rect 31407 24780 31463 24836
rect 31276 24668 31332 24724
rect 32508 25340 32564 25396
rect 32340 25282 32396 25284
rect 32340 25230 32342 25282
rect 32342 25230 32394 25282
rect 32394 25230 32396 25282
rect 32340 25228 32396 25230
rect 33572 29650 33628 29652
rect 33572 29598 33574 29650
rect 33574 29598 33626 29650
rect 33626 29598 33628 29650
rect 33572 29596 33628 29598
rect 34076 29820 34132 29876
rect 33516 29372 33572 29428
rect 33348 28866 33404 28868
rect 33348 28814 33350 28866
rect 33350 28814 33402 28866
rect 33402 28814 33404 28866
rect 33348 28812 33404 28814
rect 33068 28642 33124 28644
rect 33068 28590 33070 28642
rect 33070 28590 33122 28642
rect 33122 28590 33124 28642
rect 33068 28588 33124 28590
rect 33516 28588 33572 28644
rect 33628 29260 33684 29316
rect 32956 24892 33012 24948
rect 32788 24780 32844 24836
rect 31164 23884 31220 23940
rect 31612 24668 31668 24724
rect 32284 24722 32340 24724
rect 32284 24670 32286 24722
rect 32286 24670 32338 24722
rect 32338 24670 32340 24722
rect 32284 24668 32340 24670
rect 32620 23996 32676 24052
rect 33404 27858 33460 27860
rect 33404 27806 33406 27858
rect 33406 27806 33458 27858
rect 33458 27806 33460 27858
rect 33404 27804 33460 27806
rect 34300 30044 34356 30100
rect 34300 29596 34356 29652
rect 34300 29401 34302 29428
rect 34302 29401 34354 29428
rect 34354 29401 34356 29428
rect 34300 29372 34356 29401
rect 34636 29426 34692 29428
rect 34636 29374 34638 29426
rect 34638 29374 34690 29426
rect 34690 29374 34692 29426
rect 34636 29372 34692 29374
rect 34188 29260 34244 29316
rect 33852 28364 33908 28420
rect 33964 28700 34020 28756
rect 34524 28603 34580 28644
rect 34524 28588 34526 28603
rect 34526 28588 34578 28603
rect 34578 28588 34580 28603
rect 33740 27858 33796 27860
rect 33740 27806 33742 27858
rect 33742 27806 33794 27858
rect 33794 27806 33796 27858
rect 33740 27804 33796 27806
rect 34244 28252 34300 28308
rect 36540 36482 36596 36484
rect 36540 36430 36542 36482
rect 36542 36430 36594 36482
rect 36594 36430 36596 36482
rect 36540 36428 36596 36430
rect 36428 35196 36484 35252
rect 37156 40572 37212 40628
rect 36764 40378 36766 40404
rect 36766 40378 36818 40404
rect 36818 40378 36820 40404
rect 36764 40348 36820 40378
rect 36988 40378 36990 40404
rect 36990 40378 37042 40404
rect 37042 40378 37044 40404
rect 36988 40348 37044 40378
rect 37436 40796 37492 40852
rect 37268 40514 37324 40516
rect 37268 40462 37270 40514
rect 37270 40462 37322 40514
rect 37322 40462 37324 40514
rect 37268 40460 37324 40462
rect 36764 40124 36820 40180
rect 36988 39583 37044 39620
rect 36988 39564 36990 39583
rect 36990 39564 37042 39583
rect 37042 39564 37044 39583
rect 36876 39116 36932 39172
rect 36764 39004 36820 39060
rect 36876 38892 36932 38948
rect 36764 38668 36820 38724
rect 36876 38050 36932 38052
rect 36876 37998 36878 38050
rect 36878 37998 36930 38050
rect 36930 37998 36932 38050
rect 36876 37996 36932 37998
rect 37100 39004 37156 39060
rect 37100 38780 37156 38836
rect 37324 40236 37380 40292
rect 37884 40572 37940 40628
rect 37548 39676 37604 39732
rect 38108 39676 38164 39732
rect 37772 39564 37828 39620
rect 37324 39004 37380 39060
rect 37100 35980 37156 36036
rect 37604 38834 37660 38836
rect 37604 38782 37606 38834
rect 37606 38782 37658 38834
rect 37658 38782 37660 38834
rect 37604 38780 37660 38782
rect 37436 38556 37492 38612
rect 37996 38834 38052 38836
rect 37996 38782 37998 38834
rect 37998 38782 38050 38834
rect 38050 38782 38052 38834
rect 37996 38780 38052 38782
rect 38332 41356 38388 41412
rect 39228 43148 39284 43204
rect 38668 42700 38724 42756
rect 40348 43596 40404 43652
rect 40460 43538 40516 43540
rect 40460 43486 40462 43538
rect 40462 43486 40514 43538
rect 40514 43486 40516 43538
rect 40460 43484 40516 43486
rect 40348 42028 40404 42084
rect 39116 41356 39172 41412
rect 39340 41858 39396 41860
rect 39340 41806 39342 41858
rect 39342 41806 39394 41858
rect 39394 41806 39396 41858
rect 39340 41804 39396 41806
rect 38780 40572 38836 40628
rect 39340 40572 39396 40628
rect 40236 41916 40292 41972
rect 39900 40908 39956 40964
rect 39676 40460 39732 40516
rect 40124 40684 40180 40740
rect 40236 40796 40292 40852
rect 38668 39788 38724 39844
rect 38444 39116 38500 39172
rect 38948 38722 39004 38724
rect 38948 38670 38950 38722
rect 38950 38670 39002 38722
rect 39002 38670 39004 38722
rect 38948 38668 39004 38670
rect 39116 37772 39172 37828
rect 37828 35980 37884 36036
rect 37324 35698 37380 35700
rect 37324 35646 37326 35698
rect 37326 35646 37378 35698
rect 37378 35646 37380 35698
rect 37324 35644 37380 35646
rect 37324 35420 37380 35476
rect 36932 34748 36988 34804
rect 36764 34412 36820 34468
rect 36652 34300 36708 34356
rect 37100 33740 37156 33796
rect 36372 33122 36428 33124
rect 36372 33070 36374 33122
rect 36374 33070 36426 33122
rect 36426 33070 36428 33122
rect 36372 33068 36428 33070
rect 36540 33068 36596 33124
rect 36316 32732 36372 32788
rect 35756 31388 35812 31444
rect 35476 30770 35532 30772
rect 35476 30718 35478 30770
rect 35478 30718 35530 30770
rect 35530 30718 35532 30770
rect 35476 30716 35532 30718
rect 36764 32956 36820 33012
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 34972 29932 35028 29988
rect 35308 30156 35364 30212
rect 35532 30044 35588 30100
rect 35364 29650 35420 29652
rect 35364 29598 35366 29650
rect 35366 29598 35418 29650
rect 35418 29598 35420 29650
rect 35364 29596 35420 29598
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35644 28812 35700 28868
rect 34972 28364 35028 28420
rect 33852 27692 33908 27748
rect 33292 27020 33348 27076
rect 33516 27074 33572 27076
rect 33516 27022 33518 27074
rect 33518 27022 33570 27074
rect 33570 27022 33572 27074
rect 33516 27020 33572 27022
rect 34188 27074 34244 27076
rect 34188 27022 34190 27074
rect 34190 27022 34242 27074
rect 34242 27022 34244 27074
rect 34188 27020 34244 27022
rect 34468 27074 34524 27076
rect 34468 27022 34470 27074
rect 34470 27022 34522 27074
rect 34522 27022 34524 27074
rect 34468 27020 34524 27022
rect 34076 26908 34132 26964
rect 34748 27074 34804 27076
rect 34748 27022 34750 27074
rect 34750 27022 34802 27074
rect 34802 27022 34804 27074
rect 34748 27020 34804 27022
rect 33852 26796 33908 26852
rect 33572 26066 33628 26068
rect 33572 26014 33574 26066
rect 33574 26014 33626 26066
rect 33626 26014 33628 26066
rect 33572 26012 33628 26014
rect 34188 26684 34244 26740
rect 34076 26276 34078 26292
rect 34078 26276 34130 26292
rect 34130 26276 34132 26292
rect 34076 26236 34132 26276
rect 33516 25340 33572 25396
rect 33180 25228 33236 25284
rect 35084 27692 35140 27748
rect 34860 26684 34916 26740
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35084 26908 35140 26964
rect 33180 24946 33236 24948
rect 33180 24894 33182 24946
rect 33182 24894 33234 24946
rect 33234 24894 33236 24946
rect 33180 24892 33236 24894
rect 34076 24722 34132 24724
rect 34076 24670 34078 24722
rect 34078 24670 34130 24722
rect 34130 24670 34132 24722
rect 34076 24668 34132 24670
rect 34748 25506 34804 25508
rect 34748 25454 34750 25506
rect 34750 25454 34802 25506
rect 34802 25454 34804 25506
rect 34748 25452 34804 25454
rect 35084 26012 35140 26068
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35308 25506 35364 25508
rect 35308 25454 35310 25506
rect 35310 25454 35362 25506
rect 35362 25454 35364 25506
rect 35308 25452 35364 25454
rect 34916 25340 34972 25396
rect 35308 25228 35364 25284
rect 34636 24668 34692 24724
rect 33516 24444 33572 24500
rect 34076 24050 34132 24052
rect 34076 23998 34078 24050
rect 34078 23998 34130 24050
rect 34130 23998 34132 24050
rect 34076 23996 34132 23998
rect 31724 23436 31780 23492
rect 32172 23324 32228 23380
rect 32956 23324 33012 23380
rect 31668 23154 31724 23156
rect 31668 23102 31670 23154
rect 31670 23102 31722 23154
rect 31722 23102 31724 23154
rect 31668 23100 31724 23102
rect 32396 23212 32452 23268
rect 32620 23212 32676 23268
rect 32956 23154 33012 23156
rect 31164 22988 31220 23044
rect 32956 23102 32958 23154
rect 32958 23102 33010 23154
rect 33010 23102 33012 23154
rect 32956 23100 33012 23102
rect 33516 23100 33572 23156
rect 31948 22988 32004 23044
rect 31500 22876 31556 22932
rect 30716 20860 30772 20916
rect 29596 19404 29652 19460
rect 29708 19740 29764 19796
rect 29484 19292 29540 19348
rect 29260 19206 29316 19236
rect 29260 19180 29262 19206
rect 29262 19180 29314 19206
rect 29314 19180 29316 19206
rect 30380 19740 30436 19796
rect 30156 19628 30212 19684
rect 30156 19404 30212 19460
rect 28588 19068 28644 19124
rect 27916 18508 27972 18564
rect 28028 18732 28084 18788
rect 27356 18284 27412 18340
rect 27692 18338 27748 18340
rect 27692 18286 27694 18338
rect 27694 18286 27746 18338
rect 27746 18286 27748 18338
rect 27692 18284 27748 18286
rect 26348 17724 26404 17780
rect 25564 17164 25620 17220
rect 25676 16156 25732 16212
rect 25788 17388 25844 17444
rect 25116 15932 25172 15988
rect 24668 15596 24724 15652
rect 24500 15538 24556 15540
rect 24500 15486 24502 15538
rect 24502 15486 24554 15538
rect 24554 15486 24556 15538
rect 24500 15484 24556 15486
rect 24332 15372 24388 15428
rect 24668 13692 24724 13748
rect 24108 13468 24164 13524
rect 24892 15148 24948 15204
rect 25564 16044 25620 16100
rect 25452 15090 25508 15092
rect 25452 15038 25454 15090
rect 25454 15038 25506 15090
rect 25506 15038 25508 15090
rect 25452 15036 25508 15038
rect 26796 17666 26852 17668
rect 26796 17614 26798 17666
rect 26798 17614 26850 17666
rect 26850 17614 26852 17666
rect 26796 17612 26852 17614
rect 26630 17276 26686 17332
rect 27020 17612 27076 17668
rect 27244 17388 27300 17444
rect 27020 17052 27076 17108
rect 27132 17164 27188 17220
rect 26796 16882 26852 16884
rect 26796 16830 26798 16882
rect 26798 16830 26850 16882
rect 26850 16830 26852 16882
rect 26796 16828 26852 16830
rect 26964 16882 27020 16884
rect 26964 16830 26966 16882
rect 26966 16830 27018 16882
rect 27018 16830 27020 16882
rect 26964 16828 27020 16830
rect 27542 17276 27598 17332
rect 27356 17052 27412 17108
rect 27692 17164 27748 17220
rect 27916 16828 27972 16884
rect 26012 15260 26068 15316
rect 26236 15314 26292 15316
rect 26236 15262 26238 15314
rect 26238 15262 26290 15314
rect 26290 15262 26292 15314
rect 26236 15260 26292 15262
rect 25340 13746 25396 13748
rect 25340 13694 25342 13746
rect 25342 13694 25394 13746
rect 25394 13694 25396 13746
rect 25340 13692 25396 13694
rect 25228 13356 25284 13412
rect 24780 13244 24836 13300
rect 25452 13020 25508 13076
rect 21084 11564 21140 11620
rect 21980 11394 22036 11396
rect 21980 11342 21982 11394
rect 21982 11342 22034 11394
rect 22034 11342 22036 11394
rect 21980 11340 22036 11342
rect 22092 11228 22148 11284
rect 21678 10780 21734 10836
rect 20972 10668 21028 10724
rect 21532 10668 21588 10724
rect 20636 10610 20692 10612
rect 20636 10558 20638 10610
rect 20638 10558 20690 10610
rect 20690 10558 20692 10610
rect 20636 10556 20692 10558
rect 19292 10444 19348 10500
rect 21420 10444 21476 10500
rect 19292 9826 19348 9828
rect 19292 9774 19294 9826
rect 19294 9774 19346 9826
rect 19346 9774 19348 9826
rect 19292 9772 19348 9774
rect 20412 10332 20468 10388
rect 21980 10668 22036 10724
rect 20188 10220 20244 10276
rect 22652 9884 22708 9940
rect 22092 9826 22148 9828
rect 22092 9774 22094 9826
rect 22094 9774 22146 9826
rect 22146 9774 22148 9826
rect 22092 9772 22148 9774
rect 19516 9714 19572 9716
rect 19516 9662 19518 9714
rect 19518 9662 19570 9714
rect 19570 9662 19572 9714
rect 19516 9660 19572 9662
rect 20636 9714 20692 9716
rect 20636 9662 20638 9714
rect 20638 9662 20690 9714
rect 20690 9662 20692 9714
rect 20636 9660 20692 9662
rect 21308 9660 21364 9716
rect 19404 9212 19460 9268
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 20636 9436 20692 9492
rect 18284 8876 18340 8932
rect 17612 8540 17668 8596
rect 15932 5869 15934 5908
rect 15934 5869 15986 5908
rect 15986 5869 15988 5908
rect 15932 5852 15988 5869
rect 14028 5122 14084 5124
rect 14028 5070 14030 5122
rect 14030 5070 14082 5122
rect 14082 5070 14084 5122
rect 14028 5068 14084 5070
rect 15372 4844 15428 4900
rect 14364 4508 14420 4564
rect 8316 4284 8372 4340
rect 15708 4396 15764 4452
rect 16268 5404 16324 5460
rect 16380 5292 16436 5348
rect 16492 5906 16548 5908
rect 16492 5854 16494 5906
rect 16494 5854 16546 5906
rect 16546 5854 16548 5906
rect 16492 5852 16548 5854
rect 15036 4338 15092 4340
rect 15036 4286 15038 4338
rect 15038 4286 15090 4338
rect 15090 4286 15092 4338
rect 15036 4284 15092 4286
rect 16940 6076 16996 6132
rect 16828 5628 16884 5684
rect 16604 5404 16660 5460
rect 16716 5292 16772 5348
rect 17500 6076 17556 6132
rect 17612 6690 17668 6692
rect 17612 6638 17614 6690
rect 17614 6638 17666 6690
rect 17666 6638 17668 6690
rect 17612 6636 17668 6638
rect 17500 5628 17556 5684
rect 19908 9100 19964 9156
rect 19740 9042 19796 9044
rect 18620 8230 18676 8260
rect 18620 8204 18622 8230
rect 18622 8204 18674 8230
rect 18674 8204 18676 8230
rect 18396 7980 18452 8036
rect 19740 8990 19742 9042
rect 19742 8990 19794 9042
rect 19794 8990 19796 9042
rect 19740 8988 19796 8990
rect 19404 8316 19460 8372
rect 20188 8316 20244 8372
rect 19852 8092 19908 8148
rect 20412 8092 20468 8148
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19404 6748 19460 6804
rect 18116 6578 18172 6580
rect 18116 6526 18118 6578
rect 18118 6526 18170 6578
rect 18170 6526 18172 6578
rect 18116 6524 18172 6526
rect 19740 7420 19796 7476
rect 19628 6690 19684 6692
rect 19628 6638 19630 6690
rect 19630 6638 19682 6690
rect 19682 6638 19684 6690
rect 19628 6636 19684 6638
rect 20300 7586 20356 7588
rect 20300 7534 20302 7586
rect 20302 7534 20354 7586
rect 20354 7534 20356 7586
rect 20300 7532 20356 7534
rect 19852 6636 19908 6692
rect 19068 6300 19124 6356
rect 20300 6690 20356 6692
rect 20300 6638 20302 6690
rect 20302 6638 20354 6690
rect 20354 6638 20356 6690
rect 20300 6636 20356 6638
rect 20524 8034 20580 8036
rect 20524 7982 20526 8034
rect 20526 7982 20578 8034
rect 20578 7982 20580 8034
rect 20524 7980 20580 7982
rect 24780 12684 24836 12740
rect 22876 10610 22932 10612
rect 22876 10558 22878 10610
rect 22878 10558 22930 10610
rect 22930 10558 22932 10610
rect 22876 10556 22932 10558
rect 24668 11676 24724 11732
rect 24174 10780 24230 10836
rect 24332 10668 24388 10724
rect 24444 10610 24500 10612
rect 24444 10558 24446 10610
rect 24446 10558 24498 10610
rect 24498 10558 24500 10610
rect 24444 10556 24500 10558
rect 25900 13522 25956 13524
rect 25900 13470 25902 13522
rect 25902 13470 25954 13522
rect 25954 13470 25956 13522
rect 25900 13468 25956 13470
rect 26572 13356 26628 13412
rect 25900 13244 25956 13300
rect 25788 12178 25844 12180
rect 25788 12126 25790 12178
rect 25790 12126 25842 12178
rect 25842 12126 25844 12178
rect 25788 12124 25844 12126
rect 25340 11564 25396 11620
rect 25452 11506 25508 11508
rect 25452 11454 25454 11506
rect 25454 11454 25506 11506
rect 25506 11454 25508 11506
rect 25452 11452 25508 11454
rect 24780 10780 24836 10836
rect 23100 10220 23156 10276
rect 23660 9938 23716 9940
rect 23660 9886 23662 9938
rect 23662 9886 23714 9938
rect 23714 9886 23716 9938
rect 23660 9884 23716 9886
rect 22316 9436 22372 9492
rect 22876 9436 22932 9492
rect 23324 9436 23380 9492
rect 21924 8482 21980 8484
rect 21924 8430 21926 8482
rect 21926 8430 21978 8482
rect 21978 8430 21980 8482
rect 21924 8428 21980 8430
rect 21588 8258 21644 8260
rect 21588 8206 21590 8258
rect 21590 8206 21642 8258
rect 21642 8206 21644 8258
rect 21588 8204 21644 8206
rect 25340 11340 25396 11396
rect 25452 10610 25508 10612
rect 25452 10558 25454 10610
rect 25454 10558 25506 10610
rect 25506 10558 25508 10610
rect 25452 10556 25508 10558
rect 25676 11452 25732 11508
rect 27916 16210 27972 16212
rect 27916 16158 27918 16210
rect 27918 16158 27970 16210
rect 27970 16158 27972 16210
rect 27916 16156 27972 16158
rect 27804 16044 27860 16100
rect 29988 18732 30044 18788
rect 28924 18338 28980 18340
rect 28924 18286 28926 18338
rect 28926 18286 28978 18338
rect 28978 18286 28980 18338
rect 28924 18284 28980 18286
rect 30772 19852 30828 19908
rect 31052 19964 31108 20020
rect 30828 19628 30884 19684
rect 31276 21644 31332 21700
rect 31276 21474 31332 21476
rect 31276 21422 31278 21474
rect 31278 21422 31330 21474
rect 31330 21422 31332 21474
rect 31276 21420 31332 21422
rect 31388 21308 31444 21364
rect 33404 21756 33460 21812
rect 31612 21586 31668 21588
rect 31612 21534 31614 21586
rect 31614 21534 31666 21586
rect 31666 21534 31668 21586
rect 31612 21532 31668 21534
rect 32956 21532 33012 21588
rect 32396 21420 32452 21476
rect 31276 20018 31332 20020
rect 31276 19966 31278 20018
rect 31278 19966 31330 20018
rect 31330 19966 31332 20018
rect 32060 20748 32116 20804
rect 32564 21084 32620 21140
rect 32060 20188 32116 20244
rect 31948 20018 32004 20020
rect 31276 19964 31332 19966
rect 31948 19966 31950 20018
rect 31950 19966 32002 20018
rect 32002 19966 32004 20018
rect 31948 19964 32004 19966
rect 31612 19906 31668 19908
rect 31612 19854 31614 19906
rect 31614 19854 31666 19906
rect 31666 19854 31668 19906
rect 31612 19852 31668 19854
rect 31388 19628 31444 19684
rect 31164 19234 31220 19236
rect 31164 19182 31166 19234
rect 31166 19182 31218 19234
rect 31218 19182 31220 19234
rect 31164 19180 31220 19182
rect 28588 17500 28644 17556
rect 28924 16882 28980 16884
rect 28924 16830 28926 16882
rect 28926 16830 28978 16882
rect 28978 16830 28980 16882
rect 28924 16828 28980 16830
rect 31052 17612 31108 17668
rect 30156 17052 30212 17108
rect 29260 16828 29316 16884
rect 28252 16044 28308 16100
rect 28700 16098 28756 16100
rect 28700 16046 28702 16098
rect 28702 16046 28754 16098
rect 28754 16046 28756 16098
rect 28700 16044 28756 16046
rect 29484 15596 29540 15652
rect 29260 15484 29316 15540
rect 26796 15036 26852 15092
rect 26796 13244 26852 13300
rect 29372 14530 29428 14532
rect 29372 14478 29374 14530
rect 29374 14478 29426 14530
rect 29426 14478 29428 14530
rect 29372 14476 29428 14478
rect 30044 16828 30100 16884
rect 30380 16940 30436 16996
rect 31164 17164 31220 17220
rect 31388 19180 31444 19236
rect 32452 19404 32508 19460
rect 32956 19628 33012 19684
rect 33068 20300 33124 20356
rect 31948 18425 31950 18452
rect 31950 18425 32002 18452
rect 32002 18425 32004 18452
rect 31948 18396 32004 18425
rect 32284 17836 32340 17892
rect 31948 17666 32004 17668
rect 31948 17614 31950 17666
rect 31950 17614 32002 17666
rect 32002 17614 32004 17666
rect 31948 17612 32004 17614
rect 31612 17052 31668 17108
rect 32844 18396 32900 18452
rect 33236 20130 33292 20132
rect 33236 20078 33238 20130
rect 33238 20078 33290 20130
rect 33290 20078 33292 20130
rect 33236 20076 33292 20078
rect 33908 23154 33964 23156
rect 33908 23102 33910 23154
rect 33910 23102 33962 23154
rect 33962 23102 33964 23154
rect 33908 23100 33964 23102
rect 34076 22428 34132 22484
rect 33740 22316 33796 22372
rect 33740 21756 33796 21812
rect 33852 21532 33908 21588
rect 33628 20972 33684 21028
rect 34580 24332 34636 24388
rect 34580 23884 34636 23940
rect 34916 24668 34972 24724
rect 34748 23772 34804 23828
rect 35588 25506 35644 25508
rect 35588 25454 35590 25506
rect 35590 25454 35642 25506
rect 35642 25454 35644 25506
rect 35588 25452 35644 25454
rect 37324 33740 37380 33796
rect 37660 35586 37716 35588
rect 37660 35534 37662 35586
rect 37662 35534 37714 35586
rect 37714 35534 37716 35586
rect 37660 35532 37716 35534
rect 37884 35308 37940 35364
rect 37660 34914 37716 34916
rect 37660 34862 37662 34914
rect 37662 34862 37714 34914
rect 37714 34862 37716 34914
rect 37660 34860 37716 34862
rect 37772 34748 37828 34804
rect 40460 42364 40516 42420
rect 40684 46620 40740 46676
rect 41468 46674 41524 46676
rect 41468 46622 41470 46674
rect 41470 46622 41522 46674
rect 41522 46622 41524 46674
rect 41468 46620 41524 46622
rect 42364 47346 42420 47348
rect 42364 47294 42366 47346
rect 42366 47294 42418 47346
rect 42418 47294 42420 47346
rect 42364 47292 42420 47294
rect 42980 47292 43036 47348
rect 41804 45890 41860 45892
rect 41804 45838 41806 45890
rect 41806 45838 41858 45890
rect 41858 45838 41860 45890
rect 41804 45836 41860 45838
rect 41356 45724 41412 45780
rect 42140 46620 42196 46676
rect 42140 45612 42196 45668
rect 40908 45106 40964 45108
rect 40908 45054 40910 45106
rect 40910 45054 40962 45106
rect 40962 45054 40964 45106
rect 40908 45052 40964 45054
rect 40684 44492 40740 44548
rect 41784 45106 41840 45108
rect 41784 45054 41786 45106
rect 41786 45054 41838 45106
rect 41838 45054 41840 45106
rect 41784 45052 41840 45054
rect 41244 44604 41300 44660
rect 41244 44322 41300 44324
rect 41244 44270 41246 44322
rect 41246 44270 41298 44322
rect 41298 44270 41300 44322
rect 41244 44268 41300 44270
rect 41468 44434 41524 44436
rect 41468 44382 41470 44434
rect 41470 44382 41522 44434
rect 41522 44382 41524 44434
rect 41468 44380 41524 44382
rect 41804 44492 41860 44548
rect 42364 46508 42420 46564
rect 42364 45388 42420 45444
rect 42700 45890 42756 45892
rect 42700 45838 42702 45890
rect 42702 45838 42754 45890
rect 42754 45838 42756 45890
rect 42700 45836 42756 45838
rect 44492 47516 44548 47572
rect 43820 46844 43876 46900
rect 44268 47180 44324 47236
rect 46396 47570 46452 47572
rect 46396 47518 46398 47570
rect 46398 47518 46450 47570
rect 46450 47518 46452 47570
rect 46396 47516 46452 47518
rect 45724 47292 45780 47348
rect 45276 46844 45332 46900
rect 43576 45612 43632 45668
rect 44044 45500 44100 45556
rect 42476 45164 42532 45220
rect 42364 45052 42420 45108
rect 42700 45106 42756 45108
rect 42700 45054 42702 45106
rect 42702 45054 42754 45106
rect 42754 45054 42756 45106
rect 42700 45052 42756 45054
rect 42140 44380 42196 44436
rect 41692 43596 41748 43652
rect 42924 44492 42980 44548
rect 42812 44380 42868 44436
rect 43148 45164 43204 45220
rect 43596 44940 43652 44996
rect 43484 44546 43540 44548
rect 43484 44494 43486 44546
rect 43486 44494 43538 44546
rect 43538 44494 43540 44546
rect 43484 44492 43540 44494
rect 43260 44268 43316 44324
rect 42700 43596 42756 43652
rect 42252 43314 42308 43316
rect 42252 43262 42254 43314
rect 42254 43262 42306 43314
rect 42306 43262 42308 43314
rect 42252 43260 42308 43262
rect 42924 43820 42980 43876
rect 44492 45276 44548 45332
rect 44380 44322 44436 44324
rect 44380 44270 44382 44322
rect 44382 44270 44434 44322
rect 44434 44270 44436 44322
rect 44380 44268 44436 44270
rect 43932 44044 43988 44100
rect 43372 43260 43428 43316
rect 40908 42476 40964 42532
rect 41580 41916 41636 41972
rect 41784 42028 41840 42084
rect 43036 43036 43092 43092
rect 42868 42700 42924 42756
rect 42868 42140 42924 42196
rect 42868 41970 42924 41972
rect 42868 41918 42870 41970
rect 42870 41918 42922 41970
rect 42922 41918 42924 41970
rect 42868 41916 42924 41918
rect 43708 42924 43764 42980
rect 44380 43820 44436 43876
rect 43540 42812 43596 42868
rect 43820 42754 43876 42756
rect 43820 42702 43822 42754
rect 43822 42702 43874 42754
rect 43874 42702 43876 42754
rect 43820 42700 43876 42702
rect 43484 42140 43540 42196
rect 44156 43538 44212 43540
rect 44156 43486 44158 43538
rect 44158 43486 44210 43538
rect 44210 43486 44212 43538
rect 44156 43484 44212 43486
rect 44100 42978 44156 42980
rect 44100 42926 44102 42978
rect 44102 42926 44154 42978
rect 44154 42926 44156 42978
rect 44100 42924 44156 42926
rect 44716 45388 44772 45444
rect 44828 44044 44884 44100
rect 45276 45276 45332 45332
rect 45500 45836 45556 45892
rect 45500 44492 45556 44548
rect 46508 47180 46564 47236
rect 45836 46956 45892 47012
rect 49308 47628 49364 47684
rect 47628 47234 47684 47236
rect 47628 47182 47630 47234
rect 47630 47182 47682 47234
rect 47682 47182 47684 47234
rect 47628 47180 47684 47182
rect 46060 46620 46116 46676
rect 45948 45890 46004 45892
rect 45948 45838 45950 45890
rect 45950 45838 46002 45890
rect 46002 45838 46004 45890
rect 45948 45836 46004 45838
rect 46172 46562 46228 46564
rect 46172 46510 46174 46562
rect 46174 46510 46226 46562
rect 46226 46510 46228 46562
rect 46172 46508 46228 46510
rect 46284 46396 46340 46452
rect 46172 45724 46228 45780
rect 45724 45089 45726 45108
rect 45726 45089 45778 45108
rect 45778 45089 45780 45108
rect 45724 45052 45780 45089
rect 46060 44940 46116 44996
rect 45388 44156 45444 44212
rect 44940 43932 44996 43988
rect 45052 43820 45108 43876
rect 44716 43036 44772 43092
rect 43820 41970 43876 41972
rect 43820 41918 43822 41970
rect 43822 41918 43874 41970
rect 43874 41918 43876 41970
rect 43820 41916 43876 41918
rect 44268 41916 44324 41972
rect 44492 41244 44548 41300
rect 40572 40908 40628 40964
rect 41076 40962 41132 40964
rect 41076 40910 41078 40962
rect 41078 40910 41130 40962
rect 41130 40910 41132 40962
rect 41076 40908 41132 40910
rect 40460 40460 40516 40516
rect 40796 40348 40852 40404
rect 40460 38556 40516 38612
rect 40684 39340 40740 39396
rect 40348 37772 40404 37828
rect 40572 37996 40628 38052
rect 39116 37378 39172 37380
rect 39116 37326 39118 37378
rect 39118 37326 39170 37378
rect 39170 37326 39172 37378
rect 39116 37324 39172 37326
rect 40404 37378 40460 37380
rect 40404 37326 40406 37378
rect 40406 37326 40458 37378
rect 40458 37326 40460 37378
rect 40404 37324 40460 37326
rect 38556 36876 38612 36932
rect 39732 36876 39788 36932
rect 40236 36988 40292 37044
rect 38220 35308 38276 35364
rect 37884 34524 37940 34580
rect 37996 34636 38052 34692
rect 37996 34242 38052 34244
rect 37996 34190 37998 34242
rect 37998 34190 38050 34242
rect 38050 34190 38052 34242
rect 37996 34188 38052 34190
rect 37212 32620 37268 32676
rect 38108 32732 38164 32788
rect 38220 32396 38276 32452
rect 38108 32172 38164 32228
rect 36876 30268 36932 30324
rect 35868 29372 35924 29428
rect 35980 29596 36036 29652
rect 36876 29372 36932 29428
rect 35868 28700 35924 28756
rect 36036 28812 36092 28868
rect 36876 28812 36932 28868
rect 36484 28642 36540 28644
rect 36484 28590 36486 28642
rect 36486 28590 36538 28642
rect 36538 28590 36540 28642
rect 36484 28588 36540 28590
rect 36876 28476 36932 28532
rect 36988 29484 37044 29540
rect 36764 28364 36820 28420
rect 36148 28082 36204 28084
rect 36148 28030 36150 28082
rect 36150 28030 36202 28082
rect 36202 28030 36204 28082
rect 36148 28028 36204 28030
rect 35868 26850 35924 26852
rect 35868 26798 35870 26850
rect 35870 26798 35922 26850
rect 35922 26798 35924 26850
rect 35868 26796 35924 26798
rect 35868 25506 35924 25508
rect 35868 25454 35870 25506
rect 35870 25454 35922 25506
rect 35922 25454 35924 25506
rect 35868 25452 35924 25454
rect 35756 25116 35812 25172
rect 35196 24330 35252 24332
rect 34972 24220 35028 24276
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 34860 23660 34916 23716
rect 34916 23436 34972 23492
rect 34468 23378 34524 23380
rect 34468 23326 34470 23378
rect 34470 23326 34522 23378
rect 34522 23326 34524 23378
rect 34468 23324 34524 23326
rect 35420 23938 35476 23940
rect 35420 23886 35422 23938
rect 35422 23886 35474 23938
rect 35474 23886 35476 23938
rect 35420 23884 35476 23886
rect 35308 23436 35364 23492
rect 34636 22428 34692 22484
rect 34300 22204 34356 22260
rect 34860 22342 34916 22372
rect 34860 22316 34862 22342
rect 34862 22316 34914 22342
rect 34914 22316 34916 22342
rect 35084 23324 35140 23380
rect 35308 23042 35364 23044
rect 35308 22990 35310 23042
rect 35310 22990 35362 23042
rect 35362 22990 35364 23042
rect 35308 22988 35364 22990
rect 35420 22876 35476 22932
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35420 22342 35476 22372
rect 35420 22316 35422 22342
rect 35422 22316 35474 22342
rect 35474 22316 35476 22342
rect 34972 21868 35028 21924
rect 34412 21756 34468 21812
rect 35308 21308 35364 21364
rect 34188 21084 34244 21140
rect 34300 21196 34356 21252
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 34860 20972 34916 21028
rect 34356 20188 34412 20244
rect 33852 20076 33908 20132
rect 35868 22988 35924 23044
rect 35644 22428 35700 22484
rect 35868 21308 35924 21364
rect 35532 20972 35588 21028
rect 35196 20524 35252 20580
rect 34748 20076 34804 20132
rect 35140 20018 35196 20020
rect 35140 19966 35142 20018
rect 35142 19966 35194 20018
rect 35194 19966 35196 20018
rect 35140 19964 35196 19966
rect 34860 19740 34916 19796
rect 34636 19516 34692 19572
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 33628 18426 33630 18452
rect 33630 18426 33682 18452
rect 33682 18426 33684 18452
rect 33628 18396 33684 18426
rect 33908 18620 33964 18676
rect 35756 19346 35812 19348
rect 35756 19294 35758 19346
rect 35758 19294 35810 19346
rect 35810 19294 35812 19346
rect 35756 19292 35812 19294
rect 35532 18620 35588 18676
rect 37212 28642 37268 28644
rect 37212 28590 37214 28642
rect 37214 28590 37266 28642
rect 37266 28590 37268 28642
rect 37212 28588 37268 28590
rect 37436 30182 37492 30212
rect 37436 30156 37438 30182
rect 37438 30156 37490 30182
rect 37490 30156 37492 30182
rect 37660 30044 37716 30100
rect 37996 30716 38052 30772
rect 37884 30268 37940 30324
rect 37548 28642 37604 28644
rect 37548 28590 37550 28642
rect 37550 28590 37602 28642
rect 37602 28590 37604 28642
rect 37548 28588 37604 28590
rect 37436 28028 37492 28084
rect 37268 27634 37324 27636
rect 37268 27582 37270 27634
rect 37270 27582 37322 27634
rect 37322 27582 37324 27634
rect 37268 27580 37324 27582
rect 36484 26962 36540 26964
rect 36484 26910 36486 26962
rect 36486 26910 36538 26962
rect 36538 26910 36540 26962
rect 36484 26908 36540 26910
rect 37436 27244 37492 27300
rect 37324 27132 37380 27188
rect 36988 27020 37044 27076
rect 37772 29148 37828 29204
rect 37884 28754 37940 28756
rect 37884 28702 37886 28754
rect 37886 28702 37938 28754
rect 37938 28702 37940 28754
rect 37884 28700 37940 28702
rect 37772 27804 37828 27860
rect 37884 28028 37940 28084
rect 39340 36204 39396 36260
rect 39620 35922 39676 35924
rect 39620 35870 39622 35922
rect 39622 35870 39674 35922
rect 39674 35870 39676 35922
rect 39620 35868 39676 35870
rect 38892 35474 38948 35476
rect 38892 35422 38894 35474
rect 38894 35422 38946 35474
rect 38946 35422 38948 35474
rect 38892 35420 38948 35422
rect 38444 34860 38500 34916
rect 38892 34748 38948 34804
rect 40348 35868 40404 35924
rect 41692 40908 41748 40964
rect 42364 40908 42420 40964
rect 41524 40684 41580 40740
rect 41356 40402 41412 40404
rect 41356 40350 41358 40402
rect 41358 40350 41410 40402
rect 41410 40350 41412 40402
rect 41356 40348 41412 40350
rect 41804 40460 41860 40516
rect 42924 40460 42980 40516
rect 42588 40402 42644 40404
rect 42588 40350 42590 40402
rect 42590 40350 42642 40402
rect 42642 40350 42644 40402
rect 42588 40348 42644 40350
rect 41244 39340 41300 39396
rect 41636 39228 41692 39284
rect 41244 38050 41300 38052
rect 41244 37998 41246 38050
rect 41246 37998 41298 38050
rect 41298 37998 41300 38050
rect 41244 37996 41300 37998
rect 41580 38035 41636 38052
rect 41580 37996 41582 38035
rect 41582 37996 41634 38035
rect 41634 37996 41636 38035
rect 40796 37212 40852 37268
rect 41020 37436 41076 37492
rect 41356 37436 41412 37492
rect 40684 37100 40740 37156
rect 39060 34188 39116 34244
rect 38556 33628 38612 33684
rect 39004 32844 39060 32900
rect 38668 32620 38724 32676
rect 38444 30268 38500 30324
rect 38780 31948 38836 32004
rect 38332 29820 38388 29876
rect 38220 28642 38276 28644
rect 38220 28590 38222 28642
rect 38222 28590 38274 28642
rect 38274 28590 38276 28642
rect 38220 28588 38276 28590
rect 39004 31836 39060 31892
rect 38780 31164 38836 31220
rect 40236 35420 40292 35476
rect 41244 36988 41300 37044
rect 41020 36204 41076 36260
rect 40572 35980 40628 36036
rect 41580 35868 41636 35924
rect 41468 35756 41524 35812
rect 42532 39676 42588 39732
rect 42532 39394 42588 39396
rect 42532 39342 42534 39394
rect 42534 39342 42586 39394
rect 42586 39342 42588 39394
rect 44380 41020 44436 41076
rect 43876 40962 43932 40964
rect 43876 40910 43878 40962
rect 43878 40910 43930 40962
rect 43930 40910 43932 40962
rect 43876 40908 43932 40910
rect 44212 40460 44268 40516
rect 43372 40348 43428 40404
rect 42532 39340 42588 39342
rect 43260 39116 43316 39172
rect 42084 39004 42140 39060
rect 44492 40378 44494 40404
rect 44494 40378 44546 40404
rect 44546 40378 44548 40404
rect 44492 40348 44548 40378
rect 45164 43596 45220 43652
rect 45164 41970 45220 41972
rect 45164 41918 45166 41970
rect 45166 41918 45218 41970
rect 45218 41918 45220 41970
rect 45164 41916 45220 41918
rect 45388 42812 45444 42868
rect 44940 41468 44996 41524
rect 45052 40460 45108 40516
rect 43484 39788 43540 39844
rect 44492 39676 44548 39732
rect 42495 38108 42551 38164
rect 42252 38050 42308 38052
rect 42252 37998 42254 38050
rect 42254 37998 42306 38050
rect 42306 37998 42308 38050
rect 42252 37996 42308 37998
rect 43708 38162 43764 38164
rect 43708 38110 43710 38162
rect 43710 38110 43762 38162
rect 43762 38110 43764 38162
rect 43708 38108 43764 38110
rect 44156 39116 44212 39172
rect 43820 37772 43876 37828
rect 44044 38220 44100 38276
rect 44268 38108 44324 38164
rect 44156 38050 44212 38052
rect 44156 37998 44158 38050
rect 44158 37998 44210 38050
rect 44210 37998 44212 38050
rect 44156 37996 44212 37998
rect 44044 37884 44100 37940
rect 41804 37324 41860 37380
rect 42364 37266 42420 37268
rect 42364 37214 42366 37266
rect 42366 37214 42418 37266
rect 42418 37214 42420 37266
rect 42364 37212 42420 37214
rect 42364 35922 42420 35924
rect 42364 35870 42366 35922
rect 42366 35870 42418 35922
rect 42418 35870 42420 35922
rect 42364 35868 42420 35870
rect 43820 36467 43876 36484
rect 43820 36428 43822 36467
rect 43822 36428 43874 36467
rect 43874 36428 43876 36467
rect 44268 37324 44324 37380
rect 44604 39340 44660 39396
rect 44492 38780 44548 38836
rect 44604 38444 44660 38500
rect 45276 40378 45278 40404
rect 45278 40378 45330 40404
rect 45330 40378 45332 40404
rect 45276 40348 45332 40378
rect 45500 41468 45556 41524
rect 45500 41298 45556 41300
rect 45500 41246 45502 41298
rect 45502 41246 45554 41298
rect 45554 41246 45556 41298
rect 45500 41244 45556 41246
rect 48076 46396 48132 46452
rect 46172 44380 46228 44436
rect 46060 44156 46116 44212
rect 46396 44492 46452 44548
rect 46508 44380 46564 44436
rect 46508 43820 46564 43876
rect 47180 45500 47236 45556
rect 47292 45276 47348 45332
rect 46732 44716 46788 44772
rect 45948 43538 46004 43540
rect 45948 43486 45950 43538
rect 45950 43486 46002 43538
rect 46002 43486 46004 43538
rect 45948 43484 46004 43486
rect 45724 41186 45780 41188
rect 45724 41134 45726 41186
rect 45726 41134 45778 41186
rect 45778 41134 45780 41186
rect 45724 41132 45780 41134
rect 45948 41020 46004 41076
rect 46396 41916 46452 41972
rect 47180 45052 47236 45108
rect 46844 44604 46900 44660
rect 47404 45052 47460 45108
rect 46844 44156 46900 44212
rect 46732 43484 46788 43540
rect 46452 41132 46508 41188
rect 46620 41074 46676 41076
rect 46620 41022 46622 41074
rect 46622 41022 46674 41074
rect 46674 41022 46676 41074
rect 46620 41020 46676 41022
rect 46284 40402 46340 40404
rect 46284 40350 46286 40402
rect 46286 40350 46338 40402
rect 46338 40350 46340 40402
rect 46284 40348 46340 40350
rect 45612 39788 45668 39844
rect 44884 39116 44940 39172
rect 44828 38834 44884 38836
rect 44828 38782 44830 38834
rect 44830 38782 44882 38834
rect 44882 38782 44884 38834
rect 44828 38780 44884 38782
rect 45500 39564 45556 39620
rect 46004 39788 46060 39844
rect 46396 39730 46452 39732
rect 46396 39678 46398 39730
rect 46398 39678 46450 39730
rect 46450 39678 46452 39730
rect 46396 39676 46452 39678
rect 45948 39618 46004 39620
rect 45948 39566 45950 39618
rect 45950 39566 46002 39618
rect 46002 39566 46004 39618
rect 45948 39564 46004 39566
rect 45836 38892 45892 38948
rect 45276 38834 45332 38836
rect 45276 38782 45278 38834
rect 45278 38782 45330 38834
rect 45330 38782 45332 38834
rect 45276 38780 45332 38782
rect 44716 38332 44772 38388
rect 45276 38444 45332 38500
rect 44492 37996 44548 38052
rect 44940 38050 44996 38052
rect 44940 37998 44942 38050
rect 44942 37998 44994 38050
rect 44994 37998 44996 38050
rect 44940 37996 44996 37998
rect 44940 37266 44996 37268
rect 44940 37214 44942 37266
rect 44942 37214 44994 37266
rect 44994 37214 44996 37266
rect 44940 37212 44996 37214
rect 44380 36876 44436 36932
rect 44044 36204 44100 36260
rect 41244 35420 41300 35476
rect 40572 35308 40628 35364
rect 40460 35196 40516 35252
rect 39900 34300 39956 34356
rect 40684 34914 40740 34916
rect 40684 34862 40686 34914
rect 40686 34862 40738 34914
rect 40738 34862 40740 34914
rect 40684 34860 40740 34862
rect 40236 33964 40292 34020
rect 39900 33740 39956 33796
rect 39340 33292 39396 33348
rect 39452 33180 39508 33236
rect 39452 32732 39508 32788
rect 39452 31948 39508 32004
rect 40012 33122 40068 33124
rect 40012 33070 40014 33122
rect 40014 33070 40066 33122
rect 40066 33070 40068 33122
rect 40012 33068 40068 33070
rect 40012 32732 40068 32788
rect 39676 32172 39732 32228
rect 39564 31836 39620 31892
rect 39228 31052 39284 31108
rect 38668 30210 38724 30212
rect 38668 30158 38670 30210
rect 38670 30158 38722 30210
rect 38722 30158 38724 30210
rect 38668 30156 38724 30158
rect 39004 30828 39060 30884
rect 38892 30156 38948 30212
rect 38556 29596 38612 29652
rect 38892 29932 38948 29988
rect 38556 29426 38612 29428
rect 38556 29374 38558 29426
rect 38558 29374 38610 29426
rect 38610 29374 38612 29426
rect 38556 29372 38612 29374
rect 38332 28364 38388 28420
rect 38332 28028 38388 28084
rect 38108 27580 38164 27636
rect 37660 27020 37716 27076
rect 36988 26684 37044 26740
rect 36204 24892 36260 24948
rect 36372 23436 36428 23492
rect 37212 26796 37268 26852
rect 37212 24892 37268 24948
rect 37100 24162 37156 24164
rect 37100 24110 37102 24162
rect 37102 24110 37154 24162
rect 37154 24110 37156 24162
rect 37100 24108 37156 24110
rect 36988 23324 37044 23380
rect 37604 26684 37660 26740
rect 37436 26460 37492 26516
rect 38444 27858 38500 27860
rect 38444 27806 38446 27858
rect 38446 27806 38498 27858
rect 38498 27806 38500 27858
rect 38444 27804 38500 27806
rect 38220 27244 38276 27300
rect 37772 26236 37828 26292
rect 37884 27132 37940 27188
rect 38108 27132 38164 27188
rect 37772 25506 37828 25508
rect 37772 25454 37774 25506
rect 37774 25454 37826 25506
rect 37826 25454 37828 25506
rect 37772 25452 37828 25454
rect 37772 25228 37828 25284
rect 37324 23100 37380 23156
rect 36988 22988 37044 23044
rect 37436 22988 37492 23044
rect 37324 22876 37380 22932
rect 36988 21980 37044 22036
rect 37996 27020 38052 27076
rect 38780 29260 38836 29316
rect 39228 30210 39284 30212
rect 39228 30158 39230 30210
rect 39230 30158 39282 30210
rect 39282 30158 39284 30210
rect 39228 30156 39284 30158
rect 40012 31052 40068 31108
rect 39900 30156 39956 30212
rect 39116 30044 39172 30100
rect 41804 35420 41860 35476
rect 41580 35308 41636 35364
rect 41468 34972 41524 35028
rect 41692 34972 41748 35028
rect 41468 34188 41524 34244
rect 41580 34130 41636 34132
rect 41580 34078 41582 34130
rect 41582 34078 41634 34130
rect 41634 34078 41636 34130
rect 41580 34076 41636 34078
rect 40908 33307 40964 33348
rect 40908 33292 40910 33307
rect 40910 33292 40962 33307
rect 40962 33292 40964 33307
rect 40292 32562 40348 32564
rect 40292 32510 40294 32562
rect 40294 32510 40346 32562
rect 40346 32510 40348 32562
rect 40292 32508 40348 32510
rect 40796 32562 40852 32564
rect 40796 32510 40798 32562
rect 40798 32510 40850 32562
rect 40850 32510 40852 32562
rect 40796 32508 40852 32510
rect 44156 35308 44212 35364
rect 43596 35196 43652 35252
rect 42140 34972 42196 35028
rect 42028 34748 42084 34804
rect 41916 34188 41972 34244
rect 43260 34972 43316 35028
rect 42588 34914 42644 34916
rect 42588 34862 42590 34914
rect 42590 34862 42642 34914
rect 42642 34862 42644 34914
rect 42588 34860 42644 34862
rect 42756 34748 42812 34804
rect 42028 34076 42084 34132
rect 41972 33628 42028 33684
rect 41804 32844 41860 32900
rect 42028 32732 42084 32788
rect 41468 32508 41524 32564
rect 40908 30977 40910 30996
rect 40910 30977 40962 30996
rect 40962 30977 40964 30996
rect 40908 30940 40964 30977
rect 41244 30970 41246 30996
rect 41246 30970 41298 30996
rect 41298 30970 41300 30996
rect 41244 30940 41300 30970
rect 44940 36428 44996 36484
rect 42924 34130 42980 34132
rect 42924 34078 42926 34130
rect 42926 34078 42978 34130
rect 42978 34078 42980 34130
rect 42924 34076 42980 34078
rect 42588 33628 42644 33684
rect 43652 34130 43708 34132
rect 43652 34078 43654 34130
rect 43654 34078 43706 34130
rect 43706 34078 43708 34130
rect 43652 34076 43708 34078
rect 42924 33628 42980 33684
rect 43148 33404 43204 33460
rect 43820 33404 43876 33460
rect 42924 33180 42980 33236
rect 43876 33180 43932 33236
rect 42476 32732 42532 32788
rect 44492 33068 44548 33124
rect 42812 32562 42868 32564
rect 42812 32510 42814 32562
rect 42814 32510 42866 32562
rect 42866 32510 42868 32562
rect 42812 32508 42868 32510
rect 43372 32450 43428 32452
rect 43372 32398 43374 32450
rect 43374 32398 43426 32450
rect 43426 32398 43428 32450
rect 43372 32396 43428 32398
rect 42028 31948 42084 32004
rect 42588 31948 42644 32004
rect 41020 30828 41076 30884
rect 40124 30044 40180 30100
rect 41356 30156 41412 30212
rect 39284 29202 39340 29204
rect 39284 29150 39286 29202
rect 39286 29150 39338 29202
rect 39338 29150 39340 29202
rect 39284 29148 39340 29150
rect 41076 29426 41132 29428
rect 41076 29374 41078 29426
rect 41078 29374 41130 29426
rect 41130 29374 41132 29426
rect 41076 29372 41132 29374
rect 39452 29148 39508 29204
rect 41020 29148 41076 29204
rect 39004 28924 39060 28980
rect 38892 28642 38948 28644
rect 38892 28590 38894 28642
rect 38894 28590 38946 28642
rect 38946 28590 38948 28642
rect 38892 28588 38948 28590
rect 40796 28642 40852 28644
rect 40796 28590 40798 28642
rect 40798 28590 40850 28642
rect 40850 28590 40852 28642
rect 40796 28588 40852 28590
rect 39004 28252 39060 28308
rect 40236 28364 40292 28420
rect 42252 31106 42308 31108
rect 42252 31054 42254 31106
rect 42254 31054 42306 31106
rect 42306 31054 42308 31106
rect 42252 31052 42308 31054
rect 41468 29596 41524 29652
rect 41076 28082 41132 28084
rect 41076 28030 41078 28082
rect 41078 28030 41130 28082
rect 41130 28030 41132 28082
rect 41076 28028 41132 28030
rect 39150 27916 39206 27972
rect 39004 27858 39060 27860
rect 39004 27806 39006 27858
rect 39006 27806 39058 27858
rect 39058 27806 39060 27858
rect 39004 27804 39060 27806
rect 38780 27132 38836 27188
rect 41356 27858 41412 27860
rect 41356 27806 41358 27858
rect 41358 27806 41410 27858
rect 41410 27806 41412 27858
rect 41356 27804 41412 27806
rect 40796 27186 40852 27188
rect 40796 27134 40798 27186
rect 40798 27134 40850 27186
rect 40850 27134 40852 27186
rect 40796 27132 40852 27134
rect 39004 26908 39060 26964
rect 41132 27074 41188 27076
rect 41132 27022 41134 27074
rect 41134 27022 41186 27074
rect 41186 27022 41188 27074
rect 41132 27020 41188 27022
rect 42028 29596 42084 29652
rect 41916 28812 41972 28868
rect 41916 27186 41972 27188
rect 41916 27134 41918 27186
rect 41918 27134 41970 27186
rect 41970 27134 41972 27186
rect 41916 27132 41972 27134
rect 38108 26572 38164 26628
rect 38780 26460 38836 26516
rect 39340 26460 39396 26516
rect 39116 26348 39172 26404
rect 39452 26266 39454 26292
rect 39454 26266 39506 26292
rect 39506 26266 39508 26292
rect 39452 26236 39508 26266
rect 38108 25228 38164 25284
rect 38948 25730 39004 25732
rect 38948 25678 38950 25730
rect 38950 25678 39002 25730
rect 39002 25678 39004 25730
rect 38948 25676 39004 25678
rect 38668 25478 38724 25508
rect 38668 25452 38670 25478
rect 38670 25452 38722 25478
rect 38722 25452 38724 25478
rect 38332 25228 38388 25284
rect 38220 24722 38276 24724
rect 38220 24670 38222 24722
rect 38222 24670 38274 24722
rect 38274 24670 38276 24722
rect 38220 24668 38276 24670
rect 38780 25116 38836 25172
rect 39900 26348 39956 26404
rect 39564 25676 39620 25732
rect 38556 24108 38612 24164
rect 38444 23996 38500 24052
rect 37996 23884 38052 23940
rect 38332 23772 38388 23828
rect 38220 22988 38276 23044
rect 38444 23100 38500 23156
rect 37548 22204 37604 22260
rect 37212 21868 37268 21924
rect 36092 21586 36148 21588
rect 36092 21534 36094 21586
rect 36094 21534 36146 21586
rect 36146 21534 36148 21586
rect 36092 21532 36148 21534
rect 36092 21308 36148 21364
rect 36428 21532 36484 21588
rect 37436 21532 37492 21588
rect 36372 20578 36428 20580
rect 36372 20526 36374 20578
rect 36374 20526 36426 20578
rect 36426 20526 36428 20578
rect 36372 20524 36428 20526
rect 36204 20188 36260 20244
rect 35980 18732 36036 18788
rect 35868 18620 35924 18676
rect 34524 18450 34580 18452
rect 34524 18398 34526 18450
rect 34526 18398 34578 18450
rect 34578 18398 34580 18450
rect 34524 18396 34580 18398
rect 33740 17724 33796 17780
rect 33404 17612 33460 17668
rect 31276 16940 31332 16996
rect 31948 16940 32004 16996
rect 30784 16268 30840 16324
rect 30940 16098 30996 16100
rect 30940 16046 30942 16098
rect 30942 16046 30994 16098
rect 30994 16046 30996 16098
rect 30940 16044 30996 16046
rect 30604 15596 30660 15652
rect 30492 15484 30548 15540
rect 29932 14700 29988 14756
rect 27468 13244 27524 13300
rect 28364 13244 28420 13300
rect 26684 13020 26740 13076
rect 28252 12962 28308 12964
rect 28252 12910 28254 12962
rect 28254 12910 28306 12962
rect 28306 12910 28308 12962
rect 28252 12908 28308 12910
rect 29484 13244 29540 13300
rect 29260 12908 29316 12964
rect 28364 12684 28420 12740
rect 27580 12290 27636 12292
rect 27580 12238 27582 12290
rect 27582 12238 27634 12290
rect 27634 12238 27636 12290
rect 27580 12236 27636 12238
rect 26292 11954 26348 11956
rect 26292 11902 26294 11954
rect 26294 11902 26346 11954
rect 26346 11902 26348 11954
rect 26292 11900 26348 11902
rect 26124 11452 26180 11508
rect 26684 12124 26740 12180
rect 24108 8876 24164 8932
rect 25116 8876 25172 8932
rect 23324 8482 23380 8484
rect 23324 8430 23326 8482
rect 23326 8430 23378 8482
rect 23378 8430 23380 8482
rect 23324 8428 23380 8430
rect 22316 8230 22372 8260
rect 22316 8204 22318 8230
rect 22318 8204 22370 8230
rect 22370 8204 22372 8230
rect 20636 7420 20692 7476
rect 20860 8092 20916 8148
rect 21084 7532 21140 7588
rect 21756 7474 21812 7476
rect 21756 7422 21758 7474
rect 21758 7422 21810 7474
rect 21810 7422 21812 7474
rect 21756 7420 21812 7422
rect 20748 6748 20804 6804
rect 20412 6524 20468 6580
rect 18340 6130 18396 6132
rect 18340 6078 18342 6130
rect 18342 6078 18394 6130
rect 18394 6078 18396 6130
rect 18340 6076 18396 6078
rect 19068 5906 19124 5908
rect 19068 5854 19070 5906
rect 19070 5854 19122 5906
rect 19122 5854 19124 5906
rect 19404 5964 19460 6020
rect 19068 5852 19124 5854
rect 17836 5628 17892 5684
rect 19068 5628 19124 5684
rect 17500 5180 17556 5236
rect 16940 5068 16996 5124
rect 16492 4172 16548 4228
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 14700 3612 14756 3668
rect 17276 5068 17332 5124
rect 1148 3388 1204 3444
rect 1764 3388 1820 3444
rect 4732 3388 4788 3444
rect 5572 3388 5628 3444
rect 18508 5068 18564 5124
rect 18956 5068 19012 5124
rect 18732 4956 18788 5012
rect 17724 4844 17780 4900
rect 17444 4226 17500 4228
rect 17444 4174 17446 4226
rect 17446 4174 17498 4226
rect 17498 4174 17500 4226
rect 17444 4172 17500 4174
rect 17724 3666 17780 3668
rect 17724 3614 17726 3666
rect 17726 3614 17778 3666
rect 17778 3614 17780 3666
rect 17724 3612 17780 3614
rect 18508 4284 18564 4340
rect 18396 4172 18452 4228
rect 17948 3612 18004 3668
rect 19404 5068 19460 5124
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 20076 6076 20132 6132
rect 20300 5682 20356 5684
rect 20300 5630 20302 5682
rect 20302 5630 20354 5682
rect 20354 5630 20356 5682
rect 20300 5628 20356 5630
rect 20188 5180 20244 5236
rect 20636 5180 20692 5236
rect 20188 4844 20244 4900
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 19628 3666 19684 3668
rect 19628 3614 19630 3666
rect 19630 3614 19682 3666
rect 19682 3614 19684 3666
rect 19628 3612 19684 3614
rect 20748 5068 20804 5124
rect 21196 6412 21252 6468
rect 21532 6466 21588 6468
rect 21532 6414 21534 6466
rect 21534 6414 21586 6466
rect 21586 6414 21588 6466
rect 21532 6412 21588 6414
rect 22186 5906 22242 5908
rect 22186 5854 22188 5906
rect 22188 5854 22240 5906
rect 22240 5854 22242 5906
rect 22186 5852 22242 5854
rect 22186 4508 22242 4564
rect 20300 3612 20356 3668
rect 20860 3612 20916 3668
rect 20132 3388 20188 3444
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 22092 3666 22148 3668
rect 22092 3614 22094 3666
rect 22094 3614 22146 3666
rect 22146 3614 22148 3666
rect 22092 3612 22148 3614
rect 23436 6690 23492 6692
rect 23436 6638 23438 6690
rect 23438 6638 23490 6690
rect 23490 6638 23492 6690
rect 23436 6636 23492 6638
rect 22932 6412 22988 6468
rect 24332 8764 24388 8820
rect 23996 8092 24052 8148
rect 23884 6636 23940 6692
rect 25452 8818 25508 8820
rect 25452 8766 25454 8818
rect 25454 8766 25506 8818
rect 25506 8766 25508 8818
rect 25452 8764 25508 8766
rect 25116 8428 25172 8484
rect 23772 5964 23828 6020
rect 24332 6663 24388 6692
rect 24332 6636 24334 6663
rect 24334 6636 24386 6663
rect 24386 6636 24388 6663
rect 25452 8428 25508 8484
rect 25508 8146 25564 8148
rect 25508 8094 25510 8146
rect 25510 8094 25562 8146
rect 25562 8094 25564 8146
rect 25508 8092 25564 8094
rect 26572 10780 26628 10836
rect 26348 10610 26404 10612
rect 26348 10558 26350 10610
rect 26350 10558 26402 10610
rect 26402 10558 26404 10610
rect 26348 10556 26404 10558
rect 26516 10444 26572 10500
rect 27244 12178 27300 12180
rect 27244 12126 27246 12178
rect 27246 12126 27298 12178
rect 27298 12126 27300 12178
rect 27244 12124 27300 12126
rect 28812 12684 28868 12740
rect 28476 11452 28532 11508
rect 27804 10834 27860 10836
rect 27804 10782 27806 10834
rect 27806 10782 27858 10834
rect 27858 10782 27860 10834
rect 27804 10780 27860 10782
rect 28140 10610 28196 10612
rect 28140 10558 28142 10610
rect 28142 10558 28194 10610
rect 28194 10558 28196 10610
rect 28140 10556 28196 10558
rect 29372 12684 29428 12740
rect 29148 12348 29204 12404
rect 29932 13468 29988 13524
rect 30044 14476 30100 14532
rect 29596 12908 29652 12964
rect 29708 13020 29764 13076
rect 30492 13468 30548 13524
rect 30380 13074 30436 13076
rect 30380 13022 30382 13074
rect 30382 13022 30434 13074
rect 30434 13022 30436 13074
rect 30380 13020 30436 13022
rect 31724 15596 31780 15652
rect 30884 14754 30940 14756
rect 30884 14702 30886 14754
rect 30886 14702 30938 14754
rect 30938 14702 30940 14754
rect 30884 14700 30940 14702
rect 31052 14476 31108 14532
rect 31836 14812 31892 14868
rect 31948 15260 32004 15316
rect 31724 14588 31780 14644
rect 31388 14476 31444 14532
rect 31052 13244 31108 13300
rect 30716 12962 30772 12964
rect 30716 12910 30718 12962
rect 30718 12910 30770 12962
rect 30770 12910 30772 12962
rect 30716 12908 30772 12910
rect 30044 12236 30100 12292
rect 26684 8876 26740 8932
rect 27132 8428 27188 8484
rect 26964 8258 27020 8260
rect 26964 8206 26966 8258
rect 26966 8206 27018 8258
rect 27018 8206 27020 8258
rect 26964 8204 27020 8206
rect 25340 6748 25396 6804
rect 25452 6636 25508 6692
rect 25396 6412 25452 6468
rect 24556 6076 24612 6132
rect 26460 6748 26516 6804
rect 26796 6663 26852 6692
rect 26796 6636 26798 6663
rect 26798 6636 26850 6663
rect 26850 6636 26852 6663
rect 28028 8988 28084 9044
rect 28028 8428 28084 8484
rect 28252 9811 28308 9828
rect 28252 9772 28254 9811
rect 28254 9772 28306 9811
rect 28306 9772 28308 9811
rect 29260 10556 29316 10612
rect 29596 11452 29652 11508
rect 29148 9772 29204 9828
rect 28924 8876 28980 8932
rect 27468 7420 27524 7476
rect 27468 6636 27524 6692
rect 28364 7474 28420 7476
rect 28364 7422 28366 7474
rect 28366 7422 28418 7474
rect 28418 7422 28420 7474
rect 28364 7420 28420 7422
rect 31052 12124 31108 12180
rect 30828 11340 30884 11396
rect 30940 11452 30996 11508
rect 31164 11228 31220 11284
rect 31724 13468 31780 13524
rect 31500 12908 31556 12964
rect 31948 13468 32004 13524
rect 31948 12684 32004 12740
rect 32620 14812 32676 14868
rect 32284 14530 32340 14532
rect 32284 14478 32286 14530
rect 32286 14478 32338 14530
rect 32338 14478 32340 14530
rect 32284 14476 32340 14478
rect 32620 13746 32676 13748
rect 32620 13694 32622 13746
rect 32622 13694 32674 13746
rect 32674 13694 32676 13746
rect 32620 13692 32676 13694
rect 32284 13522 32340 13524
rect 32284 13470 32286 13522
rect 32286 13470 32338 13522
rect 32338 13470 32340 13522
rect 32284 13468 32340 13470
rect 32060 12348 32116 12404
rect 33236 16994 33292 16996
rect 33236 16942 33238 16994
rect 33238 16942 33290 16994
rect 33290 16942 33292 16994
rect 33236 16940 33292 16942
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35028 17890 35084 17892
rect 35028 17838 35030 17890
rect 35030 17838 35082 17890
rect 35082 17838 35084 17890
rect 35028 17836 35084 17838
rect 35420 17724 35476 17780
rect 34524 17612 34580 17668
rect 35308 17666 35364 17668
rect 35308 17614 35310 17666
rect 35310 17614 35362 17666
rect 35362 17614 35364 17666
rect 35308 17612 35364 17614
rect 34188 17388 34244 17444
rect 34412 17276 34468 17332
rect 34412 16828 34468 16884
rect 33236 16156 33292 16212
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 33124 15596 33180 15652
rect 33628 15314 33684 15316
rect 33628 15262 33630 15314
rect 33630 15262 33682 15314
rect 33682 15262 33684 15314
rect 33628 15260 33684 15262
rect 33740 15148 33796 15204
rect 33404 14588 33460 14644
rect 34076 15148 34132 15204
rect 34916 15314 34972 15316
rect 34916 15262 34918 15314
rect 34918 15262 34970 15314
rect 34970 15262 34972 15314
rect 34916 15260 34972 15262
rect 35084 15148 35140 15204
rect 34468 15090 34524 15092
rect 34468 15038 34470 15090
rect 34470 15038 34522 15090
rect 34522 15038 34524 15090
rect 34468 15036 34524 15038
rect 33516 13468 33572 13524
rect 32564 12402 32620 12404
rect 32564 12350 32566 12402
rect 32566 12350 32618 12402
rect 32618 12350 32620 12402
rect 32564 12348 32620 12350
rect 33068 12796 33124 12852
rect 32620 12012 32676 12068
rect 31724 11506 31780 11508
rect 31724 11454 31726 11506
rect 31726 11454 31778 11506
rect 31778 11454 31780 11506
rect 31724 11452 31780 11454
rect 31836 11379 31892 11396
rect 31836 11340 31838 11379
rect 31838 11340 31890 11379
rect 31890 11340 31892 11379
rect 31836 10668 31892 10724
rect 32956 12178 33012 12180
rect 32956 12126 32958 12178
rect 32958 12126 33010 12178
rect 33010 12126 33012 12178
rect 32956 12124 33012 12126
rect 33740 13692 33796 13748
rect 34300 14476 34356 14532
rect 35196 15036 35252 15092
rect 35980 17442 36036 17444
rect 35980 17390 35982 17442
rect 35982 17390 36034 17442
rect 36034 17390 36036 17442
rect 35980 17388 36036 17390
rect 35756 16716 35812 16772
rect 35756 15277 35758 15316
rect 35758 15277 35810 15316
rect 35810 15277 35812 15316
rect 35756 15260 35812 15277
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35532 14700 35588 14756
rect 35644 14588 35700 14644
rect 36652 19292 36708 19348
rect 36540 19234 36596 19236
rect 36540 19182 36542 19234
rect 36542 19182 36594 19234
rect 36594 19182 36596 19234
rect 36540 19180 36596 19182
rect 36652 18732 36708 18788
rect 36428 18450 36484 18452
rect 36428 18398 36430 18450
rect 36430 18398 36482 18450
rect 36482 18398 36484 18450
rect 36428 18396 36484 18398
rect 37100 19404 37156 19460
rect 36988 18620 37044 18676
rect 36876 18508 36932 18564
rect 36204 16268 36260 16324
rect 36764 16716 36820 16772
rect 36484 16210 36540 16212
rect 36484 16158 36486 16210
rect 36486 16158 36538 16210
rect 36538 16158 36540 16210
rect 36484 16156 36540 16158
rect 37100 19234 37156 19236
rect 37100 19182 37102 19234
rect 37102 19182 37154 19234
rect 37154 19182 37156 19234
rect 37100 19180 37156 19182
rect 37100 18508 37156 18564
rect 37548 21420 37604 21476
rect 37548 20300 37604 20356
rect 37996 21644 38052 21700
rect 37884 21474 37940 21476
rect 37884 21422 37886 21474
rect 37886 21422 37938 21474
rect 37938 21422 37940 21474
rect 37884 21420 37940 21422
rect 38668 23154 38724 23156
rect 38668 23102 38670 23154
rect 38670 23102 38722 23154
rect 38722 23102 38724 23154
rect 38668 23100 38724 23102
rect 38220 21644 38276 21700
rect 38220 21420 38276 21476
rect 37660 19964 37716 20020
rect 38108 20300 38164 20356
rect 37884 19852 37940 19908
rect 37660 18508 37716 18564
rect 38556 19981 38558 20020
rect 38558 19981 38610 20020
rect 38610 19981 38612 20020
rect 38556 19964 38612 19981
rect 38444 19906 38500 19908
rect 38444 19854 38446 19906
rect 38446 19854 38498 19906
rect 38498 19854 38500 19906
rect 38444 19852 38500 19854
rect 39172 24108 39228 24164
rect 39788 25116 39844 25172
rect 39564 23996 39620 24052
rect 39452 23938 39508 23940
rect 39452 23886 39454 23938
rect 39454 23886 39506 23938
rect 39506 23886 39508 23938
rect 39452 23884 39508 23886
rect 40012 25340 40068 25396
rect 40292 25228 40348 25284
rect 41132 25228 41188 25284
rect 42140 28924 42196 28980
rect 42700 29932 42756 29988
rect 42140 28364 42196 28420
rect 42644 28082 42700 28084
rect 42644 28030 42646 28082
rect 42646 28030 42698 28082
rect 42698 28030 42700 28082
rect 42644 28028 42700 28030
rect 42924 30156 42980 30212
rect 44268 31388 44324 31444
rect 45164 36482 45220 36484
rect 45164 36430 45166 36482
rect 45166 36430 45218 36482
rect 45218 36430 45220 36482
rect 45164 36428 45220 36430
rect 45164 35868 45220 35924
rect 45164 35196 45220 35252
rect 45276 35644 45332 35700
rect 45612 35644 45668 35700
rect 45276 35308 45332 35364
rect 45612 35196 45668 35252
rect 45444 34748 45500 34804
rect 46508 38220 46564 38276
rect 46620 38556 46676 38612
rect 46060 38108 46116 38164
rect 46956 43314 47012 43316
rect 46956 43262 46958 43314
rect 46958 43262 47010 43314
rect 47010 43262 47012 43314
rect 46956 43260 47012 43262
rect 46956 41468 47012 41524
rect 46956 40460 47012 40516
rect 47180 43036 47236 43092
rect 47068 40908 47124 40964
rect 47516 44268 47572 44324
rect 47628 44492 47684 44548
rect 47964 45106 48020 45108
rect 47964 45054 47966 45106
rect 47966 45054 48018 45106
rect 48018 45054 48020 45106
rect 47964 45052 48020 45054
rect 48972 47068 49028 47124
rect 48636 46674 48692 46676
rect 48636 46622 48638 46674
rect 48638 46622 48690 46674
rect 48690 46622 48692 46674
rect 48636 46620 48692 46622
rect 48972 46562 49028 46564
rect 48972 46510 48974 46562
rect 48974 46510 49026 46562
rect 49026 46510 49028 46562
rect 48972 46508 49028 46510
rect 49084 45276 49140 45332
rect 48636 45164 48692 45220
rect 48300 44604 48356 44660
rect 49140 45106 49196 45108
rect 49140 45054 49142 45106
rect 49142 45054 49194 45106
rect 49194 45054 49196 45106
rect 49140 45052 49196 45054
rect 48860 44492 48916 44548
rect 47516 43538 47572 43540
rect 47516 43486 47518 43538
rect 47518 43486 47570 43538
rect 47570 43486 47572 43538
rect 47516 43484 47572 43486
rect 47852 43148 47908 43204
rect 47964 43036 48020 43092
rect 47964 41970 48020 41972
rect 47964 41918 47966 41970
rect 47966 41918 48018 41970
rect 48018 41918 48020 41970
rect 47964 41916 48020 41918
rect 48300 41916 48356 41972
rect 48412 43148 48468 43204
rect 48300 41468 48356 41524
rect 47068 40348 47124 40404
rect 48076 40684 48132 40740
rect 46956 39788 47012 39844
rect 47068 39676 47124 39732
rect 47234 39228 47290 39284
rect 48524 41468 48580 41524
rect 48524 41186 48580 41188
rect 48524 41134 48526 41186
rect 48526 41134 48578 41186
rect 48578 41134 48580 41186
rect 48524 41132 48580 41134
rect 48412 40684 48468 40740
rect 48412 40460 48468 40516
rect 48300 39340 48356 39396
rect 48972 41746 49028 41748
rect 48972 41694 48974 41746
rect 48974 41694 49026 41746
rect 49026 41694 49028 41746
rect 48972 41692 49028 41694
rect 48748 41132 48804 41188
rect 48860 41020 48916 41076
rect 49084 40572 49140 40628
rect 49084 40236 49140 40292
rect 46732 38108 46788 38164
rect 46844 38834 46900 38836
rect 46844 38782 46846 38834
rect 46846 38782 46898 38834
rect 46898 38782 46900 38834
rect 46844 38780 46900 38782
rect 46284 37772 46340 37828
rect 46620 37436 46676 37492
rect 47404 38810 47406 38836
rect 47406 38810 47458 38836
rect 47458 38810 47460 38836
rect 47404 38780 47460 38810
rect 48860 38780 48916 38836
rect 47908 38444 47964 38500
rect 47740 37548 47796 37604
rect 45836 35868 45892 35924
rect 45948 36428 46004 36484
rect 46116 36370 46172 36372
rect 46116 36318 46118 36370
rect 46118 36318 46170 36370
rect 46170 36318 46172 36370
rect 46116 36316 46172 36318
rect 45836 35196 45892 35252
rect 46508 35698 46564 35700
rect 46508 35646 46510 35698
rect 46510 35646 46562 35698
rect 46562 35646 46564 35698
rect 46508 35644 46564 35646
rect 46172 34860 46228 34916
rect 46396 34914 46452 34916
rect 46396 34862 46398 34914
rect 46398 34862 46450 34914
rect 46450 34862 46452 34914
rect 46396 34860 46452 34862
rect 46284 34748 46340 34804
rect 45948 34412 46004 34468
rect 46732 36316 46788 36372
rect 46956 34972 47012 35028
rect 47180 35868 47236 35924
rect 48188 37772 48244 37828
rect 47292 35756 47348 35812
rect 47740 36204 47796 36260
rect 44716 31948 44772 32004
rect 43708 30828 43764 30884
rect 44940 30828 44996 30884
rect 45052 32562 45108 32564
rect 45052 32510 45054 32562
rect 45054 32510 45106 32562
rect 45106 32510 45108 32562
rect 45052 32508 45108 32510
rect 43260 30044 43316 30100
rect 43596 30182 43652 30212
rect 43596 30156 43598 30182
rect 43598 30156 43650 30182
rect 43650 30156 43652 30182
rect 43372 29932 43428 29988
rect 44492 29932 44548 29988
rect 44380 29484 44436 29540
rect 43932 28866 43988 28868
rect 43932 28814 43934 28866
rect 43934 28814 43986 28866
rect 43986 28814 43988 28866
rect 43932 28812 43988 28814
rect 43148 28614 43204 28644
rect 43148 28588 43150 28614
rect 43150 28588 43202 28614
rect 43202 28588 43204 28614
rect 42812 27858 42868 27860
rect 42812 27806 42814 27858
rect 42814 27806 42866 27858
rect 42866 27806 42868 27858
rect 42812 27804 42868 27806
rect 42028 26124 42084 26180
rect 40236 24050 40292 24052
rect 40236 23998 40238 24050
rect 40238 23998 40290 24050
rect 40290 23998 40292 24050
rect 40236 23996 40292 23998
rect 41356 23884 41412 23940
rect 39676 23324 39732 23380
rect 38892 22428 38948 22484
rect 40404 23378 40460 23380
rect 40404 23326 40406 23378
rect 40406 23326 40458 23378
rect 40458 23326 40460 23378
rect 40404 23324 40460 23326
rect 40908 23324 40964 23380
rect 40124 23100 40180 23156
rect 39956 23042 40012 23044
rect 39956 22990 39958 23042
rect 39958 22990 40010 23042
rect 40010 22990 40012 23042
rect 39956 22988 40012 22990
rect 40124 22316 40180 22372
rect 40348 22540 40404 22596
rect 39228 22092 39284 22148
rect 38892 21586 38948 21588
rect 38892 21534 38894 21586
rect 38894 21534 38946 21586
rect 38946 21534 38948 21586
rect 38892 21532 38948 21534
rect 38780 21308 38836 21364
rect 38892 21196 38948 21252
rect 39564 21196 39620 21252
rect 40012 21362 40068 21364
rect 40012 21310 40014 21362
rect 40014 21310 40066 21362
rect 40066 21310 40068 21362
rect 40012 21308 40068 21310
rect 38668 19740 38724 19796
rect 38892 19516 38948 19572
rect 39004 19964 39060 20020
rect 37548 16882 37604 16884
rect 37548 16830 37550 16882
rect 37550 16830 37602 16882
rect 37602 16830 37604 16882
rect 37548 16828 37604 16830
rect 36988 16156 37044 16212
rect 37660 16098 37716 16100
rect 37660 16046 37662 16098
rect 37662 16046 37714 16098
rect 37714 16046 37716 16098
rect 37660 16044 37716 16046
rect 37996 18060 38052 18116
rect 37884 17442 37940 17444
rect 37884 17390 37886 17442
rect 37886 17390 37938 17442
rect 37938 17390 37940 17442
rect 37884 17388 37940 17390
rect 38332 18508 38388 18564
rect 38780 18396 38836 18452
rect 36540 15314 36596 15316
rect 36540 15262 36542 15314
rect 36542 15262 36594 15314
rect 36594 15262 36596 15314
rect 36540 15260 36596 15262
rect 38556 16716 38612 16772
rect 39116 18396 39172 18452
rect 39900 19852 39956 19908
rect 40124 19740 40180 19796
rect 39788 19516 39844 19572
rect 39900 19404 39956 19460
rect 39564 18060 39620 18116
rect 39900 18620 39956 18676
rect 40908 22482 40964 22484
rect 40908 22430 40910 22482
rect 40910 22430 40962 22482
rect 40962 22430 40964 22482
rect 40908 22428 40964 22430
rect 41020 22652 41076 22708
rect 40348 19404 40404 19460
rect 40460 21420 40516 21476
rect 40236 18396 40292 18452
rect 41244 22540 41300 22596
rect 41916 25506 41972 25508
rect 41916 25454 41918 25506
rect 41918 25454 41970 25506
rect 41970 25454 41972 25506
rect 41916 25452 41972 25454
rect 41468 22652 41524 22708
rect 41916 23100 41972 23156
rect 42532 26178 42588 26180
rect 42532 26126 42534 26178
rect 42534 26126 42586 26178
rect 42586 26126 42588 26178
rect 42532 26124 42588 26126
rect 44716 30156 44772 30212
rect 44940 29932 44996 29988
rect 44828 29820 44884 29876
rect 45612 33180 45668 33236
rect 46620 33516 46676 33572
rect 47964 34354 48020 34356
rect 47964 34302 47966 34354
rect 47966 34302 48018 34354
rect 48018 34302 48020 34354
rect 47964 34300 48020 34302
rect 46844 33404 46900 33460
rect 45388 32396 45444 32452
rect 45220 31948 45276 32004
rect 45836 33068 45892 33124
rect 46116 33180 46172 33236
rect 45948 32508 46004 32564
rect 46844 32284 46900 32340
rect 47404 33516 47460 33572
rect 48636 38444 48692 38500
rect 48524 38162 48580 38164
rect 48524 38110 48526 38162
rect 48526 38110 48578 38162
rect 48578 38110 48580 38162
rect 48524 38108 48580 38110
rect 48524 34300 48580 34356
rect 48524 32732 48580 32788
rect 48748 37772 48804 37828
rect 49196 38108 49252 38164
rect 49308 41916 49364 41972
rect 49420 41692 49476 41748
rect 49420 40236 49476 40292
rect 49084 37436 49140 37492
rect 48860 36876 48916 36932
rect 48860 36092 48916 36148
rect 48972 35980 49028 36036
rect 48748 35868 48804 35924
rect 49084 35698 49140 35700
rect 49084 35646 49086 35698
rect 49086 35646 49138 35698
rect 49138 35646 49140 35698
rect 49084 35644 49140 35646
rect 49420 34860 49476 34916
rect 49084 34802 49140 34804
rect 49084 34750 49086 34802
rect 49086 34750 49138 34802
rect 49138 34750 49140 34802
rect 49084 34748 49140 34750
rect 48972 34018 49028 34020
rect 48972 33966 48974 34018
rect 48974 33966 49026 34018
rect 49026 33966 49028 34018
rect 48972 33964 49028 33966
rect 45724 31948 45780 32004
rect 45164 30182 45220 30212
rect 45164 30156 45166 30182
rect 45166 30156 45218 30182
rect 45218 30156 45220 30182
rect 46788 31276 46844 31332
rect 46172 31218 46228 31220
rect 46172 31166 46174 31218
rect 46174 31166 46226 31218
rect 46226 31166 46228 31218
rect 46172 31164 46228 31166
rect 45500 30882 45556 30884
rect 45500 30830 45502 30882
rect 45502 30830 45554 30882
rect 45554 30830 45556 30882
rect 45500 30828 45556 30830
rect 46396 30210 46452 30212
rect 46396 30158 46398 30210
rect 46398 30158 46450 30210
rect 46450 30158 46452 30210
rect 46396 30156 46452 30158
rect 46228 29820 46284 29876
rect 46452 29538 46508 29540
rect 46452 29486 46454 29538
rect 46454 29486 46506 29538
rect 46506 29486 46508 29538
rect 46452 29484 46508 29486
rect 47964 32562 48020 32564
rect 47964 32510 47966 32562
rect 47966 32510 48018 32562
rect 48018 32510 48020 32562
rect 47964 32508 48020 32510
rect 48636 32562 48692 32564
rect 48636 32510 48638 32562
rect 48638 32510 48690 32562
rect 48690 32510 48692 32562
rect 48636 32508 48692 32510
rect 48076 32284 48132 32340
rect 47404 31276 47460 31332
rect 47740 31164 47796 31220
rect 47908 31388 47964 31444
rect 48972 32732 49028 32788
rect 48860 32002 48916 32004
rect 48860 31950 48862 32002
rect 48862 31950 48914 32002
rect 48914 31950 48916 32002
rect 48860 31948 48916 31950
rect 49308 34130 49364 34132
rect 49308 34078 49310 34130
rect 49310 34078 49362 34130
rect 49362 34078 49364 34130
rect 49308 34076 49364 34078
rect 49308 32508 49364 32564
rect 48524 30156 48580 30212
rect 47628 29932 47684 29988
rect 44604 28588 44660 28644
rect 45500 28588 45556 28644
rect 44716 27804 44772 27860
rect 43820 26348 43876 26404
rect 48972 29820 49028 29876
rect 43036 26124 43092 26180
rect 43464 25506 43520 25508
rect 43464 25454 43466 25506
rect 43466 25454 43518 25506
rect 43518 25454 43520 25506
rect 43464 25452 43520 25454
rect 42588 25340 42644 25396
rect 43820 25116 43876 25172
rect 43708 24668 43764 24724
rect 42140 24444 42196 24500
rect 42476 24332 42532 24388
rect 42028 22876 42084 22932
rect 42980 23938 43036 23940
rect 42980 23886 42982 23938
rect 42982 23886 43034 23938
rect 43034 23886 43036 23938
rect 42980 23884 43036 23886
rect 41132 21586 41188 21588
rect 41132 21534 41134 21586
rect 41134 21534 41186 21586
rect 41186 21534 41188 21586
rect 41132 21532 41188 21534
rect 41300 21420 41356 21476
rect 40908 20972 40964 21028
rect 40908 20412 40964 20468
rect 41356 20300 41412 20356
rect 41356 19906 41412 19908
rect 41356 19854 41358 19906
rect 41358 19854 41410 19906
rect 41410 19854 41412 19906
rect 41356 19852 41412 19854
rect 40684 19516 40740 19572
rect 43484 22988 43540 23044
rect 42252 21644 42308 21700
rect 41748 21362 41804 21364
rect 41748 21310 41750 21362
rect 41750 21310 41802 21362
rect 41802 21310 41804 21362
rect 41748 21308 41804 21310
rect 41804 20412 41860 20468
rect 42140 21420 42196 21476
rect 41916 20188 41972 20244
rect 42028 19852 42084 19908
rect 43372 22204 43428 22260
rect 42700 21420 42756 21476
rect 42364 21308 42420 21364
rect 42588 21196 42644 21252
rect 42364 20076 42420 20132
rect 39900 17948 39956 18004
rect 39004 17052 39060 17108
rect 37100 15036 37156 15092
rect 36988 14642 37044 14644
rect 36988 14590 36990 14642
rect 36990 14590 37042 14642
rect 37042 14590 37044 14642
rect 36988 14588 37044 14590
rect 35980 14476 36036 14532
rect 38332 15036 38388 15092
rect 37324 14700 37380 14756
rect 37660 14530 37716 14532
rect 37660 14478 37662 14530
rect 37662 14478 37714 14530
rect 37714 14478 37716 14530
rect 37660 14476 37716 14478
rect 38668 14530 38724 14532
rect 38668 14478 38670 14530
rect 38670 14478 38722 14530
rect 38722 14478 38724 14530
rect 38668 14476 38724 14478
rect 38220 14028 38276 14084
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 37772 13074 37828 13076
rect 37772 13022 37774 13074
rect 37774 13022 37826 13074
rect 37826 13022 37828 13074
rect 37772 13020 37828 13022
rect 34300 12796 34356 12852
rect 33740 12066 33796 12068
rect 33740 12014 33742 12066
rect 33742 12014 33794 12066
rect 33794 12014 33796 12066
rect 33740 12012 33796 12014
rect 33628 11228 33684 11284
rect 32508 10332 32564 10388
rect 33180 10668 33236 10724
rect 33628 10332 33684 10388
rect 31612 9660 31668 9716
rect 30604 8988 30660 9044
rect 29260 7586 29316 7588
rect 29260 7534 29262 7586
rect 29262 7534 29314 7586
rect 29314 7534 29316 7586
rect 29260 7532 29316 7534
rect 31276 7532 31332 7588
rect 29484 7420 29540 7476
rect 30716 7474 30772 7476
rect 30716 7422 30718 7474
rect 30718 7422 30770 7474
rect 30770 7422 30772 7474
rect 30716 7420 30772 7422
rect 28644 6748 28700 6804
rect 29372 6748 29428 6804
rect 27020 6524 27076 6580
rect 25396 6130 25452 6132
rect 25396 6078 25398 6130
rect 25398 6078 25450 6130
rect 25450 6078 25452 6130
rect 25396 6076 25452 6078
rect 25844 6130 25900 6132
rect 25844 6078 25846 6130
rect 25846 6078 25898 6130
rect 25898 6078 25900 6130
rect 25844 6076 25900 6078
rect 26516 6130 26572 6132
rect 26516 6078 26518 6130
rect 26518 6078 26570 6130
rect 26570 6078 26572 6130
rect 26516 6076 26572 6078
rect 23100 5122 23156 5124
rect 23100 5070 23102 5122
rect 23102 5070 23154 5122
rect 23154 5070 23156 5122
rect 23100 5068 23156 5070
rect 22932 4620 22988 4676
rect 22540 4508 22596 4564
rect 22858 4450 22914 4452
rect 22858 4398 22860 4450
rect 22860 4398 22912 4450
rect 22912 4398 22914 4450
rect 22858 4396 22914 4398
rect 23772 5068 23828 5124
rect 23604 4620 23660 4676
rect 23772 4450 23828 4452
rect 23772 4398 23774 4450
rect 23774 4398 23826 4450
rect 23826 4398 23828 4450
rect 23772 4396 23828 4398
rect 24444 5068 24500 5124
rect 25564 5122 25620 5124
rect 25564 5070 25566 5122
rect 25566 5070 25618 5122
rect 25618 5070 25620 5122
rect 25564 5068 25620 5070
rect 25396 4620 25452 4676
rect 25228 4450 25284 4452
rect 25228 4398 25230 4450
rect 25230 4398 25282 4450
rect 25282 4398 25284 4450
rect 25228 4396 25284 4398
rect 26348 5122 26404 5124
rect 26348 5070 26350 5122
rect 26350 5070 26402 5122
rect 26402 5070 26404 5122
rect 26348 5068 26404 5070
rect 26908 5068 26964 5124
rect 25788 4396 25844 4452
rect 26142 4508 26198 4564
rect 25900 4338 25956 4340
rect 25900 4286 25902 4338
rect 25902 4286 25954 4338
rect 25954 4286 25956 4338
rect 25900 4284 25956 4286
rect 22428 3612 22484 3668
rect 24780 3666 24836 3668
rect 24780 3614 24782 3666
rect 24782 3614 24834 3666
rect 24834 3614 24836 3666
rect 24780 3612 24836 3614
rect 22652 3388 22708 3444
rect 27916 5906 27972 5908
rect 27916 5854 27918 5906
rect 27918 5854 27970 5906
rect 27970 5854 27972 5906
rect 27916 5852 27972 5854
rect 29260 5852 29316 5908
rect 29596 6076 29652 6132
rect 29932 6690 29988 6692
rect 29932 6638 29934 6690
rect 29934 6638 29986 6690
rect 29986 6638 29988 6690
rect 29932 6636 29988 6638
rect 30156 6524 30212 6580
rect 30492 6690 30548 6692
rect 30492 6638 30494 6690
rect 30494 6638 30546 6690
rect 30546 6638 30548 6690
rect 30492 6636 30548 6638
rect 31500 8428 31556 8484
rect 33292 9660 33348 9716
rect 34300 11788 34356 11844
rect 35644 11900 35700 11956
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35980 11452 36036 11508
rect 36540 11900 36596 11956
rect 34412 11228 34468 11284
rect 36204 11340 36260 11396
rect 34356 10892 34412 10948
rect 35700 10668 35756 10724
rect 34356 10108 34412 10164
rect 33180 8540 33236 8596
rect 35308 10332 35364 10388
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35252 9996 35308 10052
rect 35420 9884 35476 9940
rect 35868 9996 35924 10052
rect 32396 8258 32452 8260
rect 32396 8206 32398 8258
rect 32398 8206 32450 8258
rect 32450 8206 32452 8258
rect 32396 8204 32452 8206
rect 31612 7532 31668 7588
rect 30716 6524 30772 6580
rect 30380 6076 30436 6132
rect 30268 5906 30324 5908
rect 30268 5854 30270 5906
rect 30270 5854 30322 5906
rect 30322 5854 30324 5906
rect 30268 5852 30324 5854
rect 28196 5180 28252 5236
rect 27132 5068 27188 5124
rect 27468 5068 27524 5124
rect 27916 4956 27972 5012
rect 28476 5180 28532 5236
rect 29036 4956 29092 5012
rect 28196 4844 28252 4900
rect 28812 4844 28868 4900
rect 28812 3500 28868 3556
rect 27748 3388 27804 3444
rect 29484 5122 29540 5124
rect 29484 5070 29486 5122
rect 29486 5070 29538 5122
rect 29538 5070 29540 5122
rect 29484 5068 29540 5070
rect 29484 3612 29540 3668
rect 29148 3554 29204 3556
rect 29148 3502 29150 3554
rect 29150 3502 29202 3554
rect 29202 3502 29204 3554
rect 29148 3500 29204 3502
rect 29596 3500 29652 3556
rect 30716 5180 30772 5236
rect 30492 5122 30548 5124
rect 30492 5070 30494 5122
rect 30494 5070 30546 5122
rect 30546 5070 30548 5122
rect 30492 5068 30548 5070
rect 31388 5404 31444 5460
rect 31164 5068 31220 5124
rect 30156 3554 30212 3556
rect 30156 3502 30158 3554
rect 30158 3502 30210 3554
rect 30210 3502 30212 3554
rect 30156 3500 30212 3502
rect 30604 3666 30660 3668
rect 30604 3614 30606 3666
rect 30606 3614 30658 3666
rect 30658 3614 30660 3666
rect 30604 3612 30660 3614
rect 31780 7474 31836 7476
rect 31780 7422 31782 7474
rect 31782 7422 31834 7474
rect 31834 7422 31836 7474
rect 31780 7420 31836 7422
rect 33180 7084 33236 7140
rect 31836 6690 31892 6692
rect 31836 6638 31838 6690
rect 31838 6638 31890 6690
rect 31890 6638 31892 6690
rect 31836 6636 31892 6638
rect 32340 6690 32396 6692
rect 32340 6638 32342 6690
rect 32342 6638 32394 6690
rect 32394 6638 32396 6690
rect 32340 6636 32396 6638
rect 31612 5906 31668 5908
rect 31612 5854 31614 5906
rect 31614 5854 31666 5906
rect 31666 5854 31668 5906
rect 31612 5852 31668 5854
rect 32844 6690 32900 6692
rect 32844 6638 32846 6690
rect 32846 6638 32898 6690
rect 32898 6638 32900 6690
rect 32844 6636 32900 6638
rect 35644 8764 35700 8820
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 34188 8204 34244 8260
rect 34748 8204 34804 8260
rect 33516 8146 33572 8148
rect 33516 8094 33518 8146
rect 33518 8094 33570 8146
rect 33570 8094 33572 8146
rect 33516 8092 33572 8094
rect 34188 7644 34244 7700
rect 34916 8258 34972 8260
rect 34916 8206 34918 8258
rect 34918 8206 34970 8258
rect 34970 8206 34972 8258
rect 34916 8204 34972 8206
rect 35644 8258 35700 8260
rect 35644 8206 35646 8258
rect 35646 8206 35698 8258
rect 35698 8206 35700 8258
rect 35644 8204 35700 8206
rect 35868 8764 35924 8820
rect 35980 9884 36036 9940
rect 36876 11394 36932 11396
rect 36876 11342 36878 11394
rect 36878 11342 36930 11394
rect 36930 11342 36932 11394
rect 36876 11340 36932 11342
rect 36988 10108 37044 10164
rect 37772 11452 37828 11508
rect 37156 9996 37212 10052
rect 37772 9996 37828 10052
rect 37996 11340 38052 11396
rect 38108 13020 38164 13076
rect 37996 11116 38052 11172
rect 40124 16828 40180 16884
rect 39340 16716 39396 16772
rect 40012 16716 40068 16772
rect 39116 15484 39172 15540
rect 39228 15036 39284 15092
rect 38500 13522 38556 13524
rect 38500 13470 38502 13522
rect 38502 13470 38554 13522
rect 38554 13470 38556 13522
rect 38500 13468 38556 13470
rect 39228 14252 39284 14308
rect 40404 17836 40460 17892
rect 41244 18413 41246 18452
rect 41246 18413 41298 18452
rect 41298 18413 41300 18452
rect 41244 18396 41300 18413
rect 43148 20748 43204 20804
rect 44044 26348 44100 26404
rect 45108 26348 45164 26404
rect 44940 26290 44996 26292
rect 44940 26238 44942 26290
rect 44942 26238 44994 26290
rect 44994 26238 44996 26290
rect 44940 26236 44996 26238
rect 44324 25788 44380 25844
rect 44716 25228 44772 25284
rect 44828 25452 44884 25508
rect 44566 25116 44622 25172
rect 44380 24722 44436 24724
rect 44380 24670 44382 24722
rect 44382 24670 44434 24722
rect 44434 24670 44436 24722
rect 44380 24668 44436 24670
rect 46284 26796 46340 26852
rect 46116 26236 46172 26292
rect 47404 26962 47460 26964
rect 47404 26910 47406 26962
rect 47406 26910 47458 26962
rect 47458 26910 47460 26962
rect 47404 26908 47460 26910
rect 46620 26236 46676 26292
rect 47628 26290 47684 26292
rect 46732 25788 46788 25844
rect 47628 26238 47630 26290
rect 47630 26238 47682 26290
rect 47682 26238 47684 26290
rect 47628 26236 47684 26238
rect 45612 25116 45668 25172
rect 45388 24780 45444 24836
rect 45836 24780 45892 24836
rect 44212 23772 44268 23828
rect 44548 23212 44604 23268
rect 44828 23772 44884 23828
rect 44044 22876 44100 22932
rect 44940 23324 44996 23380
rect 45388 23154 45444 23156
rect 45388 23102 45390 23154
rect 45390 23102 45442 23154
rect 45442 23102 45444 23154
rect 45388 23100 45444 23102
rect 45108 22930 45164 22932
rect 45108 22878 45110 22930
rect 45110 22878 45162 22930
rect 45162 22878 45164 22930
rect 45108 22876 45164 22878
rect 44492 22540 44548 22596
rect 43820 21420 43876 21476
rect 43988 22316 44044 22372
rect 44156 22258 44212 22260
rect 44156 22206 44158 22258
rect 44158 22206 44210 22258
rect 44210 22206 44212 22258
rect 44156 22204 44212 22206
rect 45724 22540 45780 22596
rect 45948 23212 46004 23268
rect 44828 22204 44884 22260
rect 44604 21644 44660 21700
rect 45500 21644 45556 21700
rect 47068 25116 47124 25172
rect 46732 23938 46788 23940
rect 46732 23886 46734 23938
rect 46734 23886 46786 23938
rect 46786 23886 46788 23938
rect 46732 23884 46788 23886
rect 48860 29484 48916 29540
rect 48076 29426 48132 29428
rect 48076 29374 48078 29426
rect 48078 29374 48130 29426
rect 48130 29374 48132 29426
rect 48076 29372 48132 29374
rect 49084 29372 49140 29428
rect 49308 27580 49364 27636
rect 48244 27132 48300 27188
rect 49308 27132 49364 27188
rect 47852 25788 47908 25844
rect 47404 24668 47460 24724
rect 47628 25116 47684 25172
rect 47628 24780 47684 24836
rect 47964 24332 48020 24388
rect 47180 23884 47236 23940
rect 47628 23938 47684 23940
rect 47628 23886 47630 23938
rect 47630 23886 47682 23938
rect 47682 23886 47684 23938
rect 47628 23884 47684 23886
rect 46172 23042 46228 23044
rect 46172 22990 46174 23042
rect 46174 22990 46226 23042
rect 46226 22990 46228 23042
rect 46172 22988 46228 22990
rect 46060 21644 46116 21700
rect 44884 21586 44940 21588
rect 44884 21534 44886 21586
rect 44886 21534 44938 21586
rect 44938 21534 44940 21586
rect 44884 21532 44940 21534
rect 47740 23100 47796 23156
rect 48860 24722 48916 24724
rect 48860 24670 48862 24722
rect 48862 24670 48914 24722
rect 48914 24670 48916 24722
rect 48860 24668 48916 24670
rect 48748 24332 48804 24388
rect 48188 23884 48244 23940
rect 48580 23938 48636 23940
rect 48580 23886 48582 23938
rect 48582 23886 48634 23938
rect 48634 23886 48636 23938
rect 48580 23884 48636 23886
rect 46732 22540 46788 22596
rect 46172 21586 46228 21588
rect 46172 21534 46174 21586
rect 46174 21534 46226 21586
rect 46226 21534 46228 21586
rect 46172 21532 46228 21534
rect 43988 21196 44044 21252
rect 45276 21308 45332 21364
rect 44268 20802 44324 20804
rect 44268 20750 44270 20802
rect 44270 20750 44322 20802
rect 44322 20750 44324 20802
rect 44268 20748 44324 20750
rect 45052 20748 45108 20804
rect 45836 21196 45892 21252
rect 42700 20412 42756 20468
rect 42920 20076 42976 20132
rect 42644 19906 42700 19908
rect 42644 19854 42646 19906
rect 42646 19854 42698 19906
rect 42698 19854 42700 19906
rect 42644 19852 42700 19854
rect 46060 20242 46116 20244
rect 46060 20190 46062 20242
rect 46062 20190 46114 20242
rect 46114 20190 46116 20242
rect 46060 20188 46116 20190
rect 43596 20076 43652 20132
rect 45332 20130 45388 20132
rect 45332 20078 45334 20130
rect 45334 20078 45386 20130
rect 45386 20078 45388 20130
rect 45332 20076 45388 20078
rect 45948 20076 46004 20132
rect 43708 19964 43764 20020
rect 43484 19740 43540 19796
rect 42920 19516 42976 19572
rect 43484 19404 43540 19460
rect 41804 18450 41860 18452
rect 41804 18398 41806 18450
rect 41806 18398 41858 18450
rect 41858 18398 41860 18450
rect 41804 18396 41860 18398
rect 41356 18060 41412 18116
rect 41804 18172 41860 18228
rect 42364 18284 42420 18340
rect 41692 17388 41748 17444
rect 41076 16994 41132 16996
rect 41076 16942 41078 16994
rect 41078 16942 41130 16994
rect 41130 16942 41132 16994
rect 41076 16940 41132 16942
rect 41244 16828 41300 16884
rect 40236 16716 40292 16772
rect 40236 16098 40292 16100
rect 40236 16046 40238 16098
rect 40238 16046 40290 16098
rect 40290 16046 40292 16098
rect 40236 16044 40292 16046
rect 39900 15484 39956 15540
rect 40124 14700 40180 14756
rect 39956 14476 40012 14532
rect 39900 14252 39956 14308
rect 38892 13020 38948 13076
rect 39396 13074 39452 13076
rect 39396 13022 39398 13074
rect 39398 13022 39450 13074
rect 39450 13022 39452 13074
rect 39396 13020 39452 13022
rect 39900 13074 39956 13076
rect 39900 13022 39902 13074
rect 39902 13022 39954 13074
rect 39954 13022 39956 13074
rect 39900 13020 39956 13022
rect 38220 11452 38276 11508
rect 38108 10220 38164 10276
rect 38220 10556 38276 10612
rect 38332 9938 38388 9940
rect 38332 9886 38334 9938
rect 38334 9886 38386 9938
rect 38386 9886 38388 9938
rect 38332 9884 38388 9886
rect 37548 8652 37604 8708
rect 34860 7474 34916 7476
rect 34860 7422 34862 7474
rect 34862 7422 34914 7474
rect 34914 7422 34916 7474
rect 34860 7420 34916 7422
rect 34244 7362 34300 7364
rect 34244 7310 34246 7362
rect 34246 7310 34298 7362
rect 34298 7310 34300 7362
rect 34244 7308 34300 7310
rect 33404 6748 33460 6804
rect 33292 6636 33348 6692
rect 33404 5906 33460 5908
rect 33404 5854 33406 5906
rect 33406 5854 33458 5906
rect 33458 5854 33460 5906
rect 33404 5852 33460 5854
rect 32060 5740 32116 5796
rect 31724 5404 31780 5460
rect 33628 5122 33684 5124
rect 33628 5070 33630 5122
rect 33630 5070 33682 5122
rect 33682 5070 33684 5122
rect 33628 5068 33684 5070
rect 31500 4844 31556 4900
rect 32508 4956 32564 5012
rect 34188 5869 34190 5908
rect 34190 5869 34242 5908
rect 34242 5869 34244 5908
rect 34188 5852 34244 5869
rect 35420 7474 35476 7476
rect 35420 7422 35422 7474
rect 35422 7422 35474 7474
rect 35474 7422 35476 7474
rect 35420 7420 35476 7422
rect 34972 7084 35028 7140
rect 38108 8258 38164 8260
rect 38108 8206 38110 8258
rect 38110 8206 38162 8258
rect 38162 8206 38164 8258
rect 38108 8204 38164 8206
rect 39564 12962 39620 12964
rect 39564 12910 39566 12962
rect 39566 12910 39618 12962
rect 39618 12910 39620 12962
rect 39564 12908 39620 12910
rect 39508 11954 39564 11956
rect 39508 11902 39510 11954
rect 39510 11902 39562 11954
rect 39562 11902 39564 11954
rect 39508 11900 39564 11902
rect 38668 11116 38724 11172
rect 38556 10332 38612 10388
rect 38892 10668 38948 10724
rect 39676 10668 39732 10724
rect 42588 18172 42644 18228
rect 43820 18060 43876 18116
rect 43708 17948 43764 18004
rect 41804 16492 41860 16548
rect 42476 16882 42532 16884
rect 42476 16830 42478 16882
rect 42478 16830 42530 16882
rect 42530 16830 42532 16882
rect 42476 16828 42532 16830
rect 42700 16882 42756 16884
rect 42700 16830 42702 16882
rect 42702 16830 42754 16882
rect 42754 16830 42756 16882
rect 42700 16828 42756 16830
rect 43484 16828 43540 16884
rect 42084 16658 42140 16660
rect 42084 16606 42086 16658
rect 42086 16606 42138 16658
rect 42138 16606 42140 16658
rect 42084 16604 42140 16606
rect 41804 15372 41860 15428
rect 41636 15202 41692 15204
rect 41636 15150 41638 15202
rect 41638 15150 41690 15202
rect 41690 15150 41692 15202
rect 41636 15148 41692 15150
rect 42364 15596 42420 15652
rect 42252 15277 42254 15316
rect 42254 15277 42306 15316
rect 42306 15277 42308 15316
rect 42252 15260 42308 15277
rect 42476 15484 42532 15540
rect 41468 14028 41524 14084
rect 40236 13970 40292 13972
rect 40236 13918 40238 13970
rect 40238 13918 40290 13970
rect 40290 13918 40292 13970
rect 40236 13916 40292 13918
rect 41692 13916 41748 13972
rect 41972 14028 42028 14084
rect 41244 13020 41300 13076
rect 40516 12908 40572 12964
rect 40012 10668 40068 10724
rect 39340 10444 39396 10500
rect 38668 10108 38724 10164
rect 38780 8988 38836 9044
rect 38500 8258 38556 8260
rect 38500 8206 38502 8258
rect 38502 8206 38554 8258
rect 38554 8206 38556 8258
rect 38500 8204 38556 8206
rect 38220 8092 38276 8148
rect 38556 7980 38612 8036
rect 36316 7420 36372 7476
rect 36540 7474 36596 7476
rect 36540 7422 36542 7474
rect 36542 7422 36594 7474
rect 36594 7422 36596 7474
rect 36540 7420 36596 7422
rect 37044 7420 37100 7476
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 34748 5906 34804 5908
rect 34748 5854 34750 5906
rect 34750 5854 34802 5906
rect 34802 5854 34804 5906
rect 34748 5852 34804 5854
rect 34972 6748 35028 6804
rect 34300 5794 34356 5796
rect 34300 5742 34302 5794
rect 34302 5742 34354 5794
rect 34354 5742 34356 5794
rect 34300 5740 34356 5742
rect 37044 6860 37100 6916
rect 37660 6972 37716 7028
rect 36092 6748 36148 6804
rect 35756 6636 35812 6692
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 33964 4956 34020 5012
rect 35084 4844 35140 4900
rect 33180 4338 33236 4340
rect 33180 4286 33182 4338
rect 33182 4286 33234 4338
rect 33234 4286 33236 4338
rect 33180 4284 33236 4286
rect 34636 3948 34692 4004
rect 33404 3612 33460 3668
rect 31612 3500 31668 3556
rect 29820 3388 29876 3444
rect 32396 3554 32452 3556
rect 32396 3502 32398 3554
rect 32398 3502 32450 3554
rect 32450 3502 32452 3554
rect 32396 3500 32452 3502
rect 35644 5180 35700 5236
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 35868 5068 35924 5124
rect 35084 3554 35140 3556
rect 35084 3502 35086 3554
rect 35086 3502 35138 3554
rect 35138 3502 35140 3554
rect 35084 3500 35140 3502
rect 37548 6690 37604 6692
rect 37548 6638 37550 6690
rect 37550 6638 37602 6690
rect 37602 6638 37604 6690
rect 37548 6636 37604 6638
rect 38312 7644 38368 7700
rect 38312 6972 38368 7028
rect 37436 6412 37492 6468
rect 37156 5234 37212 5236
rect 37156 5182 37158 5234
rect 37158 5182 37210 5234
rect 37210 5182 37212 5234
rect 37156 5180 37212 5182
rect 36764 4338 36820 4340
rect 36764 4286 36766 4338
rect 36766 4286 36818 4338
rect 36818 4286 36820 4338
rect 36764 4284 36820 4286
rect 37884 4172 37940 4228
rect 36988 3666 37044 3668
rect 36988 3614 36990 3666
rect 36990 3614 37042 3666
rect 37042 3614 37044 3666
rect 36988 3612 37044 3614
rect 38108 5180 38164 5236
rect 38668 7308 38724 7364
rect 38556 6690 38612 6692
rect 38556 6638 38558 6690
rect 38558 6638 38610 6690
rect 38610 6638 38612 6690
rect 38556 6636 38612 6638
rect 38444 5068 38500 5124
rect 38556 5628 38612 5684
rect 38220 4620 38276 4676
rect 39228 10332 39284 10388
rect 39004 9436 39060 9492
rect 39116 8652 39172 8708
rect 39340 10220 39396 10276
rect 39676 10108 39732 10164
rect 40012 9660 40068 9716
rect 41020 12738 41076 12740
rect 41020 12686 41022 12738
rect 41022 12686 41074 12738
rect 41074 12686 41076 12738
rect 41020 12684 41076 12686
rect 41356 12796 41412 12852
rect 41916 12947 41972 12964
rect 41916 12908 41918 12947
rect 41918 12908 41970 12947
rect 41970 12908 41972 12947
rect 42364 14924 42420 14980
rect 42700 15260 42756 15316
rect 43260 16380 43316 16436
rect 43036 15596 43092 15652
rect 42924 15484 42980 15540
rect 42812 15036 42868 15092
rect 43148 15372 43204 15428
rect 43036 14924 43092 14980
rect 44322 20018 44378 20020
rect 44322 19966 44324 20018
rect 44324 19966 44376 20018
rect 44376 19966 44378 20018
rect 44322 19964 44378 19966
rect 44996 19852 45052 19908
rect 44716 19628 44772 19684
rect 45444 19404 45500 19460
rect 47348 21474 47404 21476
rect 47348 21422 47350 21474
rect 47350 21422 47402 21474
rect 47402 21422 47404 21474
rect 47348 21420 47404 21422
rect 47740 21420 47796 21476
rect 47852 21532 47908 21588
rect 46844 20412 46900 20468
rect 46620 20300 46676 20356
rect 46956 20188 47012 20244
rect 47740 20802 47796 20804
rect 47740 20750 47742 20802
rect 47742 20750 47794 20802
rect 47794 20750 47796 20802
rect 47740 20748 47796 20750
rect 48636 23154 48692 23156
rect 48636 23102 48638 23154
rect 48638 23102 48690 23154
rect 48690 23102 48692 23154
rect 48636 23100 48692 23102
rect 48524 21420 48580 21476
rect 48636 21308 48692 21364
rect 47068 20018 47124 20020
rect 47068 19966 47070 20018
rect 47070 19966 47122 20018
rect 47122 19966 47124 20018
rect 47068 19964 47124 19966
rect 46956 19740 47012 19796
rect 46396 19234 46452 19236
rect 46396 19182 46398 19234
rect 46398 19182 46450 19234
rect 46450 19182 46452 19234
rect 46396 19180 46452 19182
rect 44044 18060 44100 18116
rect 43820 17651 43876 17668
rect 43820 17612 43822 17651
rect 43822 17612 43874 17651
rect 43874 17612 43876 17651
rect 44268 16882 44324 16884
rect 44268 16830 44270 16882
rect 44270 16830 44322 16882
rect 44322 16830 44324 16882
rect 44268 16828 44324 16830
rect 44548 16882 44604 16884
rect 44548 16830 44550 16882
rect 44550 16830 44602 16882
rect 44602 16830 44604 16882
rect 44548 16828 44604 16830
rect 44044 16380 44100 16436
rect 44940 16380 44996 16436
rect 43708 16156 43764 16212
rect 43372 15484 43428 15540
rect 43484 15260 43540 15316
rect 44212 16210 44268 16212
rect 44212 16158 44214 16210
rect 44214 16158 44266 16210
rect 44266 16158 44268 16210
rect 44212 16156 44268 16158
rect 43820 15484 43876 15540
rect 44716 15538 44772 15540
rect 44716 15486 44718 15538
rect 44718 15486 44770 15538
rect 44770 15486 44772 15538
rect 44716 15484 44772 15486
rect 43484 14924 43540 14980
rect 41692 12684 41748 12740
rect 41916 12124 41972 12180
rect 41412 12066 41468 12068
rect 41412 12014 41414 12066
rect 41414 12014 41466 12066
rect 41466 12014 41468 12066
rect 41412 12012 41468 12014
rect 41020 11676 41076 11732
rect 40908 10498 40964 10500
rect 40908 10446 40910 10498
rect 40910 10446 40962 10498
rect 40962 10446 40964 10498
rect 40908 10444 40964 10446
rect 41244 10610 41300 10612
rect 41244 10558 41246 10610
rect 41246 10558 41298 10610
rect 41298 10558 41300 10610
rect 41244 10556 41300 10558
rect 41020 10108 41076 10164
rect 40292 9938 40348 9940
rect 40292 9886 40294 9938
rect 40294 9886 40346 9938
rect 40346 9886 40348 9938
rect 40292 9884 40348 9886
rect 40124 9212 40180 9268
rect 41020 9826 41076 9828
rect 41020 9774 41022 9826
rect 41022 9774 41074 9826
rect 41074 9774 41076 9826
rect 41020 9772 41076 9774
rect 42140 12012 42196 12068
rect 42588 13468 42644 13524
rect 42756 12850 42812 12852
rect 42756 12798 42758 12850
rect 42758 12798 42810 12850
rect 42810 12798 42812 12850
rect 42756 12796 42812 12798
rect 42588 12236 42644 12292
rect 42364 11788 42420 11844
rect 43596 13468 43652 13524
rect 44828 14364 44884 14420
rect 44828 13692 44884 13748
rect 43932 13020 43988 13076
rect 43820 12796 43876 12852
rect 43260 12236 43316 12292
rect 42812 11900 42868 11956
rect 43372 11900 43428 11956
rect 42476 11116 42532 11172
rect 42364 10610 42420 10612
rect 42364 10558 42366 10610
rect 42366 10558 42418 10610
rect 42418 10558 42420 10610
rect 42364 10556 42420 10558
rect 41916 9884 41972 9940
rect 40852 9660 40908 9716
rect 41580 9548 41636 9604
rect 40572 9100 40628 9156
rect 41132 9212 41188 9268
rect 39788 9042 39844 9044
rect 39788 8990 39790 9042
rect 39790 8990 39842 9042
rect 39842 8990 39844 9042
rect 39788 8988 39844 8990
rect 39004 8258 39060 8260
rect 39004 8206 39006 8258
rect 39006 8206 39058 8258
rect 39058 8206 39060 8258
rect 39004 8204 39060 8206
rect 37996 3612 38052 3668
rect 38892 7084 38948 7140
rect 39172 7362 39228 7364
rect 39172 7310 39174 7362
rect 39174 7310 39226 7362
rect 39226 7310 39228 7362
rect 39172 7308 39228 7310
rect 39228 6860 39284 6916
rect 39004 6412 39060 6468
rect 39116 6748 39172 6804
rect 39788 8092 39844 8148
rect 40236 9042 40292 9044
rect 40236 8990 40238 9042
rect 40238 8990 40290 9042
rect 40290 8990 40292 9042
rect 40236 8988 40292 8990
rect 39900 7196 39956 7252
rect 39564 7084 39620 7140
rect 39340 6636 39396 6692
rect 41244 7196 41300 7252
rect 42252 9602 42308 9604
rect 42252 9550 42254 9602
rect 42254 9550 42306 9602
rect 42306 9550 42308 9602
rect 42252 9548 42308 9550
rect 42868 9996 42924 10052
rect 42476 9548 42532 9604
rect 42868 9436 42924 9492
rect 43932 12178 43988 12180
rect 43932 12126 43934 12178
rect 43934 12126 43986 12178
rect 43986 12126 43988 12178
rect 43932 12124 43988 12126
rect 43820 11788 43876 11844
rect 43708 10556 43764 10612
rect 44268 12796 44324 12852
rect 44940 13020 44996 13076
rect 44604 11788 44660 11844
rect 44380 10556 44436 10612
rect 44940 11788 44996 11844
rect 44716 11676 44772 11732
rect 43316 9826 43372 9828
rect 43316 9774 43318 9826
rect 43318 9774 43370 9826
rect 43370 9774 43372 9826
rect 43316 9772 43372 9774
rect 43148 9100 43204 9156
rect 44156 9884 44212 9940
rect 43260 9548 43316 9604
rect 43036 8370 43092 8372
rect 43036 8318 43038 8370
rect 43038 8318 43090 8370
rect 43090 8318 43092 8370
rect 43036 8316 43092 8318
rect 43036 7308 43092 7364
rect 40460 6802 40516 6804
rect 40460 6750 40462 6802
rect 40462 6750 40514 6802
rect 40514 6750 40516 6802
rect 40460 6748 40516 6750
rect 40348 6636 40404 6692
rect 41244 6690 41300 6692
rect 41244 6638 41246 6690
rect 41246 6638 41298 6690
rect 41298 6638 41300 6690
rect 41244 6636 41300 6638
rect 39228 5964 39284 6020
rect 39900 5964 39956 6020
rect 41356 6524 41412 6580
rect 39452 5628 39508 5684
rect 41356 5628 41412 5684
rect 38892 5180 38948 5236
rect 39340 5234 39396 5236
rect 39340 5182 39342 5234
rect 39342 5182 39394 5234
rect 39394 5182 39396 5234
rect 39340 5180 39396 5182
rect 39452 5068 39508 5124
rect 39004 4844 39060 4900
rect 38668 3500 38724 3556
rect 36988 3388 37044 3444
rect 39228 4396 39284 4452
rect 39116 4226 39172 4228
rect 39116 4174 39118 4226
rect 39118 4174 39170 4226
rect 39170 4174 39172 4226
rect 39116 4172 39172 4174
rect 41244 5122 41300 5124
rect 41244 5070 41246 5122
rect 41246 5070 41298 5122
rect 41298 5070 41300 5122
rect 41244 5068 41300 5070
rect 39788 4620 39844 4676
rect 40124 4338 40180 4340
rect 40124 4286 40126 4338
rect 40126 4286 40178 4338
rect 40178 4286 40180 4338
rect 40124 4284 40180 4286
rect 43484 9154 43540 9156
rect 43484 9102 43486 9154
rect 43486 9102 43538 9154
rect 43538 9102 43540 9154
rect 43484 9100 43540 9102
rect 43372 8258 43428 8260
rect 43372 8206 43374 8258
rect 43374 8206 43426 8258
rect 43426 8206 43428 8258
rect 43372 8204 43428 8206
rect 43820 9100 43876 9156
rect 44156 9660 44212 9716
rect 43988 9042 44044 9044
rect 43988 8990 43990 9042
rect 43990 8990 44042 9042
rect 44042 8990 44044 9042
rect 43988 8988 44044 8990
rect 43596 8204 43652 8260
rect 43820 8428 43876 8484
rect 43708 7532 43764 7588
rect 44268 9100 44324 9156
rect 44492 10498 44548 10500
rect 44492 10446 44494 10498
rect 44494 10446 44546 10498
rect 44546 10446 44548 10498
rect 44492 10444 44548 10446
rect 44716 10332 44772 10388
rect 44716 9884 44772 9940
rect 45612 18226 45668 18228
rect 45612 18174 45614 18226
rect 45614 18174 45666 18226
rect 45666 18174 45668 18226
rect 45612 18172 45668 18174
rect 45276 17666 45332 17668
rect 45276 17614 45278 17666
rect 45278 17614 45330 17666
rect 45330 17614 45332 17666
rect 45276 17612 45332 17614
rect 45948 17388 46004 17444
rect 45276 16882 45332 16884
rect 45276 16830 45278 16882
rect 45278 16830 45330 16882
rect 45330 16830 45332 16882
rect 45276 16828 45332 16830
rect 46452 18450 46508 18452
rect 46452 18398 46454 18450
rect 46454 18398 46506 18450
rect 46506 18398 46508 18450
rect 46452 18396 46508 18398
rect 46620 17666 46676 17668
rect 46620 17614 46622 17666
rect 46622 17614 46674 17666
rect 46674 17614 46676 17666
rect 46620 17612 46676 17614
rect 45724 16156 45780 16212
rect 46396 15314 46452 15316
rect 46396 15262 46398 15314
rect 46398 15262 46450 15314
rect 46450 15262 46452 15314
rect 46396 15260 46452 15262
rect 45183 14364 45239 14420
rect 46452 13522 46508 13524
rect 46452 13470 46454 13522
rect 46454 13470 46506 13522
rect 46506 13470 46508 13522
rect 46452 13468 46508 13470
rect 45500 12962 45556 12964
rect 45500 12910 45502 12962
rect 45502 12910 45554 12962
rect 45554 12910 45556 12962
rect 45500 12908 45556 12910
rect 48300 20300 48356 20356
rect 47292 19180 47348 19236
rect 47516 18450 47572 18452
rect 47516 18398 47518 18450
rect 47518 18398 47570 18450
rect 47570 18398 47572 18450
rect 47516 18396 47572 18398
rect 48636 20018 48692 20020
rect 48636 19966 48638 20018
rect 48638 19966 48690 20018
rect 48690 19966 48692 20018
rect 48636 19964 48692 19966
rect 48972 23042 49028 23044
rect 48972 22990 48974 23042
rect 48974 22990 49026 23042
rect 49026 22990 49028 23042
rect 48972 22988 49028 22990
rect 49420 23324 49476 23380
rect 48860 21644 48916 21700
rect 48860 21308 48916 21364
rect 48972 20748 49028 20804
rect 49308 20412 49364 20468
rect 48636 19292 48692 19348
rect 49644 34076 49700 34132
rect 49644 31836 49700 31892
rect 49532 19404 49588 19460
rect 49084 19346 49140 19348
rect 49084 19294 49086 19346
rect 49086 19294 49138 19346
rect 49138 19294 49140 19346
rect 49084 19292 49140 19294
rect 49308 19180 49364 19236
rect 48972 17836 49028 17892
rect 47068 16882 47124 16884
rect 47068 16830 47070 16882
rect 47070 16830 47122 16882
rect 47122 16830 47124 16882
rect 47068 16828 47124 16830
rect 49420 19068 49476 19124
rect 46732 15148 46788 15204
rect 47180 15820 47236 15876
rect 46284 11788 46340 11844
rect 46172 11676 46228 11732
rect 46732 12066 46788 12068
rect 46732 12014 46734 12066
rect 46734 12014 46786 12066
rect 46786 12014 46788 12066
rect 46732 12012 46788 12014
rect 45500 9996 45556 10052
rect 44996 9602 45052 9604
rect 44996 9550 44998 9602
rect 44998 9550 45050 9602
rect 45050 9550 45052 9602
rect 44996 9548 45052 9550
rect 43260 6860 43316 6916
rect 44380 7980 44436 8036
rect 42588 6188 42644 6244
rect 41580 5628 41636 5684
rect 40572 3442 40628 3444
rect 40572 3390 40574 3442
rect 40574 3390 40626 3442
rect 40626 3390 40628 3442
rect 40572 3388 40628 3390
rect 41916 5292 41972 5348
rect 41804 3724 41860 3780
rect 42028 4396 42084 4452
rect 43372 6076 43428 6132
rect 43708 5964 43764 6020
rect 43484 5852 43540 5908
rect 43484 5180 43540 5236
rect 43036 4898 43092 4900
rect 43036 4846 43038 4898
rect 43038 4846 43090 4898
rect 43090 4846 43092 4898
rect 43036 4844 43092 4846
rect 42364 4732 42420 4788
rect 42700 3778 42756 3780
rect 42700 3726 42702 3778
rect 42702 3726 42754 3778
rect 42754 3726 42756 3778
rect 42700 3724 42756 3726
rect 43820 4060 43876 4116
rect 44716 8764 44772 8820
rect 44828 8316 44884 8372
rect 44604 8092 44660 8148
rect 45276 8230 45332 8260
rect 45052 7980 45108 8036
rect 45276 8204 45278 8230
rect 45278 8204 45330 8230
rect 45330 8204 45332 8230
rect 45612 9772 45668 9828
rect 46620 11340 46676 11396
rect 46844 10668 46900 10724
rect 46060 10386 46116 10388
rect 46060 10334 46062 10386
rect 46062 10334 46114 10386
rect 46114 10334 46116 10386
rect 46060 10332 46116 10334
rect 46060 9772 46116 9828
rect 46172 10108 46228 10164
rect 47348 15314 47404 15316
rect 47348 15262 47350 15314
rect 47350 15262 47402 15314
rect 47402 15262 47404 15314
rect 47348 15260 47404 15262
rect 48076 15874 48132 15876
rect 48076 15822 48078 15874
rect 48078 15822 48130 15874
rect 48130 15822 48132 15874
rect 48076 15820 48132 15822
rect 47628 15484 47684 15540
rect 47292 14812 47348 14868
rect 47740 14924 47796 14980
rect 47628 14812 47684 14868
rect 48076 14812 48132 14868
rect 48860 14924 48916 14980
rect 48636 14812 48692 14868
rect 47852 13746 47908 13748
rect 47852 13694 47854 13746
rect 47854 13694 47906 13746
rect 47906 13694 47908 13746
rect 47852 13692 47908 13694
rect 47180 12796 47236 12852
rect 48300 13692 48356 13748
rect 45500 8092 45556 8148
rect 45500 7756 45556 7812
rect 45276 7532 45332 7588
rect 44492 7420 44548 7476
rect 44548 7250 44604 7252
rect 44548 7198 44550 7250
rect 44550 7198 44602 7250
rect 44602 7198 44604 7250
rect 44548 7196 44604 7198
rect 44604 6524 44660 6580
rect 44100 6188 44156 6244
rect 43932 3948 43988 4004
rect 44044 5404 44100 5460
rect 43764 3554 43820 3556
rect 43764 3502 43766 3554
rect 43766 3502 43818 3554
rect 43818 3502 43820 3554
rect 43764 3500 43820 3502
rect 44156 4844 44212 4900
rect 45500 6748 45556 6804
rect 46284 8092 46340 8148
rect 45724 7756 45780 7812
rect 45724 7308 45780 7364
rect 44380 5964 44436 6020
rect 44604 5964 44660 6020
rect 44492 5852 44548 5908
rect 44268 3388 44324 3444
rect 44828 5882 44830 5908
rect 44830 5882 44882 5908
rect 44882 5882 44884 5908
rect 44828 5852 44884 5882
rect 44940 5404 44996 5460
rect 44940 5234 44996 5236
rect 44940 5182 44942 5234
rect 44942 5182 44994 5234
rect 44994 5182 44996 5234
rect 44940 5180 44996 5182
rect 44716 4956 44772 5012
rect 45388 6188 45444 6244
rect 45500 6412 45556 6468
rect 45164 5964 45220 6020
rect 45388 5180 45444 5236
rect 45500 4732 45556 4788
rect 45612 5292 45668 5348
rect 46116 6466 46172 6468
rect 46116 6414 46118 6466
rect 46118 6414 46170 6466
rect 46170 6414 46172 6466
rect 46116 6412 46172 6414
rect 45836 5964 45892 6020
rect 46620 7756 46676 7812
rect 46284 5516 46340 5572
rect 46396 6748 46452 6804
rect 46620 6578 46676 6580
rect 46620 6526 46622 6578
rect 46622 6526 46674 6578
rect 46674 6526 46676 6578
rect 46620 6524 46676 6526
rect 48860 13746 48916 13748
rect 48860 13694 48862 13746
rect 48862 13694 48914 13746
rect 48914 13694 48916 13746
rect 48860 13692 48916 13694
rect 49084 14812 49140 14868
rect 49140 13634 49196 13636
rect 49140 13582 49142 13634
rect 49142 13582 49194 13634
rect 49194 13582 49196 13634
rect 49140 13580 49196 13582
rect 47404 12012 47460 12068
rect 48412 11788 48468 11844
rect 47964 11394 48020 11396
rect 47964 11342 47966 11394
rect 47966 11342 48018 11394
rect 48018 11342 48020 11394
rect 47964 11340 48020 11342
rect 47404 10585 47406 10612
rect 47406 10585 47458 10612
rect 47458 10585 47460 10612
rect 47404 10556 47460 10585
rect 47404 10332 47460 10388
rect 48244 10610 48300 10612
rect 48244 10558 48246 10610
rect 48246 10558 48298 10610
rect 48298 10558 48300 10610
rect 48244 10556 48300 10558
rect 48188 9826 48244 9828
rect 48188 9774 48190 9826
rect 48190 9774 48242 9826
rect 48242 9774 48244 9826
rect 48188 9772 48244 9774
rect 48524 10444 48580 10500
rect 48636 10108 48692 10164
rect 48636 8764 48692 8820
rect 47068 6636 47124 6692
rect 46956 6300 47012 6356
rect 47180 6076 47236 6132
rect 47292 7196 47348 7252
rect 46956 5516 47012 5572
rect 45724 5180 45780 5236
rect 46620 5180 46676 5236
rect 45948 3948 46004 4004
rect 45836 3836 45892 3892
rect 45164 3388 45220 3444
rect 45332 3442 45388 3444
rect 45332 3390 45334 3442
rect 45334 3390 45386 3442
rect 45386 3390 45388 3442
rect 45332 3388 45388 3390
rect 44716 2044 44772 2100
rect 46508 3724 46564 3780
rect 46732 4732 46788 4788
rect 46844 4172 46900 4228
rect 48300 6636 48356 6692
rect 47852 6412 47908 6468
rect 47740 6076 47796 6132
rect 47516 5906 47572 5908
rect 47516 5854 47518 5906
rect 47518 5854 47570 5906
rect 47570 5854 47572 5906
rect 47516 5852 47572 5854
rect 47068 5068 47124 5124
rect 47292 5068 47348 5124
rect 47628 5122 47684 5124
rect 47628 5070 47630 5122
rect 47630 5070 47682 5122
rect 47682 5070 47684 5122
rect 47628 5068 47684 5070
rect 48748 8204 48804 8260
rect 48972 10386 49028 10388
rect 48972 10334 48974 10386
rect 48974 10334 49026 10386
rect 49026 10334 49028 10386
rect 48972 10332 49028 10334
rect 49308 9772 49364 9828
rect 48972 8428 49028 8484
rect 48860 7868 48916 7924
rect 48412 6076 48468 6132
rect 47964 5180 48020 5236
rect 48188 5180 48244 5236
rect 48300 5068 48356 5124
rect 48412 5292 48468 5348
rect 48524 4956 48580 5012
rect 47628 3666 47684 3668
rect 47628 3614 47630 3666
rect 47630 3614 47682 3666
rect 47682 3614 47684 3666
rect 47628 3612 47684 3614
rect 46732 3388 46788 3444
rect 46620 3330 46676 3332
rect 46620 3278 46622 3330
rect 46622 3278 46674 3330
rect 46674 3278 46676 3330
rect 46620 3276 46676 3278
rect 48300 3778 48356 3780
rect 48300 3726 48302 3778
rect 48302 3726 48354 3778
rect 48354 3726 48356 3778
rect 48300 3724 48356 3726
rect 47964 3554 48020 3556
rect 47964 3502 47966 3554
rect 47966 3502 48018 3554
rect 48018 3502 48020 3554
rect 47964 3500 48020 3502
rect 49084 5852 49140 5908
rect 49196 7868 49252 7924
rect 49308 6690 49364 6692
rect 49308 6638 49310 6690
rect 49310 6638 49362 6690
rect 49362 6638 49364 6690
rect 49308 6636 49364 6638
rect 49196 6188 49252 6244
rect 49196 5180 49252 5236
rect 49140 4898 49196 4900
rect 49140 4846 49142 4898
rect 49142 4846 49194 4898
rect 49194 4846 49196 4898
rect 49140 4844 49196 4846
rect 48972 4172 49028 4228
<< metal3 >>
rect 50200 48916 51000 48944
rect 49298 48860 49308 48916
rect 49364 48860 51000 48916
rect 50200 48832 51000 48860
rect 5730 48300 5740 48356
rect 5796 48300 6300 48356
rect 6356 48300 6366 48356
rect 39274 48076 39284 48132
rect 39340 48076 44604 48132
rect 44660 48076 47292 48132
rect 47348 48076 47358 48132
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 38826 47628 38836 47684
rect 38892 47628 49308 47684
rect 49364 47628 49374 47684
rect 21074 47516 21084 47572
rect 21140 47516 22428 47572
rect 22484 47516 22494 47572
rect 32610 47516 32620 47572
rect 32676 47516 33852 47572
rect 33908 47516 33918 47572
rect 44482 47516 44492 47572
rect 44548 47516 46396 47572
rect 46452 47516 46462 47572
rect 22754 47404 22764 47460
rect 22820 47404 24892 47460
rect 24948 47404 24958 47460
rect 26618 47404 26628 47460
rect 26684 47404 29240 47460
rect 29296 47404 30492 47460
rect 30548 47404 30558 47460
rect 35186 47404 35196 47460
rect 35252 47404 38276 47460
rect 38332 47404 43708 47460
rect 43764 47404 43774 47460
rect 33954 47292 33964 47348
rect 34020 47292 38668 47348
rect 41906 47292 41916 47348
rect 41972 47292 42364 47348
rect 42420 47292 42430 47348
rect 42970 47292 42980 47348
rect 43036 47292 45724 47348
rect 45780 47292 45790 47348
rect 38612 47236 38668 47292
rect 23258 47180 23268 47236
rect 23324 47180 23884 47236
rect 23940 47180 24556 47236
rect 24612 47180 24622 47236
rect 29250 47180 29260 47236
rect 29316 47180 30212 47236
rect 30268 47180 32172 47236
rect 32228 47180 36316 47236
rect 36372 47180 36932 47236
rect 36988 47180 36998 47236
rect 38612 47180 43708 47236
rect 44258 47180 44268 47236
rect 44324 47180 46508 47236
rect 46564 47180 46574 47236
rect 47590 47180 47628 47236
rect 47684 47180 47694 47236
rect 43652 47124 43708 47180
rect 24658 47068 24668 47124
rect 24724 47068 25340 47124
rect 25396 47068 25406 47124
rect 32498 47068 32508 47124
rect 32564 47068 35420 47124
rect 35476 47068 35486 47124
rect 40562 47068 40572 47124
rect 40628 47068 41972 47124
rect 43652 47068 48972 47124
rect 49028 47068 49038 47124
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 41916 47012 41972 47068
rect 31126 46956 31164 47012
rect 31220 46956 31230 47012
rect 41916 46956 43708 47012
rect 43764 46956 45836 47012
rect 45892 46956 45902 47012
rect 43810 46844 43820 46900
rect 43876 46844 45276 46900
rect 45332 46844 45342 46900
rect 27570 46620 27580 46676
rect 27636 46620 28364 46676
rect 28420 46620 30380 46676
rect 30436 46620 32956 46676
rect 33012 46620 33022 46676
rect 40002 46620 40012 46676
rect 40068 46620 40684 46676
rect 40740 46620 40750 46676
rect 41458 46620 41468 46676
rect 41524 46620 42140 46676
rect 42196 46620 42206 46676
rect 46050 46620 46060 46676
rect 46116 46620 48636 46676
rect 48692 46620 48702 46676
rect 13570 46508 13580 46564
rect 13636 46508 16716 46564
rect 16772 46508 17836 46564
rect 17892 46508 17902 46564
rect 36642 46508 36652 46564
rect 36708 46508 42364 46564
rect 42420 46508 42430 46564
rect 46162 46508 46172 46564
rect 46228 46508 48972 46564
rect 49028 46508 49038 46564
rect 12338 46396 12348 46452
rect 12404 46396 13748 46452
rect 13804 46396 13814 46452
rect 17434 46396 17444 46452
rect 17500 46396 18172 46452
rect 18228 46396 18238 46452
rect 30874 46396 30884 46452
rect 30940 46396 31500 46452
rect 31556 46396 31566 46452
rect 46274 46396 46284 46452
rect 46340 46396 48076 46452
rect 48132 46396 48142 46452
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 11106 45948 11116 46004
rect 11172 45948 13356 46004
rect 13412 45948 13692 46004
rect 13748 45948 13758 46004
rect 30818 45948 30828 46004
rect 30884 45948 31164 46004
rect 31220 45948 31230 46004
rect 11442 45836 11452 45892
rect 11508 45836 12012 45892
rect 12068 45836 12078 45892
rect 26338 45836 26348 45892
rect 26404 45836 26684 45892
rect 26740 45836 27804 45892
rect 27860 45836 27870 45892
rect 30034 45836 30044 45892
rect 30100 45836 30268 45892
rect 30324 45836 32956 45892
rect 33012 45836 33516 45892
rect 33572 45836 33740 45892
rect 33796 45836 36316 45892
rect 36372 45836 36876 45892
rect 36932 45836 36942 45892
rect 41794 45836 41804 45892
rect 41860 45836 42700 45892
rect 42756 45836 42766 45892
rect 45490 45836 45500 45892
rect 45556 45836 45948 45892
rect 46004 45836 46014 45892
rect 11330 45724 11340 45780
rect 11396 45724 11676 45780
rect 11732 45724 13468 45780
rect 13524 45724 13534 45780
rect 17602 45724 17612 45780
rect 17668 45724 18396 45780
rect 18452 45724 18462 45780
rect 34850 45724 34860 45780
rect 34916 45724 36092 45780
rect 36148 45724 36158 45780
rect 40450 45724 40460 45780
rect 40516 45724 41356 45780
rect 41412 45724 46172 45780
rect 46228 45724 46238 45780
rect 26674 45612 26684 45668
rect 26740 45612 27356 45668
rect 27412 45612 27422 45668
rect 31714 45612 31724 45668
rect 31780 45612 32060 45668
rect 32116 45612 32732 45668
rect 32788 45612 32798 45668
rect 42130 45612 42140 45668
rect 42196 45612 43576 45668
rect 43632 45612 43642 45668
rect 44034 45500 44044 45556
rect 44100 45500 47180 45556
rect 47236 45500 47246 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 14690 45388 14700 45444
rect 14756 45388 18172 45444
rect 18228 45388 18238 45444
rect 42354 45388 42364 45444
rect 42420 45388 44716 45444
rect 44772 45388 44782 45444
rect 17938 45276 17948 45332
rect 18004 45276 18396 45332
rect 18452 45276 20188 45332
rect 20244 45276 21308 45332
rect 21364 45276 21374 45332
rect 22754 45276 22764 45332
rect 22820 45276 22830 45332
rect 36474 45276 36484 45332
rect 36540 45276 36876 45332
rect 36932 45276 38332 45332
rect 38388 45276 38398 45332
rect 39946 45276 39956 45332
rect 40012 45276 44492 45332
rect 44548 45276 45276 45332
rect 45332 45276 47292 45332
rect 47348 45276 47358 45332
rect 48636 45276 49084 45332
rect 49140 45276 49150 45332
rect 13570 45164 13580 45220
rect 13636 45164 15596 45220
rect 15652 45164 15662 45220
rect 17714 45052 17724 45108
rect 17780 45052 17948 45108
rect 18004 45052 21196 45108
rect 21252 45052 21262 45108
rect 22764 44772 22820 45276
rect 48636 45220 48692 45276
rect 36306 45164 36316 45220
rect 36372 45164 38220 45220
rect 38276 45164 38286 45220
rect 42466 45164 42476 45220
rect 42532 45164 43148 45220
rect 43204 45164 43214 45220
rect 47180 45164 48636 45220
rect 48692 45164 48702 45220
rect 47180 45108 47236 45164
rect 23874 45052 23884 45108
rect 23940 45052 25228 45108
rect 25284 45052 25294 45108
rect 26226 45052 26236 45108
rect 26292 45052 30604 45108
rect 30660 45052 30670 45108
rect 31042 45052 31052 45108
rect 31108 45052 32228 45108
rect 32284 45052 32294 45108
rect 37034 45052 37044 45108
rect 37100 45052 38556 45108
rect 38612 45052 38622 45108
rect 40226 45052 40236 45108
rect 40292 45052 40908 45108
rect 40964 45052 40974 45108
rect 41774 45052 41784 45108
rect 41840 45052 42364 45108
rect 42420 45052 42430 45108
rect 42690 45052 42700 45108
rect 42756 45052 45724 45108
rect 45780 45052 47180 45108
rect 47236 45052 47246 45108
rect 47394 45052 47404 45108
rect 47460 45052 47964 45108
rect 48020 45052 49140 45108
rect 49196 45052 49206 45108
rect 25228 44996 25284 45052
rect 25228 44940 28252 44996
rect 28308 44940 28318 44996
rect 36194 44940 36204 44996
rect 36260 44940 38668 44996
rect 43586 44940 43596 44996
rect 43652 44940 46060 44996
rect 46116 44940 46126 44996
rect 36530 44828 36540 44884
rect 36596 44828 37996 44884
rect 38052 44828 38062 44884
rect 38612 44828 38668 44940
rect 38724 44828 39508 44884
rect 39564 44828 39574 44884
rect 22754 44716 22764 44772
rect 22820 44716 22830 44772
rect 28018 44716 28028 44772
rect 28084 44716 28588 44772
rect 28644 44716 29260 44772
rect 29316 44716 29326 44772
rect 32218 44716 32228 44772
rect 32284 44716 34392 44772
rect 34448 44716 34458 44772
rect 37762 44716 37772 44772
rect 37828 44716 39340 44772
rect 39396 44716 39406 44772
rect 41804 44716 46732 44772
rect 46788 44716 46798 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 16818 44604 16828 44660
rect 16884 44604 17444 44660
rect 17500 44604 17510 44660
rect 20738 44604 20748 44660
rect 20804 44604 29372 44660
rect 29428 44604 29438 44660
rect 32386 44604 32396 44660
rect 32452 44604 32844 44660
rect 32900 44604 32910 44660
rect 39666 44604 39676 44660
rect 39732 44604 41244 44660
rect 41300 44604 41310 44660
rect 41804 44548 41860 44716
rect 46834 44604 46844 44660
rect 46900 44604 48300 44660
rect 48356 44604 48366 44660
rect 50200 44576 51000 44688
rect 9090 44492 9100 44548
rect 9156 44492 10220 44548
rect 10276 44492 10286 44548
rect 40674 44492 40684 44548
rect 40740 44492 41804 44548
rect 41860 44492 41870 44548
rect 42914 44492 42924 44548
rect 42980 44492 43484 44548
rect 43540 44492 43550 44548
rect 45490 44492 45500 44548
rect 45556 44492 46396 44548
rect 46452 44492 47628 44548
rect 47684 44492 48860 44548
rect 48916 44492 48926 44548
rect 14802 44380 14812 44436
rect 14868 44380 15820 44436
rect 15876 44380 15886 44436
rect 20514 44380 20524 44436
rect 20580 44380 20748 44436
rect 20804 44380 20814 44436
rect 21522 44380 21532 44436
rect 21588 44380 21598 44436
rect 23762 44380 23772 44436
rect 23828 44380 24780 44436
rect 24836 44380 25564 44436
rect 25620 44380 25630 44436
rect 40450 44380 40460 44436
rect 40516 44380 41468 44436
rect 41524 44380 41534 44436
rect 42130 44380 42140 44436
rect 42196 44380 42812 44436
rect 42868 44380 42878 44436
rect 46162 44380 46172 44436
rect 46228 44380 46508 44436
rect 46564 44380 46574 44436
rect 21532 44324 21588 44380
rect 8754 44268 8764 44324
rect 8820 44268 9548 44324
rect 9604 44268 9884 44324
rect 9940 44268 9950 44324
rect 16930 44268 16940 44324
rect 16996 44268 18060 44324
rect 18116 44268 18126 44324
rect 18386 44268 18396 44324
rect 18452 44268 19964 44324
rect 20020 44268 21084 44324
rect 21140 44268 21150 44324
rect 21532 44268 23436 44324
rect 23492 44268 23660 44324
rect 23716 44268 25228 44324
rect 25284 44268 25294 44324
rect 28242 44268 28252 44324
rect 28308 44268 29036 44324
rect 29092 44268 29102 44324
rect 29530 44268 29540 44324
rect 29596 44268 30268 44324
rect 30324 44268 30492 44324
rect 30548 44268 30558 44324
rect 31714 44268 31724 44324
rect 31780 44268 32732 44324
rect 32788 44268 32798 44324
rect 34382 44268 34392 44324
rect 34448 44268 35196 44324
rect 35252 44268 35262 44324
rect 41234 44268 41244 44324
rect 41300 44268 43260 44324
rect 43316 44268 43326 44324
rect 44370 44268 44380 44324
rect 44436 44268 47516 44324
rect 47572 44268 47582 44324
rect 9426 44156 9436 44212
rect 9492 44156 11340 44212
rect 11396 44156 11406 44212
rect 12114 44156 12124 44212
rect 12180 44156 12684 44212
rect 12740 44156 16268 44212
rect 16324 44156 16334 44212
rect 21644 44100 21700 44268
rect 33506 44156 33516 44212
rect 33572 44156 34748 44212
rect 34804 44156 35532 44212
rect 35588 44156 37324 44212
rect 37380 44156 37390 44212
rect 45378 44156 45388 44212
rect 45444 44156 46060 44212
rect 46116 44156 46844 44212
rect 46900 44156 46910 44212
rect 7858 44044 7868 44100
rect 7924 44044 11116 44100
rect 11172 44044 11182 44100
rect 15362 44044 15372 44100
rect 15428 44044 16156 44100
rect 16212 44044 18284 44100
rect 18340 44044 18350 44100
rect 19618 44044 19628 44100
rect 19684 44044 20636 44100
rect 20692 44044 20702 44100
rect 21634 44044 21644 44100
rect 21700 44044 21710 44100
rect 27682 44044 27692 44100
rect 27748 44044 27916 44100
rect 27972 44044 29036 44100
rect 29092 44044 29102 44100
rect 43922 44044 43932 44100
rect 43988 44044 44828 44100
rect 44884 44044 44894 44100
rect 14578 43932 14588 43988
rect 14644 43932 15932 43988
rect 15988 43932 15998 43988
rect 28018 43932 28028 43988
rect 28084 43932 29148 43988
rect 29204 43932 29214 43988
rect 42924 43932 44940 43988
rect 44996 43932 45006 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 42924 43876 42980 43932
rect 18666 43820 18676 43876
rect 18732 43820 19460 43876
rect 39330 43820 39340 43876
rect 39396 43820 42924 43876
rect 42980 43820 42990 43876
rect 44370 43820 44380 43876
rect 44436 43820 45052 43876
rect 45108 43820 46508 43876
rect 46564 43820 46574 43876
rect 19404 43764 19460 43820
rect 7196 43708 7532 43764
rect 7588 43708 7598 43764
rect 11442 43708 11452 43764
rect 11508 43708 12012 43764
rect 12068 43708 12078 43764
rect 13682 43708 13692 43764
rect 13748 43708 14364 43764
rect 14420 43708 14430 43764
rect 17602 43708 17612 43764
rect 17668 43708 18396 43764
rect 18452 43708 18462 43764
rect 19404 43708 20636 43764
rect 20692 43708 23268 43764
rect 7196 43316 7252 43708
rect 23212 43652 23268 43708
rect 30940 43708 31836 43764
rect 31892 43708 31902 43764
rect 36418 43708 36428 43764
rect 36484 43708 37100 43764
rect 37156 43708 38220 43764
rect 38276 43708 38286 43764
rect 30940 43652 30996 43708
rect 13010 43596 13020 43652
rect 13076 43596 13524 43652
rect 13580 43596 13590 43652
rect 14466 43596 14476 43652
rect 14532 43596 16604 43652
rect 16660 43596 16670 43652
rect 21858 43596 21868 43652
rect 21924 43596 22204 43652
rect 22260 43596 23007 43652
rect 23063 43596 23073 43652
rect 23212 43596 25116 43652
rect 25172 43596 25182 43652
rect 30930 43596 30940 43652
rect 30996 43596 31006 43652
rect 31490 43596 31500 43652
rect 31556 43596 32956 43652
rect 33012 43596 33404 43652
rect 33460 43596 33470 43652
rect 40338 43596 40348 43652
rect 40404 43596 41692 43652
rect 41748 43596 41758 43652
rect 42690 43596 42700 43652
rect 42756 43596 45164 43652
rect 45220 43596 45230 43652
rect 10882 43484 10892 43540
rect 10948 43484 12572 43540
rect 12628 43484 12638 43540
rect 13234 43484 13244 43540
rect 13300 43484 14028 43540
rect 14084 43484 14924 43540
rect 14980 43484 16044 43540
rect 16100 43484 16110 43540
rect 16706 43484 16716 43540
rect 16772 43484 17052 43540
rect 17108 43484 17276 43540
rect 17332 43484 17342 43540
rect 21522 43484 21532 43540
rect 21588 43484 21756 43540
rect 21812 43484 21822 43540
rect 22082 43484 22092 43540
rect 22148 43484 24220 43540
rect 24276 43484 24286 43540
rect 28578 43484 28588 43540
rect 28644 43484 29372 43540
rect 29428 43484 29820 43540
rect 29876 43484 29886 43540
rect 32162 43484 32172 43540
rect 32228 43484 35644 43540
rect 35700 43484 35710 43540
rect 38546 43484 38556 43540
rect 38612 43484 40460 43540
rect 40516 43484 40908 43540
rect 40964 43484 40974 43540
rect 44146 43484 44156 43540
rect 44212 43484 45948 43540
rect 46004 43484 46014 43540
rect 46722 43484 46732 43540
rect 46788 43484 47516 43540
rect 47572 43484 47582 43540
rect 11564 43428 11620 43484
rect 11554 43372 11564 43428
rect 11620 43372 11630 43428
rect 13794 43372 13804 43428
rect 13860 43372 14476 43428
rect 14532 43372 14542 43428
rect 20738 43372 20748 43428
rect 20804 43372 21028 43428
rect 21084 43372 26908 43428
rect 28130 43372 28140 43428
rect 28196 43372 28812 43428
rect 28868 43372 29148 43428
rect 29204 43372 29214 43428
rect 30538 43372 30548 43428
rect 30604 43372 33236 43428
rect 33292 43372 33302 43428
rect 34738 43372 34748 43428
rect 34804 43372 35756 43428
rect 35812 43372 35822 43428
rect 26852 43316 26908 43372
rect 7186 43260 7196 43316
rect 7252 43260 7262 43316
rect 8866 43260 8876 43316
rect 8932 43260 9996 43316
rect 10052 43260 16156 43316
rect 16212 43260 16222 43316
rect 17266 43260 17276 43316
rect 17332 43260 17780 43316
rect 17836 43260 17846 43316
rect 26852 43260 27468 43316
rect 27524 43260 28252 43316
rect 28308 43260 28318 43316
rect 34962 43260 34972 43316
rect 35028 43260 35532 43316
rect 35588 43260 37212 43316
rect 37268 43260 37278 43316
rect 42242 43260 42252 43316
rect 42308 43260 43372 43316
rect 43428 43260 43438 43316
rect 45938 43260 45948 43316
rect 46004 43260 46956 43316
rect 47012 43260 47022 43316
rect 27906 43148 27916 43204
rect 27972 43148 28700 43204
rect 28756 43148 28924 43204
rect 28980 43148 28990 43204
rect 32050 43148 32060 43204
rect 32116 43148 33068 43204
rect 33124 43148 33134 43204
rect 38612 43148 39228 43204
rect 39284 43148 43708 43204
rect 47842 43148 47852 43204
rect 47908 43148 48412 43204
rect 48468 43148 48478 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 7429 43036 7439 43092
rect 7495 43036 13412 43092
rect 13468 43036 13478 43092
rect 18386 43036 18396 43092
rect 18452 43036 18956 43092
rect 19012 43036 19022 43092
rect 29530 43036 29540 43092
rect 29596 43036 31052 43092
rect 31108 43036 33516 43092
rect 33572 43036 33582 43092
rect 38612 42980 38668 43148
rect 43652 43092 43708 43148
rect 42802 43036 42812 43092
rect 42868 43036 43036 43092
rect 43092 43036 43102 43092
rect 43652 43036 44716 43092
rect 44772 43036 44782 43092
rect 47170 43036 47180 43092
rect 47236 43036 47964 43092
rect 48020 43036 48030 43092
rect 12562 42924 12572 42980
rect 12628 42924 12908 42980
rect 12964 42924 12974 42980
rect 25442 42924 25452 42980
rect 25508 42924 26012 42980
rect 26068 42924 26078 42980
rect 31154 42924 31164 42980
rect 31220 42924 31836 42980
rect 31892 42924 31902 42980
rect 32610 42924 32620 42980
rect 32676 42924 33180 42980
rect 33236 42924 33246 42980
rect 37538 42924 37548 42980
rect 37604 42924 38668 42980
rect 43698 42924 43708 42980
rect 43764 42924 44100 42980
rect 44156 42924 44166 42980
rect 30706 42812 30716 42868
rect 30772 42812 31388 42868
rect 31444 42812 31454 42868
rect 32778 42812 32788 42868
rect 32844 42812 33796 42868
rect 33852 42812 33862 42868
rect 34458 42812 34468 42868
rect 34524 42812 35420 42868
rect 35476 42812 35486 42868
rect 35634 42812 35644 42868
rect 35700 42812 36988 42868
rect 37044 42812 37054 42868
rect 43530 42812 43540 42868
rect 43596 42812 45388 42868
rect 45444 42812 45454 42868
rect 35644 42756 35700 42812
rect 12198 42700 12236 42756
rect 12292 42700 12796 42756
rect 12852 42700 12862 42756
rect 13010 42700 13020 42756
rect 13076 42700 13580 42756
rect 13636 42700 13646 42756
rect 16034 42700 16044 42756
rect 16100 42700 17948 42756
rect 18004 42700 18014 42756
rect 20626 42700 20636 42756
rect 20692 42700 21196 42756
rect 21252 42700 21262 42756
rect 25778 42700 25788 42756
rect 25844 42700 27412 42756
rect 27468 42700 27478 42756
rect 27682 42700 27692 42756
rect 27748 42700 29260 42756
rect 29316 42700 29326 42756
rect 32946 42700 32956 42756
rect 33012 42700 34076 42756
rect 34132 42700 34142 42756
rect 34524 42700 35700 42756
rect 38098 42700 38108 42756
rect 38164 42700 38668 42756
rect 38724 42700 38734 42756
rect 42858 42700 42868 42756
rect 42924 42700 43820 42756
rect 43876 42700 43886 42756
rect 34524 42644 34580 42700
rect 11666 42588 11676 42644
rect 11732 42588 12124 42644
rect 12180 42588 12190 42644
rect 13458 42588 13468 42644
rect 13524 42588 14476 42644
rect 14532 42588 14542 42644
rect 15362 42588 15372 42644
rect 15428 42588 16268 42644
rect 16324 42588 18060 42644
rect 18116 42588 18126 42644
rect 24938 42588 24948 42644
rect 25004 42588 29820 42644
rect 29876 42588 30716 42644
rect 30772 42588 30782 42644
rect 34514 42588 34524 42644
rect 34580 42588 34590 42644
rect 35018 42588 35028 42644
rect 35084 42588 36092 42644
rect 36148 42588 36158 42644
rect 10770 42476 10780 42532
rect 10836 42476 12236 42532
rect 12292 42476 12302 42532
rect 17490 42476 17500 42532
rect 17556 42476 21364 42532
rect 21420 42476 21430 42532
rect 31826 42476 31836 42532
rect 31892 42476 32508 42532
rect 32564 42476 35308 42532
rect 35364 42476 35374 42532
rect 40870 42476 40908 42532
rect 40964 42476 40974 42532
rect 11218 42364 11228 42420
rect 11284 42364 11452 42420
rect 11508 42364 11518 42420
rect 34738 42364 34748 42420
rect 34804 42364 34972 42420
rect 35028 42364 35038 42420
rect 36082 42364 36092 42420
rect 36148 42364 36652 42420
rect 36708 42364 37324 42420
rect 37380 42364 40460 42420
rect 40516 42364 40526 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 29138 42252 29148 42308
rect 29204 42252 35252 42308
rect 35308 42252 35318 42308
rect 9538 42140 9548 42196
rect 9604 42140 9996 42196
rect 10052 42140 10062 42196
rect 10322 42140 10332 42196
rect 10388 42140 11228 42196
rect 11284 42140 11294 42196
rect 20066 42140 20076 42196
rect 20132 42140 20636 42196
rect 20692 42140 20702 42196
rect 21634 42140 21644 42196
rect 21700 42140 22428 42196
rect 22484 42140 22494 42196
rect 42858 42140 42868 42196
rect 42924 42140 43484 42196
rect 43540 42140 43550 42196
rect 35970 42028 35980 42084
rect 36036 42028 36540 42084
rect 36596 42028 36606 42084
rect 40338 42028 40348 42084
rect 40404 42028 41784 42084
rect 41840 42028 41850 42084
rect 6402 41916 6412 41972
rect 6468 41916 6916 41972
rect 6972 41916 7756 41972
rect 7812 41916 7822 41972
rect 8306 41916 8316 41972
rect 8372 41916 9660 41972
rect 9716 41916 9726 41972
rect 12334 41916 12344 41972
rect 12400 41916 13692 41972
rect 13748 41916 13758 41972
rect 13906 41916 13916 41972
rect 13972 41916 15372 41972
rect 15428 41916 15438 41972
rect 16426 41916 16436 41972
rect 16492 41916 18620 41972
rect 18676 41916 18686 41972
rect 22754 41916 22764 41972
rect 22820 41916 24332 41972
rect 24388 41916 25228 41972
rect 25284 41916 25294 41972
rect 25890 41916 25900 41972
rect 25956 41916 26460 41972
rect 26516 41916 26526 41972
rect 30258 41916 30268 41972
rect 30324 41916 30828 41972
rect 30884 41916 31052 41972
rect 31108 41916 31118 41972
rect 36194 41916 36204 41972
rect 36260 41916 37436 41972
rect 37492 41916 37502 41972
rect 40226 41916 40236 41972
rect 40292 41916 41580 41972
rect 41636 41916 41646 41972
rect 42858 41916 42868 41972
rect 42924 41916 43820 41972
rect 43876 41916 43886 41972
rect 44258 41916 44268 41972
rect 44324 41916 45164 41972
rect 45220 41916 45230 41972
rect 46386 41916 46396 41972
rect 46452 41916 47964 41972
rect 48020 41916 48300 41972
rect 48356 41916 49308 41972
rect 49364 41916 49374 41972
rect 6626 41804 6636 41860
rect 6692 41804 8204 41860
rect 8260 41804 8270 41860
rect 10714 41804 10724 41860
rect 10780 41804 12572 41860
rect 12628 41804 13468 41860
rect 13524 41804 13534 41860
rect 15698 41804 15708 41860
rect 15764 41804 17500 41860
rect 17556 41804 17566 41860
rect 22530 41804 22540 41860
rect 22596 41804 23212 41860
rect 23268 41804 23278 41860
rect 28466 41804 28476 41860
rect 28532 41804 28980 41860
rect 29036 41804 29046 41860
rect 35242 41804 35252 41860
rect 35308 41804 35644 41860
rect 35700 41804 35710 41860
rect 35858 41804 35868 41860
rect 35924 41804 39340 41860
rect 39396 41804 39406 41860
rect 7410 41692 7420 41748
rect 7476 41692 8316 41748
rect 8372 41692 8382 41748
rect 8586 41692 8596 41748
rect 8652 41692 10332 41748
rect 10388 41692 10398 41748
rect 16146 41692 16156 41748
rect 16212 41692 18228 41748
rect 18284 41692 18294 41748
rect 23930 41692 23940 41748
rect 23996 41692 24556 41748
rect 24612 41692 24622 41748
rect 25386 41692 25396 41748
rect 25452 41692 27916 41748
rect 27972 41692 27982 41748
rect 30706 41692 30716 41748
rect 30772 41692 31724 41748
rect 31780 41692 31790 41748
rect 34514 41692 34524 41748
rect 34580 41692 36876 41748
rect 36932 41692 36942 41748
rect 48962 41692 48972 41748
rect 49028 41692 49420 41748
rect 49476 41692 49486 41748
rect 15586 41580 15596 41636
rect 15652 41580 16604 41636
rect 16660 41580 17388 41636
rect 17444 41580 17454 41636
rect 31042 41580 31052 41636
rect 31108 41580 32004 41636
rect 32060 41580 32620 41636
rect 32676 41580 32686 41636
rect 35634 41580 35644 41636
rect 35700 41580 36988 41636
rect 37044 41580 38220 41636
rect 38276 41580 38286 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 26226 41468 26236 41524
rect 26292 41468 26302 41524
rect 36418 41468 36428 41524
rect 36484 41468 36494 41524
rect 44930 41468 44940 41524
rect 44996 41468 45500 41524
rect 45556 41468 46956 41524
rect 47012 41468 47022 41524
rect 48290 41468 48300 41524
rect 48356 41468 48524 41524
rect 48580 41468 48590 41524
rect 10098 41356 10108 41412
rect 10164 41356 10612 41412
rect 10668 41356 15932 41412
rect 15988 41356 15998 41412
rect 17490 41356 17500 41412
rect 17556 41356 18788 41412
rect 18844 41356 18854 41412
rect 26236 41300 26292 41468
rect 36428 41412 36484 41468
rect 28242 41356 28252 41412
rect 28308 41356 36484 41412
rect 38322 41356 38332 41412
rect 38388 41356 39116 41412
rect 39172 41356 39182 41412
rect 5618 41244 5628 41300
rect 5684 41244 6300 41300
rect 6356 41244 6366 41300
rect 21186 41244 21196 41300
rect 21252 41244 21756 41300
rect 21812 41244 23548 41300
rect 23604 41244 26292 41300
rect 29530 41244 29540 41300
rect 29596 41244 30156 41300
rect 30212 41244 30222 41300
rect 34066 41244 34076 41300
rect 34132 41244 35196 41300
rect 35252 41244 35262 41300
rect 44482 41244 44492 41300
rect 44548 41244 45500 41300
rect 45556 41244 45566 41300
rect 9874 41132 9884 41188
rect 9940 41132 10892 41188
rect 10948 41132 10958 41188
rect 11106 41132 11116 41188
rect 11172 41132 11340 41188
rect 11396 41132 11676 41188
rect 11732 41132 11742 41188
rect 12542 41132 12552 41188
rect 12608 41132 13804 41188
rect 13860 41132 13870 41188
rect 16482 41132 16492 41188
rect 16548 41132 17108 41188
rect 17164 41132 17174 41188
rect 20514 41132 20524 41188
rect 20580 41132 21420 41188
rect 21476 41132 21868 41188
rect 21924 41132 23324 41188
rect 23380 41132 23390 41188
rect 27906 41132 27916 41188
rect 27972 41132 29036 41188
rect 29092 41132 29102 41188
rect 29260 41132 33292 41188
rect 33348 41132 33628 41188
rect 33684 41132 33694 41188
rect 45714 41132 45724 41188
rect 45780 41132 46452 41188
rect 46508 41132 46518 41188
rect 48514 41132 48524 41188
rect 48580 41132 48748 41188
rect 48804 41132 48814 41188
rect 29260 41076 29316 41132
rect 8194 41020 8204 41076
rect 8260 41020 8652 41076
rect 8708 41020 8718 41076
rect 9034 41020 9044 41076
rect 9100 41020 15820 41076
rect 15876 41020 15886 41076
rect 23202 41020 23212 41076
rect 23268 41020 24220 41076
rect 24276 41020 24286 41076
rect 28130 41020 28140 41076
rect 28196 41020 29260 41076
rect 29316 41020 29326 41076
rect 30314 41020 30324 41076
rect 30380 41020 31052 41076
rect 31108 41020 31118 41076
rect 44370 41020 44380 41076
rect 44436 41020 45948 41076
rect 46004 41020 46620 41076
rect 46676 41020 48860 41076
rect 48916 41020 48926 41076
rect 18106 40908 18116 40964
rect 18172 40908 20356 40964
rect 20412 40908 21532 40964
rect 21588 40908 21598 40964
rect 22642 40908 22652 40964
rect 22708 40908 24108 40964
rect 24164 40908 24174 40964
rect 25890 40908 25900 40964
rect 25956 40908 26460 40964
rect 26516 40908 26526 40964
rect 39890 40908 39900 40964
rect 39956 40908 40572 40964
rect 40628 40908 41076 40964
rect 41132 40908 41692 40964
rect 41748 40908 41758 40964
rect 42252 40908 42364 40964
rect 42420 40908 42430 40964
rect 43866 40908 43876 40964
rect 43932 40908 47068 40964
rect 47124 40908 47134 40964
rect 16146 40796 16156 40852
rect 16212 40796 17276 40852
rect 17332 40796 19068 40852
rect 19124 40796 19134 40852
rect 27626 40796 27636 40852
rect 27748 40796 29932 40852
rect 29988 40796 29998 40852
rect 30818 40796 30828 40852
rect 30884 40796 32060 40852
rect 32116 40796 32126 40852
rect 37426 40796 37436 40852
rect 37492 40796 40236 40852
rect 40292 40796 40302 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 42252 40740 42308 40908
rect 10210 40684 10220 40740
rect 10276 40684 11116 40740
rect 11172 40684 11182 40740
rect 12786 40684 12796 40740
rect 12852 40684 13244 40740
rect 13300 40684 14812 40740
rect 14868 40684 14878 40740
rect 21970 40684 21980 40740
rect 22036 40684 22316 40740
rect 22372 40684 22382 40740
rect 24546 40684 24556 40740
rect 24612 40684 28476 40740
rect 28532 40684 28542 40740
rect 28690 40684 28700 40740
rect 28756 40684 29260 40740
rect 29316 40684 29326 40740
rect 35186 40684 35196 40740
rect 35252 40684 40124 40740
rect 40180 40684 40190 40740
rect 41514 40684 41524 40740
rect 41580 40684 42308 40740
rect 48066 40684 48076 40740
rect 48132 40684 48412 40740
rect 48468 40684 48478 40740
rect 6738 40572 6748 40628
rect 6804 40572 7644 40628
rect 7700 40572 7710 40628
rect 8866 40572 8876 40628
rect 8932 40572 9660 40628
rect 9716 40572 9884 40628
rect 9940 40572 9950 40628
rect 10322 40572 10332 40628
rect 10388 40572 11452 40628
rect 11508 40572 11518 40628
rect 12562 40572 12572 40628
rect 12628 40572 16044 40628
rect 16100 40572 16110 40628
rect 20748 40572 22428 40628
rect 22484 40572 23884 40628
rect 23940 40572 23950 40628
rect 25554 40572 25564 40628
rect 25620 40572 26124 40628
rect 26180 40572 28028 40628
rect 28084 40572 28094 40628
rect 28242 40572 28252 40628
rect 28308 40572 28980 40628
rect 29036 40572 29820 40628
rect 29876 40572 29886 40628
rect 30258 40572 30268 40628
rect 30324 40572 30940 40628
rect 30996 40572 31006 40628
rect 33058 40572 33068 40628
rect 33124 40572 34468 40628
rect 34580 40572 34972 40628
rect 35028 40572 35038 40628
rect 36418 40572 36428 40628
rect 36484 40572 37156 40628
rect 37212 40572 37222 40628
rect 37874 40572 37884 40628
rect 37940 40572 38780 40628
rect 38836 40572 38846 40628
rect 39330 40572 39340 40628
rect 39396 40572 43708 40628
rect 49074 40572 49084 40628
rect 49140 40572 49150 40628
rect 20748 40516 20804 40572
rect 5394 40460 5404 40516
rect 5460 40460 5964 40516
rect 6020 40460 6188 40516
rect 6244 40460 8316 40516
rect 8372 40460 10220 40516
rect 10276 40460 10286 40516
rect 20738 40460 20748 40516
rect 20804 40460 20814 40516
rect 24322 40460 24332 40516
rect 24388 40460 24668 40516
rect 24724 40460 25732 40516
rect 28130 40460 28140 40516
rect 28196 40460 30044 40516
rect 30100 40460 30110 40516
rect 37258 40460 37268 40516
rect 37324 40460 39676 40516
rect 39732 40460 39742 40516
rect 40450 40460 40460 40516
rect 40516 40460 41804 40516
rect 41860 40460 42924 40516
rect 42980 40460 42990 40516
rect 25676 40404 25732 40460
rect 43652 40404 43708 40572
rect 49084 40516 49140 40572
rect 44202 40460 44212 40516
rect 44268 40460 45052 40516
rect 45108 40460 45118 40516
rect 46946 40460 46956 40516
rect 47012 40460 48412 40516
rect 48468 40460 49140 40516
rect 50200 40404 51000 40432
rect 6626 40348 6636 40404
rect 6692 40348 8204 40404
rect 8260 40348 8270 40404
rect 9762 40348 9772 40404
rect 9828 40348 10668 40404
rect 10724 40348 10734 40404
rect 12898 40348 12908 40404
rect 12964 40348 14476 40404
rect 14532 40348 14542 40404
rect 15362 40348 15372 40404
rect 15428 40348 17724 40404
rect 17780 40348 19964 40404
rect 20020 40348 20030 40404
rect 23426 40348 23436 40404
rect 23492 40348 24444 40404
rect 24500 40348 24510 40404
rect 24938 40348 24948 40404
rect 25004 40348 25452 40404
rect 25508 40348 25518 40404
rect 25676 40348 26628 40404
rect 26684 40348 27692 40404
rect 27748 40348 27758 40404
rect 29362 40348 29372 40404
rect 29428 40348 29708 40404
rect 29764 40348 29774 40404
rect 34850 40348 34860 40404
rect 34916 40348 36764 40404
rect 36820 40348 36830 40404
rect 36978 40348 36988 40404
rect 37044 40348 40796 40404
rect 40852 40348 41356 40404
rect 41412 40348 41422 40404
rect 42578 40348 42588 40404
rect 42644 40348 43372 40404
rect 43428 40348 43438 40404
rect 43652 40348 44492 40404
rect 44548 40348 45276 40404
rect 45332 40348 46284 40404
rect 46340 40348 46350 40404
rect 47058 40348 47068 40404
rect 47124 40348 51000 40404
rect 36764 40292 36820 40348
rect 50200 40320 51000 40348
rect 5842 40236 5852 40292
rect 5908 40236 6524 40292
rect 6580 40236 6590 40292
rect 10098 40236 10108 40292
rect 10164 40236 10780 40292
rect 10836 40236 10846 40292
rect 11442 40236 11452 40292
rect 11508 40236 14252 40292
rect 14308 40236 14318 40292
rect 33058 40236 33068 40292
rect 33124 40236 33292 40292
rect 33348 40236 33358 40292
rect 35298 40236 35308 40292
rect 35364 40236 35980 40292
rect 36036 40236 36046 40292
rect 36764 40236 37324 40292
rect 37380 40236 37390 40292
rect 49074 40236 49084 40292
rect 49140 40236 49420 40292
rect 49476 40236 49486 40292
rect 30482 40124 30492 40180
rect 30548 40124 31612 40180
rect 31668 40124 31678 40180
rect 36530 40124 36540 40180
rect 36596 40124 36764 40180
rect 36820 40124 36830 40180
rect 13010 40012 13020 40068
rect 13076 40012 15148 40068
rect 21942 40012 21980 40068
rect 22036 40012 22046 40068
rect 26786 40012 26796 40068
rect 26852 40012 34076 40068
rect 34132 40012 34142 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 15092 39956 15148 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 10882 39900 10892 39956
rect 10948 39900 13076 39956
rect 15092 39900 16492 39956
rect 16548 39900 16558 39956
rect 27654 39900 27692 39956
rect 27748 39900 27758 39956
rect 13020 39844 13076 39900
rect 7298 39788 7308 39844
rect 7364 39788 11676 39844
rect 11732 39788 11742 39844
rect 13020 39788 19292 39844
rect 19348 39788 19358 39844
rect 27570 39788 27580 39844
rect 27636 39788 28476 39844
rect 28532 39788 28542 39844
rect 35410 39788 35420 39844
rect 35476 39788 38668 39844
rect 38724 39788 38734 39844
rect 43474 39788 43484 39844
rect 43540 39788 45612 39844
rect 45668 39788 45678 39844
rect 45994 39788 46004 39844
rect 46060 39788 46956 39844
rect 47012 39788 47022 39844
rect 6402 39676 6412 39732
rect 6468 39676 6860 39732
rect 6916 39676 7756 39732
rect 7812 39676 7822 39732
rect 8810 39676 8820 39732
rect 8876 39676 9212 39732
rect 9268 39676 9278 39732
rect 11442 39676 11452 39732
rect 11508 39676 12012 39732
rect 12068 39676 12078 39732
rect 15026 39676 15036 39732
rect 15092 39676 16716 39732
rect 16772 39676 16782 39732
rect 37538 39676 37548 39732
rect 37604 39676 38108 39732
rect 38164 39676 38174 39732
rect 42522 39676 42532 39732
rect 42588 39676 44492 39732
rect 44548 39676 44558 39732
rect 46386 39676 46396 39732
rect 46452 39676 47068 39732
rect 47124 39676 47134 39732
rect 37772 39620 37828 39676
rect 5954 39564 5964 39620
rect 6020 39564 11228 39620
rect 11284 39564 11294 39620
rect 14802 39564 14812 39620
rect 14868 39564 15762 39620
rect 15818 39564 15828 39620
rect 19394 39564 19404 39620
rect 19460 39564 20300 39620
rect 20356 39564 20366 39620
rect 28410 39564 28420 39620
rect 28476 39564 29876 39620
rect 29932 39564 29942 39620
rect 30034 39564 30044 39620
rect 30100 39564 30604 39620
rect 30660 39564 30670 39620
rect 33730 39564 33740 39620
rect 33796 39564 34972 39620
rect 35028 39564 35420 39620
rect 35476 39564 35486 39620
rect 36530 39564 36540 39620
rect 36596 39564 36988 39620
rect 37044 39564 37054 39620
rect 37762 39564 37772 39620
rect 37828 39564 37838 39620
rect 45490 39564 45500 39620
rect 45556 39564 45948 39620
rect 46004 39564 46014 39620
rect 6290 39452 6300 39508
rect 6356 39452 8316 39508
rect 8372 39452 8382 39508
rect 14914 39452 14924 39508
rect 14980 39452 15484 39508
rect 15540 39452 15550 39508
rect 19058 39452 19068 39508
rect 19124 39452 20188 39508
rect 20244 39452 20254 39508
rect 20514 39452 20524 39508
rect 20580 39452 21084 39508
rect 21140 39452 23436 39508
rect 23492 39452 23502 39508
rect 11778 39340 11788 39396
rect 11844 39340 15708 39396
rect 15764 39340 15774 39396
rect 18498 39340 18508 39396
rect 18564 39340 20412 39396
rect 20468 39340 20860 39396
rect 20916 39340 20926 39396
rect 40674 39340 40684 39396
rect 40740 39340 41244 39396
rect 41300 39340 42532 39396
rect 42588 39340 42598 39396
rect 44594 39340 44604 39396
rect 44660 39340 48300 39396
rect 48356 39340 48366 39396
rect 9202 39228 9212 39284
rect 9268 39228 9548 39284
rect 9604 39228 10444 39284
rect 10500 39228 10510 39284
rect 20962 39228 20972 39284
rect 21028 39228 21308 39284
rect 21364 39228 28364 39284
rect 28420 39228 28430 39284
rect 32556 39228 32566 39284
rect 32622 39228 33796 39284
rect 33852 39228 41636 39284
rect 41692 39228 47234 39284
rect 47290 39228 47300 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 11218 39116 11228 39172
rect 11284 39116 11788 39172
rect 11844 39116 11854 39172
rect 25106 39116 25116 39172
rect 25172 39116 31612 39172
rect 31668 39116 33348 39172
rect 33404 39116 36876 39172
rect 36932 39116 38444 39172
rect 38500 39116 38510 39172
rect 43250 39116 43260 39172
rect 43316 39116 44156 39172
rect 44212 39116 44884 39172
rect 44940 39116 44950 39172
rect 10434 39004 10444 39060
rect 10500 39004 12124 39060
rect 12180 39004 12190 39060
rect 18162 39004 18172 39060
rect 18228 39004 20188 39060
rect 20244 39004 20972 39060
rect 21028 39004 21038 39060
rect 23090 39004 23100 39060
rect 23156 39004 26124 39060
rect 26180 39004 26190 39060
rect 28802 39004 28812 39060
rect 28868 39004 29932 39060
rect 29988 39004 31724 39060
rect 31780 39004 33180 39060
rect 33236 39004 33246 39060
rect 36754 39004 36764 39060
rect 36820 39004 36830 39060
rect 37090 39004 37100 39060
rect 37156 39004 37324 39060
rect 37380 39004 37390 39060
rect 42074 39004 42084 39060
rect 42140 39004 47180 39060
rect 47236 39004 47246 39060
rect 36764 38948 36820 39004
rect 5730 38892 5740 38948
rect 5796 38892 6524 38948
rect 6580 38892 6590 38948
rect 8978 38892 8988 38948
rect 9044 38892 9660 38948
rect 9716 38892 9726 38948
rect 10042 38892 10052 38948
rect 10108 38892 12460 38948
rect 12516 38892 12526 38948
rect 15362 38892 15372 38948
rect 15428 38892 15876 38948
rect 15932 38892 16828 38948
rect 16884 38892 16894 38948
rect 29250 38892 29260 38948
rect 29316 38892 31948 38948
rect 32004 38892 33516 38948
rect 33572 38892 33582 38948
rect 35634 38892 35644 38948
rect 35700 38892 36876 38948
rect 36932 38892 36942 38948
rect 44828 38892 45836 38948
rect 45892 38892 45902 38948
rect 44828 38836 44884 38892
rect 5506 38780 5516 38836
rect 5572 38780 6188 38836
rect 6244 38780 6254 38836
rect 7634 38780 7644 38836
rect 7700 38780 7710 38836
rect 8586 38780 8596 38836
rect 8652 38780 11004 38836
rect 11060 38780 13580 38836
rect 13636 38780 13646 38836
rect 14634 38780 14644 38836
rect 14700 38780 15484 38836
rect 15540 38780 15550 38836
rect 23314 38780 23324 38836
rect 23380 38780 25116 38836
rect 25172 38780 25788 38836
rect 25844 38780 25854 38836
rect 32162 38780 32172 38836
rect 32228 38780 33180 38836
rect 33236 38780 33246 38836
rect 34850 38780 34860 38836
rect 34916 38780 35980 38836
rect 36036 38780 36046 38836
rect 36204 38780 37100 38836
rect 37156 38780 37166 38836
rect 37594 38780 37604 38836
rect 37660 38780 37996 38836
rect 38052 38780 38062 38836
rect 44482 38780 44492 38836
rect 44548 38780 44828 38836
rect 44884 38780 44894 38836
rect 45266 38780 45276 38836
rect 45332 38780 45342 38836
rect 46834 38780 46844 38836
rect 46900 38780 47404 38836
rect 47460 38780 48860 38836
rect 48916 38780 48926 38836
rect 7644 38724 7700 38780
rect 36204 38724 36260 38780
rect 3490 38668 3500 38724
rect 3556 38668 9772 38724
rect 9828 38668 9838 38724
rect 15586 38668 15596 38724
rect 15652 38668 16548 38724
rect 16604 38668 16614 38724
rect 19954 38668 19964 38724
rect 20020 38668 20300 38724
rect 20356 38668 20860 38724
rect 20916 38668 20926 38724
rect 22306 38668 22316 38724
rect 22372 38668 23772 38724
rect 23828 38668 25676 38724
rect 25732 38668 25742 38724
rect 26562 38668 26572 38724
rect 26628 38668 27580 38724
rect 27636 38668 27646 38724
rect 33282 38668 33292 38724
rect 33348 38668 35084 38724
rect 35140 38668 35150 38724
rect 36082 38668 36092 38724
rect 36148 38668 36260 38724
rect 36754 38668 36764 38724
rect 36820 38668 38948 38724
rect 39004 38668 39014 38724
rect 45276 38612 45332 38780
rect 8418 38556 8428 38612
rect 8484 38556 9492 38612
rect 9548 38556 9558 38612
rect 16930 38556 16940 38612
rect 16996 38556 17948 38612
rect 18004 38556 18014 38612
rect 28354 38556 28364 38612
rect 28420 38556 32004 38612
rect 33702 38556 33740 38612
rect 33796 38556 33806 38612
rect 35746 38556 35756 38612
rect 35812 38556 36316 38612
rect 36372 38556 36382 38612
rect 37426 38556 37436 38612
rect 37492 38556 40460 38612
rect 40516 38556 40526 38612
rect 45276 38556 46620 38612
rect 46676 38556 46686 38612
rect 30268 38500 30324 38556
rect 31948 38500 32004 38556
rect 9314 38444 9324 38500
rect 9380 38444 9996 38500
rect 10052 38444 10062 38500
rect 22306 38444 22316 38500
rect 22372 38444 23996 38500
rect 24052 38444 25004 38500
rect 25060 38444 25070 38500
rect 30258 38444 30268 38500
rect 30324 38444 30334 38500
rect 30818 38444 30828 38500
rect 30884 38444 31780 38500
rect 31836 38444 31846 38500
rect 31948 38444 33964 38500
rect 34020 38444 34030 38500
rect 44594 38444 44604 38500
rect 44660 38444 45276 38500
rect 45332 38444 45342 38500
rect 47898 38444 47908 38500
rect 47964 38444 48636 38500
rect 48692 38444 48702 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 14802 38332 14812 38388
rect 14868 38332 15820 38388
rect 15876 38332 15886 38388
rect 24434 38332 24444 38388
rect 24500 38332 26012 38388
rect 26068 38332 28476 38388
rect 28532 38332 31612 38388
rect 31668 38332 31678 38388
rect 44706 38332 44716 38388
rect 44772 38332 44940 38388
rect 44996 38332 45006 38388
rect 8866 38220 8876 38276
rect 8932 38220 9884 38276
rect 9940 38220 10612 38276
rect 10668 38220 10678 38276
rect 17938 38220 17948 38276
rect 18004 38220 20804 38276
rect 22194 38220 22204 38276
rect 22260 38220 23324 38276
rect 23380 38220 23390 38276
rect 28914 38220 28924 38276
rect 28980 38220 29596 38276
rect 29652 38220 29662 38276
rect 32162 38220 32172 38276
rect 32228 38220 32956 38276
rect 33012 38220 33022 38276
rect 44034 38220 44044 38276
rect 44100 38220 46508 38276
rect 46564 38220 46574 38276
rect 8194 38108 8204 38164
rect 8260 38108 8428 38164
rect 8484 38108 8494 38164
rect 9762 38108 9772 38164
rect 9828 38108 10108 38164
rect 10164 38108 10174 38164
rect 15250 38108 15260 38164
rect 15316 38108 15932 38164
rect 15988 38108 17500 38164
rect 17556 38108 17566 38164
rect 18610 38108 18620 38164
rect 18676 38108 18844 38164
rect 18900 38108 18910 38164
rect 20748 38052 20804 38220
rect 28578 38108 28588 38164
rect 28644 38108 29260 38164
rect 29316 38108 29326 38164
rect 42485 38108 42495 38164
rect 42551 38108 43708 38164
rect 43764 38108 44268 38164
rect 44324 38108 44334 38164
rect 46050 38108 46060 38164
rect 46116 38108 46732 38164
rect 46788 38108 46798 38164
rect 48514 38108 48524 38164
rect 48580 38108 49196 38164
rect 49252 38108 49262 38164
rect 9538 37996 9548 38052
rect 9604 37996 10332 38052
rect 10388 37996 10398 38052
rect 11666 37996 11676 38052
rect 11732 37996 12348 38052
rect 12404 37996 12414 38052
rect 16034 37996 16044 38052
rect 16100 37996 17388 38052
rect 17444 37996 17454 38052
rect 18386 37996 18396 38052
rect 18452 37996 19292 38052
rect 19348 37996 19358 38052
rect 20738 37996 20748 38052
rect 20804 37996 21308 38052
rect 21364 37996 21374 38052
rect 22082 37996 22092 38052
rect 22148 37996 22316 38052
rect 22372 37996 22382 38052
rect 29586 37996 29596 38052
rect 29652 37996 30604 38052
rect 30660 37996 30670 38052
rect 32498 37996 32508 38052
rect 32564 37996 32956 38052
rect 33012 37996 33022 38052
rect 36362 37996 36372 38052
rect 36428 37996 36876 38052
rect 36932 37996 36942 38052
rect 40562 37996 40572 38052
rect 40628 37996 41244 38052
rect 41300 37996 41310 38052
rect 41570 37996 41580 38052
rect 41636 37996 42252 38052
rect 42308 37996 42318 38052
rect 44146 37996 44156 38052
rect 44212 37996 44492 38052
rect 44548 37996 44558 38052
rect 44930 37996 44940 38052
rect 44996 37996 45164 38052
rect 45220 37996 45230 38052
rect 41244 37940 41300 37996
rect 19114 37884 19124 37940
rect 19180 37884 20300 37940
rect 20356 37884 20972 37940
rect 21028 37884 21038 37940
rect 21970 37884 21980 37940
rect 22036 37884 24668 37940
rect 24724 37884 24734 37940
rect 29362 37884 29372 37940
rect 29428 37884 31332 37940
rect 31388 37884 31398 37940
rect 41244 37884 44044 37940
rect 44100 37884 44110 37940
rect 12226 37772 12236 37828
rect 12292 37772 20580 37828
rect 23986 37772 23996 37828
rect 24052 37772 24220 37828
rect 24276 37772 29820 37828
rect 29876 37772 30380 37828
rect 30436 37772 30446 37828
rect 31948 37772 33908 37828
rect 34020 37772 34030 37828
rect 39106 37772 39116 37828
rect 39172 37772 40348 37828
rect 40404 37772 40414 37828
rect 43810 37772 43820 37828
rect 43876 37772 45164 37828
rect 45220 37772 45230 37828
rect 46274 37772 46284 37828
rect 46340 37772 48188 37828
rect 48244 37772 48748 37828
rect 48804 37772 48814 37828
rect 20524 37716 20580 37772
rect 31948 37716 32004 37772
rect 9174 37660 9212 37716
rect 9268 37660 9278 37716
rect 20514 37660 20524 37716
rect 20580 37660 21420 37716
rect 21476 37660 21486 37716
rect 25722 37660 25732 37716
rect 25788 37660 32004 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 11890 37548 11900 37604
rect 11956 37548 12460 37604
rect 12516 37548 12526 37604
rect 26674 37548 26684 37604
rect 26740 37548 27132 37604
rect 27188 37548 27198 37604
rect 34458 37548 34468 37604
rect 34524 37548 34860 37604
rect 34916 37548 35532 37604
rect 35588 37548 35598 37604
rect 47170 37548 47180 37604
rect 47236 37548 47740 37604
rect 47796 37548 47806 37604
rect 12226 37436 12236 37492
rect 12292 37436 12908 37492
rect 12964 37436 12974 37492
rect 18610 37436 18620 37492
rect 18676 37436 20076 37492
rect 20132 37436 20142 37492
rect 20300 37436 21924 37492
rect 24994 37436 25004 37492
rect 25060 37436 25732 37492
rect 25788 37436 25798 37492
rect 41010 37436 41020 37492
rect 41076 37436 41356 37492
rect 41412 37436 46620 37492
rect 46676 37436 49084 37492
rect 49140 37436 49150 37492
rect 20300 37380 20356 37436
rect 21868 37380 21924 37436
rect 12562 37324 12572 37380
rect 12628 37324 17500 37380
rect 17556 37324 17566 37380
rect 17733 37324 17743 37380
rect 17799 37324 17948 37380
rect 18004 37324 20356 37380
rect 21196 37324 21644 37380
rect 21700 37324 21710 37380
rect 21868 37324 31892 37380
rect 31948 37324 32396 37380
rect 32452 37324 34168 37380
rect 34224 37324 34234 37380
rect 36082 37324 36092 37380
rect 36148 37324 39116 37380
rect 39172 37324 39182 37380
rect 40394 37324 40404 37380
rect 40460 37324 41804 37380
rect 41860 37324 44268 37380
rect 44324 37324 44334 37380
rect 21196 37268 21252 37324
rect 15810 37212 15820 37268
rect 15876 37212 18620 37268
rect 18676 37212 20636 37268
rect 20692 37212 21252 37268
rect 21410 37212 21420 37268
rect 21476 37212 22204 37268
rect 22260 37212 22270 37268
rect 29026 37212 29036 37268
rect 29092 37212 29260 37268
rect 29316 37212 29326 37268
rect 29810 37212 29820 37268
rect 29876 37212 30828 37268
rect 30884 37212 30894 37268
rect 33282 37212 33292 37268
rect 33348 37212 33358 37268
rect 40786 37212 40796 37268
rect 40852 37212 42364 37268
rect 42420 37212 42430 37268
rect 44902 37212 44940 37268
rect 44996 37212 45006 37268
rect 33292 37156 33348 37212
rect 33292 37100 33908 37156
rect 35298 37100 35308 37156
rect 35364 37100 36148 37156
rect 36204 37100 40684 37156
rect 40740 37100 40750 37156
rect 12114 36988 12124 37044
rect 12180 36988 17836 37044
rect 17892 36988 18956 37044
rect 19012 36988 19022 37044
rect 23930 36988 23940 37044
rect 23996 36988 24444 37044
rect 24500 36988 24510 37044
rect 26878 36988 26888 37044
rect 26944 36988 27748 37044
rect 27804 36988 32060 37044
rect 32116 36988 32620 37044
rect 32676 36988 33348 37044
rect 33292 36932 33348 36988
rect 7858 36876 7868 36932
rect 7924 36876 8428 36932
rect 8484 36876 8494 36932
rect 24658 36876 24668 36932
rect 24724 36876 30380 36932
rect 30436 36876 30446 36932
rect 33282 36876 33292 36932
rect 33348 36876 33358 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 33852 36820 33908 37100
rect 35186 36988 35196 37044
rect 35252 36988 35644 37044
rect 35700 36988 35710 37044
rect 40226 36988 40236 37044
rect 40292 36988 41244 37044
rect 41300 36988 41310 37044
rect 38546 36876 38556 36932
rect 38612 36876 39732 36932
rect 39788 36876 39798 36932
rect 44370 36876 44380 36932
rect 44436 36876 48860 36932
rect 48916 36876 48926 36932
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 33842 36764 33852 36820
rect 33908 36764 33918 36820
rect 20794 36652 20804 36708
rect 20860 36652 22652 36708
rect 22708 36652 32284 36708
rect 32340 36652 32350 36708
rect 30482 36540 30492 36596
rect 30548 36540 31724 36596
rect 31780 36540 31790 36596
rect 6626 36428 6636 36484
rect 6692 36428 10780 36484
rect 10836 36428 10846 36484
rect 12562 36428 12572 36484
rect 12628 36428 15372 36484
rect 15428 36428 16716 36484
rect 16772 36428 19516 36484
rect 19572 36428 19582 36484
rect 20962 36428 20972 36484
rect 21028 36428 23660 36484
rect 23716 36428 23726 36484
rect 27356 36428 28028 36484
rect 28084 36428 29596 36484
rect 29652 36428 29662 36484
rect 33170 36428 33180 36484
rect 33236 36428 33964 36484
rect 34020 36428 34030 36484
rect 35634 36428 35644 36484
rect 35700 36428 36540 36484
rect 36596 36428 36606 36484
rect 43810 36428 43820 36484
rect 43876 36428 44940 36484
rect 44996 36428 45006 36484
rect 45126 36428 45164 36484
rect 45220 36428 45948 36484
rect 46004 36428 46014 36484
rect 27356 36372 27412 36428
rect 27346 36316 27356 36372
rect 27412 36316 27422 36372
rect 28028 36316 28364 36372
rect 28420 36316 29316 36372
rect 29372 36316 29382 36372
rect 46106 36316 46116 36372
rect 46172 36316 46732 36372
rect 46788 36316 46798 36372
rect 28028 36260 28084 36316
rect 28018 36204 28028 36260
rect 28084 36204 28094 36260
rect 39330 36204 39340 36260
rect 39396 36204 41020 36260
rect 41076 36204 41086 36260
rect 44034 36204 44044 36260
rect 44100 36204 47740 36260
rect 47796 36204 47806 36260
rect 50200 36148 51000 36176
rect 20514 36092 20524 36148
rect 20580 36092 21196 36148
rect 21252 36092 23772 36148
rect 23828 36092 31612 36148
rect 31668 36092 33628 36148
rect 33684 36092 33694 36148
rect 35522 36092 35532 36148
rect 35588 36092 36204 36148
rect 36260 36092 36270 36148
rect 36428 36092 38668 36148
rect 48850 36092 48860 36148
rect 48916 36092 51000 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 36428 36036 36484 36092
rect 38612 36036 38668 36092
rect 50200 36064 51000 36092
rect 26114 35980 26124 36036
rect 26180 35980 27524 36036
rect 27580 35980 27590 36036
rect 30370 35980 30380 36036
rect 30436 35980 31220 36036
rect 31276 35980 32060 36036
rect 32116 35980 36484 36036
rect 37090 35980 37100 36036
rect 37156 35980 37828 36036
rect 37884 35924 37940 36036
rect 38612 35980 40572 36036
rect 40628 35980 40638 36036
rect 45836 35980 48972 36036
rect 49028 35980 49038 36036
rect 45836 35924 45892 35980
rect 8082 35868 8092 35924
rect 8148 35868 8764 35924
rect 8820 35868 8830 35924
rect 16482 35868 16492 35924
rect 16548 35868 18396 35924
rect 18452 35868 18462 35924
rect 25106 35868 25116 35924
rect 25172 35868 25788 35924
rect 25844 35868 25854 35924
rect 32498 35868 32508 35924
rect 32564 35868 35420 35924
rect 35476 35868 35486 35924
rect 37884 35868 39620 35924
rect 39676 35868 40348 35924
rect 40404 35868 40414 35924
rect 41570 35868 41580 35924
rect 41636 35868 42364 35924
rect 42420 35868 42430 35924
rect 45154 35868 45164 35924
rect 45220 35868 45836 35924
rect 45892 35868 45902 35924
rect 47170 35868 47180 35924
rect 47236 35868 48748 35924
rect 48804 35868 48814 35924
rect 7858 35756 7868 35812
rect 7924 35756 11116 35812
rect 11172 35756 11182 35812
rect 17210 35756 17220 35812
rect 17276 35756 18844 35812
rect 18900 35756 18910 35812
rect 27682 35756 27692 35812
rect 27748 35756 28140 35812
rect 28196 35756 34860 35812
rect 34916 35756 34926 35812
rect 41430 35756 41468 35812
rect 41524 35756 41534 35812
rect 47254 35756 47292 35812
rect 47348 35756 47358 35812
rect 20290 35644 20300 35700
rect 20356 35644 20804 35700
rect 20860 35644 20870 35700
rect 22866 35644 22876 35700
rect 22932 35644 25396 35700
rect 25452 35644 25462 35700
rect 27122 35644 27132 35700
rect 27188 35644 28476 35700
rect 28532 35644 28542 35700
rect 32722 35644 32732 35700
rect 32788 35644 33180 35700
rect 33236 35644 33404 35700
rect 33460 35644 37324 35700
rect 37380 35644 37390 35700
rect 45266 35644 45276 35700
rect 45332 35644 45612 35700
rect 45668 35644 46508 35700
rect 46564 35644 49084 35700
rect 49140 35644 49150 35700
rect 10546 35532 10556 35588
rect 10612 35532 10948 35588
rect 11004 35532 16380 35588
rect 16436 35532 16446 35588
rect 18722 35532 18732 35588
rect 18788 35532 20188 35588
rect 20244 35532 25564 35588
rect 25620 35532 25630 35588
rect 29250 35532 29260 35588
rect 29316 35532 30660 35588
rect 30716 35532 30726 35588
rect 34972 35532 37660 35588
rect 37716 35532 37726 35588
rect 14242 35420 14252 35476
rect 14308 35420 15932 35476
rect 15988 35420 15998 35476
rect 23650 35420 23660 35476
rect 23716 35420 24612 35476
rect 24668 35420 26516 35476
rect 26572 35420 26908 35476
rect 27570 35420 27580 35476
rect 27636 35420 28364 35476
rect 28420 35420 28924 35476
rect 28980 35420 29372 35476
rect 29428 35420 29438 35476
rect 26852 35364 26908 35420
rect 12674 35308 12684 35364
rect 12740 35308 12908 35364
rect 12964 35308 15148 35364
rect 15204 35308 16492 35364
rect 16548 35308 16558 35364
rect 16874 35308 16884 35364
rect 16940 35308 17500 35364
rect 17556 35308 22876 35364
rect 22932 35308 22942 35364
rect 23202 35308 23212 35364
rect 23268 35308 23436 35364
rect 23492 35308 24220 35364
rect 24276 35308 24286 35364
rect 26852 35308 34412 35364
rect 34468 35308 34916 35364
rect 34972 35308 35028 35532
rect 37314 35420 37324 35476
rect 37380 35420 38892 35476
rect 38948 35420 38958 35476
rect 40226 35420 40236 35476
rect 40292 35420 41244 35476
rect 41300 35420 41804 35476
rect 41860 35420 41870 35476
rect 37874 35308 37884 35364
rect 37940 35308 38220 35364
rect 38276 35308 38286 35364
rect 40562 35308 40572 35364
rect 40628 35308 41580 35364
rect 41636 35308 41646 35364
rect 44146 35308 44156 35364
rect 44212 35308 45276 35364
rect 45332 35308 45342 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 14914 35196 14924 35252
rect 14980 35196 15372 35252
rect 15428 35196 15438 35252
rect 21634 35196 21644 35252
rect 21700 35196 22204 35252
rect 22260 35196 22270 35252
rect 36418 35196 36428 35252
rect 36484 35196 40460 35252
rect 40516 35196 40526 35252
rect 41458 35196 41468 35252
rect 41524 35196 43596 35252
rect 43652 35196 45164 35252
rect 45220 35196 45230 35252
rect 45602 35196 45612 35252
rect 45668 35196 45836 35252
rect 45892 35196 45902 35252
rect 20066 35084 20076 35140
rect 20132 35084 20972 35140
rect 21028 35084 21038 35140
rect 21298 35084 21308 35140
rect 21364 35084 21980 35140
rect 22036 35084 22046 35140
rect 31938 34972 31948 35028
rect 32004 34972 32396 35028
rect 32452 34972 32956 35028
rect 33012 34972 33516 35028
rect 33572 34972 33740 35028
rect 33796 34972 33806 35028
rect 34066 34972 34076 35028
rect 34132 34972 35532 35028
rect 35588 34972 41468 35028
rect 41524 34972 41692 35028
rect 41748 34972 41758 35028
rect 42130 34972 42140 35028
rect 42196 34972 43260 35028
rect 43316 34972 46956 35028
rect 47012 34972 47022 35028
rect 4834 34860 4844 34916
rect 4900 34860 5180 34916
rect 5236 34860 5516 34916
rect 5572 34860 5582 34916
rect 7410 34860 7420 34916
rect 7476 34860 10108 34916
rect 10164 34860 10174 34916
rect 17686 34860 17724 34916
rect 17780 34860 17790 34916
rect 37650 34860 37660 34916
rect 37716 34860 38444 34916
rect 38500 34860 38510 34916
rect 40674 34860 40684 34916
rect 40740 34860 42588 34916
rect 42644 34860 42654 34916
rect 46060 34860 46172 34916
rect 46228 34860 46238 34916
rect 46386 34860 46396 34916
rect 46452 34860 49420 34916
rect 49476 34860 49486 34916
rect 46060 34804 46116 34860
rect 12226 34748 12236 34804
rect 12292 34748 12796 34804
rect 12852 34748 12862 34804
rect 18162 34748 18172 34804
rect 18228 34748 21420 34804
rect 21476 34748 21486 34804
rect 29362 34748 29372 34804
rect 29428 34748 31500 34804
rect 31556 34748 31724 34804
rect 31780 34748 31790 34804
rect 33506 34748 33516 34804
rect 33572 34748 33852 34804
rect 33908 34748 34076 34804
rect 34132 34748 36932 34804
rect 36988 34748 36998 34804
rect 37762 34748 37772 34804
rect 37828 34748 38892 34804
rect 38948 34748 38958 34804
rect 42018 34748 42028 34804
rect 42084 34748 42756 34804
rect 42812 34748 42822 34804
rect 45434 34748 45444 34804
rect 45500 34748 46116 34804
rect 46274 34748 46284 34804
rect 46340 34748 49084 34804
rect 49140 34748 49150 34804
rect 6626 34636 6636 34692
rect 6692 34636 8316 34692
rect 8372 34636 9212 34692
rect 9268 34636 9380 34692
rect 9436 34636 9446 34692
rect 11666 34636 11676 34692
rect 11732 34636 12684 34692
rect 12740 34636 12750 34692
rect 12898 34636 12908 34692
rect 12964 34636 15260 34692
rect 15316 34636 16156 34692
rect 16212 34636 16222 34692
rect 16482 34636 16492 34692
rect 16548 34636 16772 34692
rect 16828 34636 21756 34692
rect 21812 34636 21822 34692
rect 25554 34636 25564 34692
rect 25620 34636 27020 34692
rect 27076 34636 27086 34692
rect 33394 34636 33404 34692
rect 33460 34636 34300 34692
rect 34356 34636 37996 34692
rect 38052 34636 38062 34692
rect 18582 34524 18620 34580
rect 18676 34524 18686 34580
rect 26450 34524 26460 34580
rect 26516 34524 37884 34580
rect 37940 34524 37950 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 45948 34468 46004 34748
rect 6178 34412 6188 34468
rect 6244 34412 9604 34468
rect 9660 34412 9670 34468
rect 9986 34412 9996 34468
rect 10052 34412 10444 34468
rect 10500 34412 13356 34468
rect 13412 34412 13422 34468
rect 18022 34412 18060 34468
rect 18116 34412 18126 34468
rect 28802 34412 28812 34468
rect 28868 34412 30044 34468
rect 30100 34412 31668 34468
rect 31724 34412 36764 34468
rect 36820 34412 36830 34468
rect 45938 34412 45948 34468
rect 46004 34412 46014 34468
rect 10882 34300 10892 34356
rect 10948 34300 12236 34356
rect 12292 34300 12302 34356
rect 26562 34300 26572 34356
rect 26628 34300 27244 34356
rect 27300 34300 27310 34356
rect 29138 34300 29148 34356
rect 29204 34300 29596 34356
rect 29652 34300 29662 34356
rect 29810 34300 29820 34356
rect 29876 34300 30268 34356
rect 30324 34300 30334 34356
rect 33842 34300 33852 34356
rect 33908 34300 33918 34356
rect 36642 34300 36652 34356
rect 36708 34300 36718 34356
rect 39890 34300 39900 34356
rect 39956 34300 42868 34356
rect 47954 34300 47964 34356
rect 48020 34300 48524 34356
rect 48580 34300 48590 34356
rect 16706 34188 16716 34244
rect 16772 34188 17500 34244
rect 17556 34188 17566 34244
rect 18470 34188 18508 34244
rect 18564 34188 18574 34244
rect 27682 34188 27692 34244
rect 27748 34188 32452 34244
rect 32508 34188 32518 34244
rect 5842 34076 5852 34132
rect 5908 34076 6300 34132
rect 6356 34076 6366 34132
rect 8194 34076 8204 34132
rect 8260 34076 9884 34132
rect 9940 34076 9950 34132
rect 13010 34076 13020 34132
rect 13076 34076 13468 34132
rect 13524 34076 15820 34132
rect 15876 34076 15886 34132
rect 16930 34076 16940 34132
rect 16996 34076 17743 34132
rect 17799 34076 19012 34132
rect 19068 34076 19078 34132
rect 20626 34076 20636 34132
rect 20692 34076 21420 34132
rect 21476 34076 21486 34132
rect 24434 34076 24444 34132
rect 24500 34076 26516 34132
rect 26572 34076 26582 34132
rect 33852 34020 33908 34300
rect 36652 34020 36708 34300
rect 37986 34188 37996 34244
rect 38052 34188 39060 34244
rect 39116 34188 39126 34244
rect 41458 34188 41468 34244
rect 41524 34188 41916 34244
rect 41972 34188 41982 34244
rect 42812 34132 42868 34300
rect 41570 34076 41580 34132
rect 41636 34076 42028 34132
rect 42084 34076 42094 34132
rect 42812 34076 42924 34132
rect 42980 34076 42990 34132
rect 43642 34076 43652 34132
rect 43708 34076 49308 34132
rect 49364 34076 49644 34132
rect 49700 34076 49710 34132
rect 20514 33964 20524 34020
rect 20580 33964 20972 34020
rect 21028 33964 21038 34020
rect 33730 33964 33740 34020
rect 33796 33964 33908 34020
rect 33964 33964 34412 34020
rect 34468 33964 34478 34020
rect 35634 33964 35644 34020
rect 35700 33964 38668 34020
rect 40226 33964 40236 34020
rect 40292 33964 48972 34020
rect 49028 33964 49038 34020
rect 33964 33908 34020 33964
rect 7746 33852 7756 33908
rect 7812 33852 8764 33908
rect 8820 33852 8830 33908
rect 16370 33852 16380 33908
rect 16436 33852 19740 33908
rect 19796 33852 19806 33908
rect 20850 33852 20860 33908
rect 20916 33852 21644 33908
rect 21700 33852 21710 33908
rect 33842 33852 33852 33908
rect 33908 33852 34020 33908
rect 34122 33852 34132 33908
rect 34188 33852 35196 33908
rect 35252 33852 35262 33908
rect 38612 33796 38668 33964
rect 12898 33740 12908 33796
rect 12964 33740 13804 33796
rect 13860 33740 13870 33796
rect 17378 33740 17388 33796
rect 17444 33740 17836 33796
rect 17892 33740 17902 33796
rect 37090 33740 37100 33796
rect 37156 33740 37324 33796
rect 37380 33740 37390 33796
rect 38612 33740 39900 33796
rect 39956 33740 39966 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 5506 33628 5516 33684
rect 5572 33628 6972 33684
rect 7028 33628 7420 33684
rect 7476 33628 7486 33684
rect 18050 33628 18060 33684
rect 18116 33628 18172 33684
rect 18228 33628 18238 33684
rect 22876 33628 23884 33684
rect 23940 33628 24780 33684
rect 24836 33628 24846 33684
rect 24994 33628 25004 33684
rect 25060 33628 25070 33684
rect 38546 33628 38556 33684
rect 38612 33628 41972 33684
rect 42028 33628 42038 33684
rect 42578 33628 42588 33684
rect 42644 33628 42924 33684
rect 42980 33628 42990 33684
rect 22876 33572 22932 33628
rect 25004 33572 25060 33628
rect 9090 33516 9100 33572
rect 9156 33516 10164 33572
rect 10220 33516 10230 33572
rect 10322 33516 10332 33572
rect 10388 33516 11564 33572
rect 11620 33516 11630 33572
rect 19394 33516 19404 33572
rect 19460 33516 21532 33572
rect 21588 33516 22652 33572
rect 22708 33516 22718 33572
rect 22866 33516 22876 33572
rect 22932 33516 22942 33572
rect 23762 33516 23772 33572
rect 23828 33516 25060 33572
rect 35634 33516 35644 33572
rect 35700 33516 35756 33572
rect 35812 33516 35822 33572
rect 46610 33516 46620 33572
rect 46676 33516 47292 33572
rect 47348 33516 47404 33572
rect 47460 33516 47470 33572
rect 9986 33404 9996 33460
rect 10052 33404 10668 33460
rect 10724 33404 10734 33460
rect 11004 33404 12684 33460
rect 12740 33404 12750 33460
rect 18498 33404 18508 33460
rect 18564 33404 18620 33460
rect 18676 33404 20188 33460
rect 20244 33404 20254 33460
rect 43138 33404 43148 33460
rect 43204 33404 43820 33460
rect 43876 33404 46844 33460
rect 46900 33404 46910 33460
rect 8978 33292 8988 33348
rect 9044 33292 9660 33348
rect 9716 33292 10444 33348
rect 10500 33292 10510 33348
rect 11004 33236 11060 33404
rect 12786 33292 12796 33348
rect 12852 33292 13580 33348
rect 13636 33292 13646 33348
rect 15138 33292 15148 33348
rect 15204 33292 17724 33348
rect 17780 33292 17790 33348
rect 17938 33292 17948 33348
rect 18004 33292 19740 33348
rect 19796 33292 19806 33348
rect 23202 33292 23212 33348
rect 23268 33292 24108 33348
rect 24164 33292 24174 33348
rect 25778 33292 25788 33348
rect 25844 33292 26460 33348
rect 26516 33292 28700 33348
rect 28756 33292 29036 33348
rect 29092 33292 29708 33348
rect 29764 33292 29774 33348
rect 39330 33292 39340 33348
rect 39396 33292 40908 33348
rect 40964 33292 40974 33348
rect 10994 33180 11004 33236
rect 11060 33180 11070 33236
rect 11890 33180 11900 33236
rect 11956 33180 12460 33236
rect 12516 33180 16380 33236
rect 16436 33180 16446 33236
rect 19226 33180 19236 33236
rect 19292 33180 19964 33236
rect 20020 33180 20300 33236
rect 20356 33180 20366 33236
rect 20524 33180 23772 33236
rect 23828 33180 23838 33236
rect 26842 33180 26852 33236
rect 26908 33180 35644 33236
rect 35700 33180 35710 33236
rect 39442 33180 39452 33236
rect 39508 33180 40292 33236
rect 42914 33180 42924 33236
rect 42980 33180 43876 33236
rect 43932 33180 43942 33236
rect 45602 33180 45612 33236
rect 45668 33180 46116 33236
rect 46172 33180 46182 33236
rect 20524 33124 20580 33180
rect 26852 33124 26908 33180
rect 40236 33124 40292 33180
rect 13570 33068 13580 33124
rect 13636 33068 14700 33124
rect 14756 33068 15484 33124
rect 15540 33068 17388 33124
rect 17444 33068 17454 33124
rect 17714 33068 17724 33124
rect 17780 33068 20580 33124
rect 21746 33068 21756 33124
rect 21812 33068 22540 33124
rect 22596 33068 22606 33124
rect 25106 33068 25116 33124
rect 25172 33068 26908 33124
rect 33954 33068 33964 33124
rect 34020 33068 36372 33124
rect 36428 33068 36438 33124
rect 36530 33068 36540 33124
rect 36596 33068 40012 33124
rect 40068 33068 40078 33124
rect 40236 33068 44492 33124
rect 44548 33068 45836 33124
rect 45892 33068 45902 33124
rect 36316 33012 36372 33068
rect 15698 32956 15708 33012
rect 15764 32956 19628 33012
rect 19684 32956 19694 33012
rect 36316 32956 36764 33012
rect 36820 32956 36830 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 34850 32844 34860 32900
rect 34916 32844 35756 32900
rect 35812 32844 35822 32900
rect 38994 32844 39004 32900
rect 39060 32844 41804 32900
rect 41860 32844 41870 32900
rect 8754 32732 8764 32788
rect 8820 32732 10332 32788
rect 10388 32732 10892 32788
rect 10948 32732 10958 32788
rect 11666 32732 11676 32788
rect 11732 32732 11900 32788
rect 11956 32732 11966 32788
rect 23090 32732 23100 32788
rect 23156 32732 23660 32788
rect 23716 32732 24556 32788
rect 24612 32732 25340 32788
rect 25396 32732 25406 32788
rect 31602 32732 31612 32788
rect 31668 32732 33124 32788
rect 33180 32732 33190 32788
rect 33618 32732 33628 32788
rect 33684 32732 33852 32788
rect 33908 32732 34412 32788
rect 34468 32732 34478 32788
rect 35522 32732 35532 32788
rect 35588 32732 36316 32788
rect 36372 32732 38108 32788
rect 38164 32732 38174 32788
rect 38444 32732 39452 32788
rect 39508 32732 39518 32788
rect 40002 32732 40012 32788
rect 40068 32732 42028 32788
rect 42084 32732 42476 32788
rect 42532 32732 42542 32788
rect 48514 32732 48524 32788
rect 48580 32732 48972 32788
rect 49028 32732 49038 32788
rect 38444 32676 38500 32732
rect 14242 32620 14252 32676
rect 14308 32620 15036 32676
rect 15092 32620 15102 32676
rect 29250 32620 29260 32676
rect 29316 32620 31052 32676
rect 31108 32620 32564 32676
rect 32620 32620 37212 32676
rect 37268 32620 38668 32676
rect 38724 32620 38734 32676
rect 9314 32508 9324 32564
rect 9380 32508 9996 32564
rect 10052 32508 13020 32564
rect 13076 32508 13086 32564
rect 14354 32508 14364 32564
rect 14420 32508 15148 32564
rect 15810 32508 15820 32564
rect 15876 32508 16268 32564
rect 16324 32508 17164 32564
rect 17220 32508 17230 32564
rect 18498 32508 18508 32564
rect 18564 32508 19404 32564
rect 19460 32508 19470 32564
rect 33618 32508 33628 32564
rect 33684 32508 34188 32564
rect 34244 32508 34636 32564
rect 34692 32508 34702 32564
rect 40282 32508 40292 32564
rect 40348 32508 40796 32564
rect 40852 32508 40862 32564
rect 41458 32508 41468 32564
rect 41524 32508 42812 32564
rect 42868 32508 42878 32564
rect 45042 32508 45052 32564
rect 45108 32508 45948 32564
rect 46004 32508 46014 32564
rect 47954 32508 47964 32564
rect 48020 32508 48636 32564
rect 48692 32508 49308 32564
rect 49364 32508 49374 32564
rect 15092 32452 15148 32508
rect 15092 32396 16492 32452
rect 16548 32396 16558 32452
rect 26562 32396 26572 32452
rect 26628 32396 27916 32452
rect 27972 32396 27982 32452
rect 38182 32396 38220 32452
rect 38276 32396 38286 32452
rect 43362 32396 43372 32452
rect 43428 32396 45388 32452
rect 45444 32396 45454 32452
rect 13234 32284 13244 32340
rect 13300 32284 13804 32340
rect 13860 32284 19516 32340
rect 19572 32284 19582 32340
rect 29810 32284 29820 32340
rect 29876 32284 31948 32340
rect 32004 32284 32014 32340
rect 32162 32284 32172 32340
rect 32228 32284 32396 32340
rect 32452 32284 32462 32340
rect 34290 32284 34300 32340
rect 34356 32284 35812 32340
rect 46834 32284 46844 32340
rect 46900 32284 48076 32340
rect 48132 32284 48142 32340
rect 9650 32172 9660 32228
rect 9716 32172 10668 32228
rect 10724 32172 10734 32228
rect 10892 32172 27860 32228
rect 27916 32172 27926 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 10892 32116 10948 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 7522 32060 7532 32116
rect 7588 32060 7598 32116
rect 9090 32060 9100 32116
rect 9156 32060 9772 32116
rect 9828 32060 10332 32116
rect 10388 32060 10948 32116
rect 19142 32060 19180 32116
rect 19236 32060 19246 32116
rect 21522 32060 21532 32116
rect 21588 32060 22652 32116
rect 22708 32060 23212 32116
rect 23268 32060 24444 32116
rect 24500 32060 24510 32116
rect 30370 32060 30380 32116
rect 30436 32060 30446 32116
rect 34262 32060 34300 32116
rect 34356 32060 34366 32116
rect 7532 31892 7588 32060
rect 16370 31948 16380 32004
rect 16436 31948 17836 32004
rect 17892 31948 17902 32004
rect 20514 31948 20524 32004
rect 20580 31948 20860 32004
rect 20916 31948 20926 32004
rect 22306 31948 22316 32004
rect 22372 31948 22932 32004
rect 22988 31948 22998 32004
rect 26002 31948 26012 32004
rect 26068 31948 26078 32004
rect 26012 31892 26068 31948
rect 7532 31836 8540 31892
rect 8596 31836 8606 31892
rect 14466 31836 14476 31892
rect 14532 31836 21420 31892
rect 21476 31836 21486 31892
rect 21634 31836 21644 31892
rect 21700 31836 25676 31892
rect 25732 31836 26068 31892
rect 2034 31724 2044 31780
rect 2100 31724 3164 31780
rect 3220 31724 7084 31780
rect 7140 31724 7150 31780
rect 10098 31724 10108 31780
rect 10164 31724 10612 31780
rect 10668 31724 10678 31780
rect 11237 31724 11247 31780
rect 11303 31724 12796 31780
rect 12852 31724 13132 31780
rect 13188 31724 13198 31780
rect 18274 31724 18284 31780
rect 18340 31724 21308 31780
rect 21364 31724 22484 31780
rect 22540 31724 22550 31780
rect 22838 31724 22876 31780
rect 22932 31724 22942 31780
rect 23426 31724 23436 31780
rect 23492 31724 23884 31780
rect 23940 31724 25452 31780
rect 25508 31724 25518 31780
rect 27570 31724 27580 31780
rect 27636 31724 28364 31780
rect 28420 31724 28430 31780
rect 11676 31612 12516 31668
rect 12572 31612 12582 31668
rect 13010 31612 13020 31668
rect 13076 31612 13916 31668
rect 13972 31612 15596 31668
rect 15652 31612 15662 31668
rect 20738 31612 20748 31668
rect 20804 31612 22092 31668
rect 22148 31612 22158 31668
rect 24434 31612 24444 31668
rect 24500 31612 25564 31668
rect 25620 31612 25630 31668
rect 11676 31444 11732 31612
rect 13020 31556 13076 31612
rect 30380 31556 30436 32060
rect 35756 32004 35812 32284
rect 38098 32172 38108 32228
rect 38164 32172 39676 32228
rect 39732 32172 39742 32228
rect 33058 31948 33068 32004
rect 33124 31948 35532 32004
rect 35588 31948 35598 32004
rect 35756 31948 38780 32004
rect 38836 31948 39452 32004
rect 39508 31948 39518 32004
rect 42018 31948 42028 32004
rect 42084 31948 42588 32004
rect 42644 31948 42654 32004
rect 44706 31948 44716 32004
rect 44772 31948 45220 32004
rect 45276 31948 45286 32004
rect 45714 31948 45724 32004
rect 45780 31948 48860 32004
rect 48916 31948 48926 32004
rect 50200 31892 51000 31920
rect 32162 31836 32172 31892
rect 32228 31836 34076 31892
rect 34132 31836 34142 31892
rect 38994 31836 39004 31892
rect 39060 31836 39564 31892
rect 39620 31836 39630 31892
rect 49634 31836 49644 31892
rect 49700 31836 51000 31892
rect 50200 31808 51000 31836
rect 12114 31500 12124 31556
rect 12180 31500 13076 31556
rect 20178 31500 20188 31556
rect 20244 31500 21812 31556
rect 21868 31500 21878 31556
rect 30370 31500 30380 31556
rect 30436 31500 30446 31556
rect 11666 31388 11676 31444
rect 11732 31388 11742 31444
rect 12338 31388 12348 31444
rect 12404 31388 13356 31444
rect 13412 31388 13422 31444
rect 32386 31388 32396 31444
rect 32452 31388 33404 31444
rect 33460 31388 33470 31444
rect 34178 31388 34188 31444
rect 34244 31388 35756 31444
rect 35812 31388 35822 31444
rect 44258 31388 44268 31444
rect 44324 31388 47908 31444
rect 47964 31388 47974 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 16706 31276 16716 31332
rect 16772 31276 17388 31332
rect 17444 31276 19684 31332
rect 26114 31276 26124 31332
rect 26180 31276 26628 31332
rect 26684 31276 29484 31332
rect 29540 31276 29550 31332
rect 46778 31276 46788 31332
rect 46844 31276 47180 31332
rect 47236 31276 47404 31332
rect 47460 31276 47470 31332
rect 19628 31220 19684 31276
rect 2370 31164 2380 31220
rect 2436 31164 4172 31220
rect 4228 31164 4956 31220
rect 5012 31164 5022 31220
rect 5394 31164 5404 31220
rect 5460 31164 6300 31220
rect 6356 31164 6366 31220
rect 14018 31164 14028 31220
rect 14084 31164 14924 31220
rect 14980 31164 15820 31220
rect 15876 31164 15886 31220
rect 16594 31164 16604 31220
rect 16660 31164 18620 31220
rect 18676 31164 18686 31220
rect 19628 31164 21196 31220
rect 21252 31164 21262 31220
rect 24770 31164 24780 31220
rect 24836 31164 25788 31220
rect 25844 31164 30380 31220
rect 30436 31164 30446 31220
rect 32386 31164 32396 31220
rect 32452 31164 38108 31220
rect 38164 31164 38780 31220
rect 38836 31164 38846 31220
rect 46162 31164 46172 31220
rect 46228 31164 47740 31220
rect 47796 31164 47806 31220
rect 4722 31052 4732 31108
rect 4788 31052 5684 31108
rect 5740 31052 5750 31108
rect 12506 31052 12516 31108
rect 12572 31052 15148 31108
rect 16034 31052 16044 31108
rect 16100 31052 18956 31108
rect 19012 31052 19022 31108
rect 19114 31052 19124 31108
rect 19180 31052 20412 31108
rect 20468 31052 20478 31108
rect 20850 31052 20860 31108
rect 20916 31052 22764 31108
rect 22820 31052 22830 31108
rect 33618 31052 33628 31108
rect 33684 31052 34748 31108
rect 34804 31052 38668 31108
rect 39218 31052 39228 31108
rect 39284 31052 40012 31108
rect 40068 31052 42252 31108
rect 42308 31052 42318 31108
rect 15092 30996 15148 31052
rect 38612 30996 38668 31052
rect 41244 30996 41300 31052
rect 4050 30940 4060 30996
rect 4116 30940 5404 30996
rect 5460 30940 5470 30996
rect 5842 30940 5852 30996
rect 5908 30940 7064 30996
rect 7120 30940 7130 30996
rect 13346 30940 13356 30996
rect 13412 30940 13524 30996
rect 13580 30940 14812 30996
rect 14868 30940 14878 30996
rect 15092 30940 19404 30996
rect 19460 30940 19470 30996
rect 19618 30940 19628 30996
rect 19684 30940 20188 30996
rect 20244 30940 20254 30996
rect 21130 30940 21140 30996
rect 21196 30940 22428 30996
rect 22484 30940 22494 30996
rect 24546 30940 24556 30996
rect 24612 30940 25788 30996
rect 25844 30940 26460 30996
rect 26516 30940 26526 30996
rect 27346 30940 27356 30996
rect 27412 30940 29036 30996
rect 29092 30940 29102 30996
rect 32274 30940 32284 30996
rect 32340 30940 32508 30996
rect 32564 30940 33516 30996
rect 33572 30940 33582 30996
rect 38612 30940 40908 30996
rect 40964 30940 40974 30996
rect 41234 30940 41244 30996
rect 41300 30940 41310 30996
rect 4274 30828 4284 30884
rect 4340 30828 5124 30884
rect 5180 30828 5516 30884
rect 5572 30828 5582 30884
rect 12674 30828 12684 30884
rect 12740 30828 13692 30884
rect 13748 30828 13758 30884
rect 18610 30828 18620 30884
rect 18676 30828 18844 30884
rect 18900 30828 18910 30884
rect 20626 30828 20636 30884
rect 20692 30828 22988 30884
rect 23044 30828 24668 30884
rect 24724 30828 24734 30884
rect 27738 30828 27748 30884
rect 27804 30828 28588 30884
rect 28644 30828 30044 30884
rect 30100 30828 30110 30884
rect 38994 30828 39004 30884
rect 39060 30828 41020 30884
rect 41076 30828 41086 30884
rect 43698 30828 43708 30884
rect 43764 30828 44940 30884
rect 44996 30828 45500 30884
rect 45556 30828 45566 30884
rect 13010 30716 13020 30772
rect 13076 30716 13916 30772
rect 13972 30716 13982 30772
rect 15092 30716 21644 30772
rect 21700 30716 21710 30772
rect 24770 30716 24780 30772
rect 24836 30716 25284 30772
rect 25340 30716 25350 30772
rect 35466 30716 35476 30772
rect 35532 30716 37996 30772
rect 38052 30716 38062 30772
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 15092 30436 15148 30716
rect 16818 30604 16828 30660
rect 16884 30604 17276 30660
rect 17332 30604 17342 30660
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 15474 30492 15484 30548
rect 15540 30492 16716 30548
rect 16772 30492 16782 30548
rect 17378 30492 17388 30548
rect 17444 30492 17724 30548
rect 17780 30492 17790 30548
rect 19058 30492 19068 30548
rect 19124 30492 20244 30548
rect 20402 30492 20412 30548
rect 20468 30492 22540 30548
rect 22596 30492 23268 30548
rect 23324 30492 23334 30548
rect 20188 30436 20244 30492
rect 13234 30380 13244 30436
rect 13300 30380 14588 30436
rect 14644 30380 15148 30436
rect 15204 30380 15214 30436
rect 16930 30380 16940 30436
rect 16996 30380 19348 30436
rect 19404 30380 19414 30436
rect 20188 30380 22596 30436
rect 22540 30324 22596 30380
rect 2930 30268 2940 30324
rect 2996 30268 4956 30324
rect 5012 30268 6188 30324
rect 6244 30268 6254 30324
rect 10658 30268 10668 30324
rect 10724 30268 11676 30324
rect 11732 30268 11742 30324
rect 17798 30268 17836 30324
rect 17892 30268 17902 30324
rect 20486 30268 20524 30324
rect 20580 30268 20590 30324
rect 22306 30268 22316 30324
rect 22372 30268 22382 30324
rect 22540 30268 23604 30324
rect 26618 30268 26628 30324
rect 26684 30268 26796 30324
rect 26852 30268 26862 30324
rect 33394 30268 33404 30324
rect 33460 30268 36876 30324
rect 36932 30268 36942 30324
rect 37874 30268 37884 30324
rect 37940 30268 38444 30324
rect 38500 30268 38510 30324
rect 22316 30212 22372 30268
rect 2818 30156 2828 30212
rect 2884 30156 5740 30212
rect 5796 30156 5806 30212
rect 6962 30156 6972 30212
rect 7028 30156 8316 30212
rect 8372 30156 8382 30212
rect 10994 30156 11004 30212
rect 11060 30156 12236 30212
rect 12292 30156 12302 30212
rect 17602 30156 17612 30212
rect 17668 30156 18172 30212
rect 18228 30156 18238 30212
rect 18386 30156 18396 30212
rect 18452 30156 19908 30212
rect 19964 30156 19974 30212
rect 21186 30156 21196 30212
rect 21252 30156 22372 30212
rect 23548 30212 23604 30268
rect 23548 30156 26012 30212
rect 26068 30156 26740 30212
rect 28130 30156 28140 30212
rect 28196 30156 28700 30212
rect 28756 30156 28766 30212
rect 33282 30156 33292 30212
rect 33348 30156 35308 30212
rect 35364 30156 35374 30212
rect 37426 30156 37436 30212
rect 37492 30156 38668 30212
rect 38724 30156 38892 30212
rect 38948 30156 38958 30212
rect 39218 30156 39228 30212
rect 39284 30156 39900 30212
rect 39956 30156 41356 30212
rect 41412 30156 41422 30212
rect 42914 30156 42924 30212
rect 42980 30156 43596 30212
rect 43652 30156 44716 30212
rect 44772 30156 45164 30212
rect 45220 30156 45230 30212
rect 46386 30156 46396 30212
rect 46452 30156 48524 30212
rect 48580 30156 48590 30212
rect 3938 30044 3948 30100
rect 4004 30044 5292 30100
rect 5348 30044 5358 30100
rect 6290 30044 6300 30100
rect 6356 30044 7084 30100
rect 7140 30044 7150 30100
rect 14074 30044 14084 30100
rect 14140 30044 15260 30100
rect 15316 30044 15820 30100
rect 15876 30044 15886 30100
rect 18274 30044 18284 30100
rect 18340 30044 19180 30100
rect 19236 30044 19246 30100
rect 4722 29932 4732 29988
rect 4788 29932 7532 29988
rect 7588 29932 7598 29988
rect 11442 29932 11452 29988
rect 11508 29932 15372 29988
rect 15428 29932 15708 29988
rect 15764 29932 15774 29988
rect 18610 29932 18620 29988
rect 18676 29932 19292 29988
rect 19348 29932 19358 29988
rect 19516 29876 19572 30156
rect 26684 30100 26740 30156
rect 26674 30044 26684 30100
rect 26740 30044 26750 30100
rect 34290 30044 34300 30100
rect 34356 30044 35532 30100
rect 35588 30044 35598 30100
rect 37650 30044 37660 30100
rect 37716 30044 39116 30100
rect 39172 30044 39182 30100
rect 40114 30044 40124 30100
rect 40180 30044 43260 30100
rect 43316 30044 43326 30100
rect 40124 29988 40180 30044
rect 47628 29988 47684 30156
rect 20066 29932 20076 29988
rect 20132 29932 21868 29988
rect 21924 29932 21934 29988
rect 31714 29932 31724 29988
rect 31780 29932 34972 29988
rect 35028 29932 35038 29988
rect 38882 29932 38892 29988
rect 38948 29932 40180 29988
rect 42690 29932 42700 29988
rect 42756 29932 43372 29988
rect 43428 29932 44492 29988
rect 44548 29932 44940 29988
rect 44996 29932 45006 29988
rect 47618 29932 47628 29988
rect 47684 29932 47694 29988
rect 5058 29820 5068 29876
rect 5124 29820 6860 29876
rect 6916 29820 6926 29876
rect 9090 29820 9100 29876
rect 9156 29820 9548 29876
rect 9604 29820 9614 29876
rect 12786 29820 12796 29876
rect 12852 29820 16940 29876
rect 16996 29820 17500 29876
rect 17556 29820 18844 29876
rect 18900 29820 18910 29876
rect 19394 29820 19404 29876
rect 19460 29820 19572 29876
rect 27794 29820 27804 29876
rect 27860 29820 28924 29876
rect 28980 29820 30604 29876
rect 30660 29820 31836 29876
rect 31892 29820 34076 29876
rect 34132 29820 34142 29876
rect 38322 29820 38332 29876
rect 38388 29820 44828 29876
rect 44884 29820 46228 29876
rect 46284 29820 48972 29876
rect 49028 29820 49038 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 5282 29708 5292 29764
rect 5348 29708 7196 29764
rect 7252 29708 7868 29764
rect 7924 29708 7934 29764
rect 31938 29708 31948 29764
rect 32004 29708 32732 29764
rect 32788 29708 32798 29764
rect 3826 29596 3836 29652
rect 3892 29596 5628 29652
rect 5684 29596 6636 29652
rect 6692 29596 6702 29652
rect 23538 29596 23548 29652
rect 23604 29596 24444 29652
rect 24500 29596 24510 29652
rect 26114 29596 26124 29652
rect 26180 29596 28588 29652
rect 28644 29596 28654 29652
rect 33562 29596 33572 29652
rect 33628 29596 34300 29652
rect 34356 29596 34366 29652
rect 35354 29596 35364 29652
rect 35420 29596 35980 29652
rect 36036 29596 38556 29652
rect 38612 29596 41468 29652
rect 41524 29596 42028 29652
rect 42084 29596 42094 29652
rect 9650 29484 9660 29540
rect 9716 29484 10444 29540
rect 10500 29484 10510 29540
rect 16370 29484 16380 29540
rect 16436 29484 21084 29540
rect 21140 29484 21150 29540
rect 36978 29484 36988 29540
rect 37044 29484 38220 29540
rect 38276 29484 44380 29540
rect 44436 29484 46452 29540
rect 46508 29484 48860 29540
rect 48916 29484 48926 29540
rect 8372 29372 9212 29428
rect 9268 29372 15932 29428
rect 15988 29372 16492 29428
rect 16548 29372 16828 29428
rect 16884 29372 16894 29428
rect 19618 29372 19628 29428
rect 19684 29372 19964 29428
rect 20020 29372 21420 29428
rect 21476 29372 21486 29428
rect 22530 29372 22540 29428
rect 22596 29372 22876 29428
rect 22932 29372 22942 29428
rect 25330 29372 25340 29428
rect 25396 29372 25676 29428
rect 25732 29372 27524 29428
rect 27580 29372 27590 29428
rect 33506 29372 33516 29428
rect 33572 29372 34300 29428
rect 34356 29372 34366 29428
rect 34626 29372 34636 29428
rect 34692 29372 35868 29428
rect 35924 29372 35934 29428
rect 36866 29372 36876 29428
rect 36932 29372 38556 29428
rect 38612 29372 41076 29428
rect 41132 29372 41142 29428
rect 48066 29372 48076 29428
rect 48132 29372 49084 29428
rect 49140 29372 49150 29428
rect 8372 29316 8428 29372
rect 7522 29260 7532 29316
rect 7588 29260 8428 29316
rect 8530 29260 8540 29316
rect 8596 29260 9996 29316
rect 10052 29260 10062 29316
rect 20962 29260 20972 29316
rect 21028 29260 23100 29316
rect 23156 29260 23166 29316
rect 27906 29260 27916 29316
rect 27972 29260 28364 29316
rect 28420 29260 33628 29316
rect 33684 29260 34188 29316
rect 34244 29260 34254 29316
rect 38770 29260 38780 29316
rect 38836 29260 39508 29316
rect 39452 29204 39508 29260
rect 12674 29148 12684 29204
rect 12740 29148 13356 29204
rect 13412 29148 13422 29204
rect 15250 29148 15260 29204
rect 15316 29148 23380 29204
rect 23436 29148 23446 29204
rect 26450 29148 26460 29204
rect 26516 29148 28476 29204
rect 28532 29148 28542 29204
rect 37762 29148 37772 29204
rect 37828 29148 39284 29204
rect 39340 29148 39350 29204
rect 39442 29148 39452 29204
rect 39508 29148 41020 29204
rect 41076 29148 41086 29204
rect 11554 29036 11564 29092
rect 11620 29036 11900 29092
rect 11956 29036 11966 29092
rect 21858 29036 21868 29092
rect 21924 29036 22316 29092
rect 22372 29036 22382 29092
rect 24434 29036 24444 29092
rect 24500 29036 30324 29092
rect 30380 29036 30390 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 18050 28924 18060 28980
rect 18116 28924 18396 28980
rect 18452 28924 18462 28980
rect 21298 28924 21308 28980
rect 21364 28924 23324 28980
rect 23380 28924 23390 28980
rect 26898 28924 26908 28980
rect 26964 28924 28140 28980
rect 28196 28924 28206 28980
rect 28466 28924 28476 28980
rect 28532 28924 29372 28980
rect 29428 28924 29438 28980
rect 38994 28924 39004 28980
rect 39060 28924 42140 28980
rect 42196 28924 42206 28980
rect 2930 28812 2940 28868
rect 2996 28812 5964 28868
rect 6020 28812 6030 28868
rect 10210 28812 10220 28868
rect 10276 28812 11396 28868
rect 11452 28812 12348 28868
rect 12404 28812 12414 28868
rect 15092 28812 16940 28868
rect 16996 28812 18508 28868
rect 18564 28812 18574 28868
rect 21522 28812 21532 28868
rect 21588 28812 24276 28868
rect 26226 28812 26236 28868
rect 26292 28812 26460 28868
rect 26516 28812 26526 28868
rect 28242 28812 28252 28868
rect 28308 28812 29708 28868
rect 29764 28812 31836 28868
rect 31892 28812 31902 28868
rect 33338 28812 33348 28868
rect 33404 28812 35644 28868
rect 35700 28812 35710 28868
rect 36026 28812 36036 28868
rect 36092 28812 36876 28868
rect 36932 28812 36942 28868
rect 41906 28812 41916 28868
rect 41972 28812 43932 28868
rect 43988 28812 43998 28868
rect 15092 28756 15148 28812
rect 4834 28700 4844 28756
rect 4900 28700 5740 28756
rect 5796 28700 5806 28756
rect 9202 28700 9212 28756
rect 9268 28700 9996 28756
rect 10052 28700 15148 28756
rect 16258 28700 16268 28756
rect 16324 28700 20300 28756
rect 20356 28700 20366 28756
rect 21410 28700 21420 28756
rect 21476 28700 22484 28756
rect 22428 28644 22484 28700
rect 24220 28644 24276 28812
rect 25722 28700 25732 28756
rect 25788 28700 26796 28756
rect 26852 28700 26862 28756
rect 28130 28700 28140 28756
rect 28196 28700 30940 28756
rect 30996 28700 32844 28756
rect 32900 28700 32910 28756
rect 33068 28700 33964 28756
rect 34020 28700 34030 28756
rect 35858 28700 35868 28756
rect 35924 28700 37884 28756
rect 37940 28700 37950 28756
rect 33068 28644 33124 28700
rect 1586 28588 1596 28644
rect 1652 28588 4060 28644
rect 4116 28588 5292 28644
rect 5348 28588 6972 28644
rect 7028 28588 7038 28644
rect 7970 28588 7980 28644
rect 8036 28588 10220 28644
rect 10276 28588 10286 28644
rect 11666 28588 11676 28644
rect 11732 28588 12236 28644
rect 12292 28588 12302 28644
rect 13234 28588 13244 28644
rect 13300 28588 13692 28644
rect 13748 28588 13758 28644
rect 14466 28588 14476 28644
rect 14532 28588 14812 28644
rect 14868 28588 14878 28644
rect 15260 28588 15932 28644
rect 15988 28588 15998 28644
rect 17714 28588 17724 28644
rect 17780 28588 18060 28644
rect 18116 28588 18126 28644
rect 22418 28588 22428 28644
rect 22484 28588 22494 28644
rect 24210 28588 24220 28644
rect 24276 28588 25956 28644
rect 26114 28588 26124 28644
rect 26180 28588 27132 28644
rect 27188 28588 27198 28644
rect 27356 28588 27636 28644
rect 27692 28588 27702 28644
rect 28802 28588 28812 28644
rect 28868 28588 29484 28644
rect 29540 28588 33068 28644
rect 33124 28588 33134 28644
rect 33506 28588 33516 28644
rect 33572 28588 34524 28644
rect 34580 28588 34590 28644
rect 36474 28588 36484 28644
rect 36540 28588 36988 28644
rect 37044 28588 37212 28644
rect 37268 28588 37278 28644
rect 37436 28588 37548 28644
rect 37604 28588 37614 28644
rect 38210 28588 38220 28644
rect 38276 28588 38892 28644
rect 38948 28588 38958 28644
rect 40236 28588 40796 28644
rect 40852 28588 40862 28644
rect 2706 28476 2716 28532
rect 2772 28476 3612 28532
rect 3668 28476 3678 28532
rect 11890 28476 11900 28532
rect 11956 28476 12460 28532
rect 12516 28476 12526 28532
rect 5954 28252 5964 28308
rect 6020 28252 6188 28308
rect 6244 28252 7252 28308
rect 7308 28252 7318 28308
rect 14802 28140 14812 28196
rect 14868 28140 15036 28196
rect 15092 28140 15102 28196
rect 15260 27972 15316 28588
rect 25900 28532 25956 28588
rect 25900 28476 26012 28532
rect 26068 28476 26078 28532
rect 26226 28476 26236 28532
rect 26292 28476 26684 28532
rect 26740 28476 26750 28532
rect 26758 28364 26796 28420
rect 26852 28364 26862 28420
rect 27356 28308 27412 28588
rect 37436 28532 37492 28588
rect 36866 28476 36876 28532
rect 36932 28476 37492 28532
rect 40236 28420 40292 28588
rect 42140 28420 42196 28812
rect 43138 28588 43148 28644
rect 43204 28588 44604 28644
rect 44660 28588 45500 28644
rect 45556 28588 45566 28644
rect 28914 28364 28924 28420
rect 28980 28364 32620 28420
rect 32676 28364 32686 28420
rect 33842 28364 33852 28420
rect 33908 28364 34972 28420
rect 35028 28364 35038 28420
rect 36754 28364 36764 28420
rect 36820 28364 38332 28420
rect 38388 28364 38398 28420
rect 40226 28364 40236 28420
rect 40292 28364 40302 28420
rect 42130 28364 42140 28420
rect 42196 28364 42206 28420
rect 26674 28252 26684 28308
rect 26740 28252 27412 28308
rect 34234 28252 34244 28308
rect 34300 28252 39004 28308
rect 39060 28252 39070 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 29026 28140 29036 28196
rect 29092 28140 29372 28196
rect 29428 28140 29438 28196
rect 30034 28140 30044 28196
rect 30100 28140 31164 28196
rect 31220 28140 32508 28196
rect 32564 28140 32574 28196
rect 17826 28028 17836 28084
rect 17892 28028 18284 28084
rect 18340 28028 20412 28084
rect 20468 28028 20478 28084
rect 27906 28028 27916 28084
rect 27972 28028 36148 28084
rect 36204 28028 37436 28084
rect 37492 28028 37502 28084
rect 37874 28028 37884 28084
rect 37940 28028 38332 28084
rect 38388 28028 38398 28084
rect 41066 28028 41076 28084
rect 41132 28028 42644 28084
rect 42700 28028 47628 28084
rect 47684 28028 47694 28084
rect 8978 27916 8988 27972
rect 9044 27916 9884 27972
rect 9940 27916 9950 27972
rect 14354 27916 14364 27972
rect 14420 27916 15036 27972
rect 15092 27916 15316 27972
rect 19618 27916 19628 27972
rect 19684 27916 20524 27972
rect 20580 27916 20590 27972
rect 30370 27916 30380 27972
rect 30436 27916 31388 27972
rect 31444 27916 31454 27972
rect 37772 27916 39150 27972
rect 39206 27916 39216 27972
rect 37772 27860 37828 27916
rect 3826 27804 3836 27860
rect 3892 27804 4284 27860
rect 4340 27804 4350 27860
rect 6738 27804 6748 27860
rect 6804 27804 7084 27860
rect 7140 27804 7150 27860
rect 9314 27804 9324 27860
rect 9380 27804 14028 27860
rect 14084 27804 14094 27860
rect 16034 27804 16044 27860
rect 16100 27804 17052 27860
rect 17108 27804 17118 27860
rect 18050 27804 18060 27860
rect 18116 27804 18732 27860
rect 18788 27804 18798 27860
rect 19954 27804 19964 27860
rect 20020 27804 20860 27860
rect 20916 27804 21644 27860
rect 21700 27804 21710 27860
rect 22418 27804 22428 27860
rect 22484 27804 23436 27860
rect 23492 27804 23502 27860
rect 31266 27804 31276 27860
rect 31332 27804 32060 27860
rect 32116 27804 32126 27860
rect 33394 27804 33404 27860
rect 33460 27804 33740 27860
rect 33796 27804 33806 27860
rect 37762 27804 37772 27860
rect 37828 27804 37838 27860
rect 38434 27804 38444 27860
rect 38500 27804 39004 27860
rect 39060 27804 39070 27860
rect 41346 27804 41356 27860
rect 41412 27804 42812 27860
rect 42868 27804 44716 27860
rect 44772 27804 44782 27860
rect 33404 27748 33460 27804
rect 37772 27748 37828 27804
rect 6066 27692 6076 27748
rect 6132 27692 25396 27748
rect 25452 27692 25676 27748
rect 25732 27692 25742 27748
rect 30818 27692 30828 27748
rect 30884 27692 31612 27748
rect 31668 27692 33460 27748
rect 33842 27692 33852 27748
rect 33908 27692 35084 27748
rect 35140 27692 37828 27748
rect 50200 27636 51000 27664
rect 18050 27580 18060 27636
rect 18116 27580 27916 27636
rect 27972 27580 27982 27636
rect 37258 27580 37268 27636
rect 37324 27580 38108 27636
rect 38164 27580 38174 27636
rect 49298 27580 49308 27636
rect 49364 27580 51000 27636
rect 50200 27552 51000 27580
rect 11666 27468 11676 27524
rect 11732 27468 14980 27524
rect 21970 27468 21980 27524
rect 22036 27468 22744 27524
rect 22800 27468 22810 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 11330 27356 11340 27412
rect 11396 27356 11900 27412
rect 11956 27356 12460 27412
rect 12516 27356 14028 27412
rect 14084 27356 14094 27412
rect 14924 27300 14980 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 15138 27356 15148 27412
rect 15204 27356 16324 27412
rect 16380 27356 16390 27412
rect 18946 27356 18956 27412
rect 19012 27356 19516 27412
rect 19572 27356 19582 27412
rect 12842 27244 12852 27300
rect 12908 27244 14700 27300
rect 14756 27244 14766 27300
rect 14924 27244 15596 27300
rect 15652 27244 15820 27300
rect 15876 27244 15886 27300
rect 17378 27244 17388 27300
rect 17444 27244 17612 27300
rect 17668 27244 17678 27300
rect 17826 27244 17836 27300
rect 17892 27244 18340 27300
rect 18396 27244 27804 27300
rect 27860 27244 27870 27300
rect 29698 27244 29708 27300
rect 29764 27244 30772 27300
rect 30828 27244 30838 27300
rect 37426 27244 37436 27300
rect 37492 27244 38220 27300
rect 38276 27244 38286 27300
rect 10098 27132 10108 27188
rect 10164 27132 13468 27188
rect 13524 27132 13534 27188
rect 17490 27132 17500 27188
rect 17556 27132 17668 27188
rect 23090 27132 23100 27188
rect 23156 27132 24220 27188
rect 24276 27132 24286 27188
rect 28578 27132 28588 27188
rect 28644 27132 32340 27188
rect 32396 27132 32406 27188
rect 37314 27132 37324 27188
rect 37380 27132 37884 27188
rect 37940 27132 37950 27188
rect 38098 27132 38108 27188
rect 38164 27132 38780 27188
rect 38836 27132 38846 27188
rect 40786 27132 40796 27188
rect 40852 27132 41916 27188
rect 41972 27132 41982 27188
rect 48234 27132 48244 27188
rect 48300 27132 49308 27188
rect 49364 27132 49374 27188
rect 4778 27020 4788 27076
rect 4844 27020 5628 27076
rect 5684 27020 5694 27076
rect 10882 27020 10892 27076
rect 10948 27020 11788 27076
rect 11844 27020 11854 27076
rect 12562 27020 12572 27076
rect 12628 27020 13300 27076
rect 13356 27020 13804 27076
rect 13860 27020 13870 27076
rect 10892 26964 10948 27020
rect 8316 26908 9660 26964
rect 9716 26908 9726 26964
rect 10332 26908 10948 26964
rect 11946 26908 11956 26964
rect 12012 26908 13580 26964
rect 13636 26908 13646 26964
rect 16258 26908 16268 26964
rect 16324 26908 17388 26964
rect 17444 26908 17454 26964
rect 8316 26852 8372 26908
rect 2594 26796 2604 26852
rect 2660 26796 5404 26852
rect 5460 26796 5470 26852
rect 8306 26796 8316 26852
rect 8372 26796 8382 26852
rect 10266 26796 10276 26852
rect 10332 26796 10388 26908
rect 17612 26740 17668 27132
rect 25452 27020 27356 27076
rect 27412 27020 27422 27076
rect 28074 27020 28084 27076
rect 28140 27020 29036 27076
rect 29092 27020 29102 27076
rect 31826 27020 31836 27076
rect 31892 27020 32620 27076
rect 32676 27020 33292 27076
rect 33348 27020 33516 27076
rect 33572 27020 34188 27076
rect 34244 27020 34254 27076
rect 34458 27020 34468 27076
rect 34524 27020 34748 27076
rect 34804 27020 34814 27076
rect 36978 27020 36988 27076
rect 37044 27020 37660 27076
rect 37716 27020 37726 27076
rect 37986 27020 37996 27076
rect 38052 27020 41132 27076
rect 41188 27020 41198 27076
rect 25452 26852 25508 27020
rect 26002 26908 26012 26964
rect 26068 26908 27020 26964
rect 27076 26908 27086 26964
rect 28364 26908 29372 26964
rect 29428 26908 29438 26964
rect 34066 26908 34076 26964
rect 34132 26908 35084 26964
rect 35140 26908 35150 26964
rect 36474 26908 36484 26964
rect 36540 26908 39004 26964
rect 39060 26908 39070 26964
rect 46284 26908 47404 26964
rect 47460 26908 47470 26964
rect 28364 26852 28420 26908
rect 46284 26852 46340 26908
rect 19170 26796 19180 26852
rect 19236 26796 21532 26852
rect 21588 26796 22372 26852
rect 25442 26796 25452 26852
rect 25508 26796 25518 26852
rect 28354 26796 28364 26852
rect 28420 26796 28430 26852
rect 33842 26796 33852 26852
rect 33908 26796 34300 26852
rect 34356 26796 34366 26852
rect 35858 26796 35868 26852
rect 35924 26796 37212 26852
rect 37268 26796 37278 26852
rect 46274 26796 46284 26852
rect 46340 26796 46350 26852
rect 22316 26740 22372 26796
rect 17602 26684 17612 26740
rect 17668 26684 17678 26740
rect 22306 26684 22316 26740
rect 22372 26684 22382 26740
rect 34178 26684 34188 26740
rect 34244 26684 34860 26740
rect 34916 26684 34926 26740
rect 36978 26684 36988 26740
rect 37044 26684 37604 26740
rect 37660 26684 37670 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 6402 26572 6412 26628
rect 6468 26572 6972 26628
rect 7028 26572 7038 26628
rect 11106 26572 11116 26628
rect 11172 26572 11788 26628
rect 11844 26572 11854 26628
rect 25330 26572 25340 26628
rect 25396 26572 25900 26628
rect 25956 26572 25966 26628
rect 31378 26572 31388 26628
rect 31444 26572 38108 26628
rect 38164 26572 38174 26628
rect 10434 26460 10444 26516
rect 10500 26460 11228 26516
rect 11284 26460 11452 26516
rect 11508 26460 11518 26516
rect 13682 26460 13692 26516
rect 13748 26460 15764 26516
rect 15820 26460 16604 26516
rect 16660 26460 16670 26516
rect 17154 26460 17164 26516
rect 17220 26460 17500 26516
rect 17556 26460 17566 26516
rect 37426 26460 37436 26516
rect 37492 26460 38780 26516
rect 38836 26460 39340 26516
rect 39396 26460 39406 26516
rect 22754 26348 22764 26404
rect 22820 26348 25788 26404
rect 25844 26348 25854 26404
rect 31042 26348 31052 26404
rect 31108 26348 32284 26404
rect 32340 26348 32350 26404
rect 39106 26348 39116 26404
rect 39172 26348 39182 26404
rect 39890 26348 39900 26404
rect 39956 26348 43820 26404
rect 43876 26348 44044 26404
rect 44100 26348 45108 26404
rect 45164 26348 45174 26404
rect 39116 26292 39172 26348
rect 5142 26236 5180 26292
rect 5236 26236 5246 26292
rect 9986 26236 9996 26292
rect 10052 26236 11508 26292
rect 11564 26236 11574 26292
rect 24714 26236 24724 26292
rect 24780 26236 25228 26292
rect 25284 26236 25294 26292
rect 27794 26236 27804 26292
rect 27860 26236 31724 26292
rect 31780 26236 34076 26292
rect 34132 26236 34142 26292
rect 37762 26236 37772 26292
rect 37828 26236 38668 26292
rect 38724 26236 39452 26292
rect 39508 26236 39518 26292
rect 44930 26236 44940 26292
rect 44996 26236 46116 26292
rect 46172 26236 46182 26292
rect 46610 26236 46620 26292
rect 46676 26236 47628 26292
rect 47684 26236 47694 26292
rect 3154 26124 3164 26180
rect 3220 26124 3724 26180
rect 3780 26124 3790 26180
rect 6178 26124 6188 26180
rect 6244 26124 6860 26180
rect 6916 26124 6926 26180
rect 11218 26124 11228 26180
rect 11284 26124 14364 26180
rect 14420 26124 14430 26180
rect 16650 26124 16660 26180
rect 16716 26124 24276 26180
rect 24332 26124 27020 26180
rect 27076 26124 27916 26180
rect 27972 26124 27982 26180
rect 42018 26124 42028 26180
rect 42084 26124 42532 26180
rect 42588 26124 43036 26180
rect 43092 26124 43102 26180
rect 17714 26012 17724 26068
rect 17780 26012 18284 26068
rect 18340 26012 18350 26068
rect 33562 26012 33572 26068
rect 33628 26012 35084 26068
rect 35140 26012 35150 26068
rect 18498 25900 18508 25956
rect 18564 25900 20188 25956
rect 20244 25900 20254 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 30594 25788 30604 25844
rect 30660 25788 31164 25844
rect 31220 25788 31230 25844
rect 44314 25788 44324 25844
rect 44380 25788 46732 25844
rect 46788 25788 46798 25844
rect 47842 25788 47852 25844
rect 47908 25788 47918 25844
rect 19842 25676 19852 25732
rect 19908 25676 20300 25732
rect 20356 25676 20366 25732
rect 38938 25676 38948 25732
rect 39004 25676 39564 25732
rect 39620 25676 39630 25732
rect 19170 25564 19180 25620
rect 19236 25564 19628 25620
rect 19684 25564 19694 25620
rect 22754 25564 22764 25620
rect 22820 25564 23436 25620
rect 23492 25564 23502 25620
rect 44828 25508 44884 25788
rect 4498 25452 4508 25508
rect 4564 25452 7980 25508
rect 8036 25452 8316 25508
rect 8372 25452 8382 25508
rect 26114 25452 26124 25508
rect 26180 25452 26348 25508
rect 26404 25452 27580 25508
rect 27636 25452 29036 25508
rect 29092 25452 29102 25508
rect 34738 25452 34748 25508
rect 34804 25452 35308 25508
rect 35364 25452 35374 25508
rect 35578 25452 35588 25508
rect 35644 25452 35868 25508
rect 35924 25452 35934 25508
rect 37734 25452 37772 25508
rect 37828 25452 37838 25508
rect 38658 25452 38668 25508
rect 38724 25452 41916 25508
rect 41972 25452 43464 25508
rect 43520 25452 43530 25508
rect 44818 25452 44828 25508
rect 44884 25452 44894 25508
rect 5730 25340 5740 25396
rect 5796 25340 6412 25396
rect 6468 25340 6636 25396
rect 6692 25340 6702 25396
rect 28914 25340 28924 25396
rect 28980 25340 30044 25396
rect 30100 25340 30110 25396
rect 30930 25340 30940 25396
rect 30996 25340 32508 25396
rect 32564 25340 33516 25396
rect 33572 25340 34916 25396
rect 34972 25340 34982 25396
rect 40002 25340 40012 25396
rect 40068 25340 42588 25396
rect 42644 25340 42654 25396
rect 42588 25284 42644 25340
rect 5394 25228 5404 25284
rect 5460 25228 6076 25284
rect 6132 25228 7196 25284
rect 7252 25228 7262 25284
rect 12338 25228 12348 25284
rect 12404 25228 12852 25284
rect 12908 25228 13356 25284
rect 13412 25228 13422 25284
rect 30706 25228 30716 25284
rect 30772 25228 31052 25284
rect 31108 25228 32340 25284
rect 32396 25228 32406 25284
rect 33170 25228 33180 25284
rect 33236 25228 35308 25284
rect 35364 25228 35374 25284
rect 37762 25228 37772 25284
rect 37828 25228 38108 25284
rect 38164 25228 38174 25284
rect 38322 25228 38332 25284
rect 38388 25228 38668 25284
rect 38724 25228 38734 25284
rect 40282 25228 40292 25284
rect 40348 25228 41132 25284
rect 41188 25228 41198 25284
rect 42588 25228 44716 25284
rect 44772 25228 44782 25284
rect 43820 25172 43876 25228
rect 47852 25172 47908 25788
rect 10658 25116 10668 25172
rect 10724 25116 12012 25172
rect 12068 25116 12236 25172
rect 12292 25116 14140 25172
rect 14196 25116 14206 25172
rect 17042 25116 17052 25172
rect 17108 25116 17612 25172
rect 17668 25116 17678 25172
rect 26786 25116 26796 25172
rect 26852 25116 27244 25172
rect 27300 25116 27310 25172
rect 29474 25116 29484 25172
rect 29540 25116 30044 25172
rect 30100 25116 35756 25172
rect 35812 25116 35822 25172
rect 38770 25116 38780 25172
rect 38836 25116 39788 25172
rect 39844 25116 39854 25172
rect 43810 25116 43820 25172
rect 43876 25116 43886 25172
rect 44556 25116 44566 25172
rect 44622 25116 45612 25172
rect 45668 25116 47068 25172
rect 47124 25116 47134 25172
rect 47618 25116 47628 25172
rect 47684 25116 47908 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 4834 25004 4844 25060
rect 4900 25004 6188 25060
rect 6244 25004 6524 25060
rect 6580 25004 6590 25060
rect 10882 25004 10892 25060
rect 10948 25004 12460 25060
rect 12516 25004 13244 25060
rect 13300 25004 13804 25060
rect 13860 25004 15260 25060
rect 15316 25004 15326 25060
rect 25890 25004 25900 25060
rect 25956 25004 26572 25060
rect 26628 25004 26638 25060
rect 6290 24892 6300 24948
rect 6356 24892 7308 24948
rect 7364 24892 7374 24948
rect 12002 24892 12012 24948
rect 12068 24892 12572 24948
rect 12628 24892 12638 24948
rect 23090 24892 23100 24948
rect 23156 24892 23884 24948
rect 23940 24892 23950 24948
rect 25442 24892 25452 24948
rect 25508 24892 26684 24948
rect 26740 24892 26750 24948
rect 29922 24892 29932 24948
rect 29988 24892 32956 24948
rect 33012 24892 33180 24948
rect 33236 24892 33246 24948
rect 36194 24892 36204 24948
rect 36260 24892 37212 24948
rect 37268 24892 37278 24948
rect 3490 24780 3500 24836
rect 3556 24780 3948 24836
rect 4004 24780 4014 24836
rect 4554 24780 4564 24836
rect 4620 24780 4956 24836
rect 5012 24780 5852 24836
rect 5908 24780 5918 24836
rect 10994 24780 11004 24836
rect 11060 24780 11676 24836
rect 11732 24780 11742 24836
rect 14466 24780 14476 24836
rect 14532 24780 15596 24836
rect 15652 24780 24220 24836
rect 24276 24780 24286 24836
rect 30930 24780 30940 24836
rect 30996 24780 31164 24836
rect 31220 24780 31230 24836
rect 31397 24780 31407 24836
rect 31463 24780 32788 24836
rect 32844 24780 32854 24836
rect 45378 24780 45388 24836
rect 45444 24780 45836 24836
rect 45892 24780 47628 24836
rect 47684 24780 47694 24836
rect 1810 24668 1820 24724
rect 1876 24668 2268 24724
rect 2324 24668 2828 24724
rect 2884 24668 2894 24724
rect 9090 24668 9100 24724
rect 9156 24668 10164 24724
rect 10220 24668 10230 24724
rect 11330 24668 11340 24724
rect 11396 24668 14700 24724
rect 14756 24668 14766 24724
rect 20402 24668 20412 24724
rect 20468 24668 21756 24724
rect 21812 24668 21822 24724
rect 31266 24668 31276 24724
rect 31332 24668 31612 24724
rect 31668 24668 32284 24724
rect 32340 24668 32350 24724
rect 34066 24668 34076 24724
rect 34132 24668 34636 24724
rect 34692 24668 34702 24724
rect 34906 24668 34916 24724
rect 34972 24668 38220 24724
rect 38276 24668 38286 24724
rect 43698 24668 43708 24724
rect 43764 24668 44380 24724
rect 44436 24668 44446 24724
rect 47394 24668 47404 24724
rect 47460 24668 48860 24724
rect 48916 24668 48926 24724
rect 23762 24556 23772 24612
rect 23828 24556 24444 24612
rect 24500 24556 27132 24612
rect 27188 24556 27198 24612
rect 16706 24444 16716 24500
rect 16772 24444 17500 24500
rect 17556 24444 17566 24500
rect 18554 24444 18564 24500
rect 18620 24444 18844 24500
rect 18900 24444 18910 24500
rect 28522 24444 28532 24500
rect 28588 24444 29708 24500
rect 29764 24444 29774 24500
rect 33506 24444 33516 24500
rect 33572 24444 42140 24500
rect 42196 24444 42532 24500
rect 42476 24388 42532 24444
rect 12338 24332 12348 24388
rect 12404 24332 13468 24388
rect 13524 24332 13916 24388
rect 13972 24332 13982 24388
rect 15092 24332 34580 24388
rect 34636 24332 34646 24388
rect 42466 24332 42476 24388
rect 42532 24332 42542 24388
rect 47954 24332 47964 24388
rect 48020 24332 48748 24388
rect 48804 24332 48814 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 15092 24164 15148 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 15978 24220 15988 24276
rect 16044 24220 17724 24276
rect 17780 24220 17790 24276
rect 25890 24220 25900 24276
rect 25956 24220 34860 24276
rect 34916 24220 34972 24276
rect 35028 24220 35038 24276
rect 13906 24108 13916 24164
rect 13972 24108 15148 24164
rect 16986 24108 16996 24164
rect 17052 24108 18284 24164
rect 18340 24108 18350 24164
rect 26674 24108 26684 24164
rect 26740 24108 27244 24164
rect 27300 24108 37100 24164
rect 37156 24108 37166 24164
rect 37324 24108 37772 24164
rect 37828 24108 38556 24164
rect 38612 24108 39172 24164
rect 39228 24108 39238 24164
rect 37324 24052 37380 24108
rect 11666 23996 11676 24052
rect 11732 23996 12460 24052
rect 12516 23996 13580 24052
rect 13636 23996 13646 24052
rect 17602 23996 17612 24052
rect 17668 23996 22671 24052
rect 22727 23996 22737 24052
rect 25218 23996 25228 24052
rect 25284 23996 25732 24052
rect 25788 23996 25798 24052
rect 25900 23996 28140 24052
rect 28196 23996 28206 24052
rect 32610 23996 32620 24052
rect 32676 23996 34076 24052
rect 34132 23996 34142 24052
rect 35420 23996 37380 24052
rect 38434 23996 38444 24052
rect 38500 23996 39564 24052
rect 39620 23996 40236 24052
rect 40292 23996 40302 24052
rect 25900 23940 25956 23996
rect 35420 23940 35476 23996
rect 12226 23884 12236 23940
rect 12292 23884 12572 23940
rect 12628 23884 12638 23940
rect 12786 23884 12796 23940
rect 12852 23884 13244 23940
rect 13300 23884 13310 23940
rect 16594 23884 16604 23940
rect 16660 23884 17948 23940
rect 18004 23884 18956 23940
rect 19012 23884 20412 23940
rect 20468 23884 20478 23940
rect 22418 23884 22428 23940
rect 22484 23884 24220 23940
rect 24276 23884 24286 23940
rect 24434 23884 24444 23940
rect 24500 23884 25956 23940
rect 26562 23884 26572 23940
rect 26628 23884 27356 23940
rect 27412 23884 27422 23940
rect 28242 23884 28252 23940
rect 28308 23884 31164 23940
rect 31220 23884 31230 23940
rect 34570 23884 34580 23940
rect 34636 23884 35420 23940
rect 35476 23884 35486 23940
rect 37986 23884 37996 23940
rect 38052 23884 39452 23940
rect 39508 23884 41356 23940
rect 41412 23884 41422 23940
rect 42970 23884 42980 23940
rect 43036 23884 46732 23940
rect 46788 23884 47180 23940
rect 47236 23884 47246 23940
rect 47618 23884 47628 23940
rect 47684 23884 48188 23940
rect 48244 23884 48580 23940
rect 48636 23884 48646 23940
rect 11106 23772 11116 23828
rect 11172 23772 11732 23828
rect 11788 23772 12908 23828
rect 12964 23772 12974 23828
rect 13122 23772 13132 23828
rect 13188 23772 15988 23828
rect 16044 23772 16054 23828
rect 16370 23772 16380 23828
rect 16436 23772 17388 23828
rect 17444 23772 17454 23828
rect 17546 23772 17556 23828
rect 17612 23772 18284 23828
rect 18340 23772 18350 23828
rect 34738 23772 34748 23828
rect 34804 23772 38332 23828
rect 38388 23772 38398 23828
rect 44202 23772 44212 23828
rect 44268 23772 44828 23828
rect 44884 23772 44894 23828
rect 12908 23716 12964 23772
rect 12908 23660 21420 23716
rect 21476 23660 21486 23716
rect 25218 23660 25228 23716
rect 25284 23660 34860 23716
rect 34916 23660 34926 23716
rect 18722 23548 18732 23604
rect 18788 23548 19292 23604
rect 19348 23548 19358 23604
rect 26852 23548 27188 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 26684 23492 26908 23548
rect 3938 23436 3948 23492
rect 4004 23436 4284 23492
rect 4340 23436 5180 23492
rect 5236 23436 5628 23492
rect 5684 23436 5694 23492
rect 13346 23436 13356 23492
rect 13412 23436 14252 23492
rect 14308 23436 14318 23492
rect 26338 23436 26348 23492
rect 26404 23436 26740 23492
rect 27132 23380 27188 23548
rect 28130 23436 28140 23492
rect 28196 23436 28588 23492
rect 28644 23436 28654 23492
rect 29586 23436 29596 23492
rect 29652 23436 30380 23492
rect 30436 23436 31724 23492
rect 31780 23436 31790 23492
rect 34906 23436 34916 23492
rect 35028 23436 35038 23492
rect 35298 23436 35308 23492
rect 35364 23436 36372 23492
rect 36428 23436 38668 23492
rect 2482 23324 2492 23380
rect 2548 23324 9660 23380
rect 9716 23324 9726 23380
rect 13178 23324 13188 23380
rect 13244 23324 13916 23380
rect 13972 23324 13982 23380
rect 18778 23324 18788 23380
rect 18844 23324 21084 23380
rect 21140 23324 21150 23380
rect 27132 23324 29820 23380
rect 29876 23324 32172 23380
rect 32228 23324 32238 23380
rect 32396 23324 32956 23380
rect 33012 23324 33022 23380
rect 34458 23324 34468 23380
rect 34524 23324 35084 23380
rect 35140 23324 36988 23380
rect 37044 23324 37054 23380
rect 32396 23268 32452 23324
rect 5338 23212 5348 23268
rect 5404 23212 5516 23268
rect 5572 23212 6636 23268
rect 6692 23212 6702 23268
rect 11386 23212 11396 23268
rect 11452 23212 14588 23268
rect 14644 23212 14654 23268
rect 17266 23212 17276 23268
rect 17332 23212 17612 23268
rect 17668 23212 17678 23268
rect 18330 23212 18340 23268
rect 18396 23212 20916 23268
rect 20972 23212 20982 23268
rect 26450 23212 26460 23268
rect 26516 23212 30044 23268
rect 30100 23212 32396 23268
rect 32452 23212 32462 23268
rect 32610 23212 32620 23268
rect 32676 23212 33572 23268
rect 33516 23156 33572 23212
rect 2706 23100 2716 23156
rect 2772 23100 3612 23156
rect 3668 23100 3678 23156
rect 6850 23100 6860 23156
rect 6916 23100 10836 23156
rect 10892 23100 13020 23156
rect 13076 23100 13086 23156
rect 15474 23100 15484 23156
rect 15540 23100 16156 23156
rect 16212 23100 19908 23156
rect 19964 23100 19974 23156
rect 24770 23100 24780 23156
rect 24836 23100 25732 23156
rect 25788 23100 25798 23156
rect 26002 23100 26012 23156
rect 26068 23100 27020 23156
rect 27076 23100 27086 23156
rect 28690 23100 28700 23156
rect 28756 23100 29708 23156
rect 29764 23100 29774 23156
rect 31658 23100 31668 23156
rect 31724 23100 32956 23156
rect 33012 23100 33022 23156
rect 33506 23100 33516 23156
rect 33572 23100 33908 23156
rect 33964 23100 37324 23156
rect 37380 23100 38444 23156
rect 38500 23100 38510 23156
rect 38612 23100 38668 23436
rect 50200 23380 51000 23408
rect 39666 23324 39676 23380
rect 39732 23324 40404 23380
rect 40460 23324 40470 23380
rect 40898 23324 40908 23380
rect 40964 23324 44940 23380
rect 44996 23324 45006 23380
rect 49410 23324 49420 23380
rect 49476 23324 51000 23380
rect 50200 23296 51000 23324
rect 44538 23212 44548 23268
rect 44604 23212 45948 23268
rect 46004 23212 46014 23268
rect 38724 23100 40124 23156
rect 40180 23100 40190 23156
rect 41906 23100 41916 23156
rect 41972 23100 45388 23156
rect 45444 23100 45454 23156
rect 47730 23100 47740 23156
rect 47796 23100 48636 23156
rect 48692 23100 48702 23156
rect 17714 22988 17724 23044
rect 17780 22988 18172 23044
rect 18228 22988 18238 23044
rect 20626 22988 20636 23044
rect 20692 22988 21084 23044
rect 21140 22988 26796 23044
rect 26852 22988 26862 23044
rect 31154 22988 31164 23044
rect 31220 22988 31948 23044
rect 32004 22988 32014 23044
rect 35298 22988 35308 23044
rect 35364 22988 35868 23044
rect 35924 22988 35934 23044
rect 36978 22988 36988 23044
rect 37044 22988 37436 23044
rect 37492 22988 38220 23044
rect 38276 22988 39956 23044
rect 40012 22988 43484 23044
rect 43540 22988 43550 23044
rect 46162 22988 46172 23044
rect 46228 22988 48972 23044
rect 49028 22988 49038 23044
rect 10882 22876 10892 22932
rect 10948 22876 11732 22932
rect 11788 22876 11798 22932
rect 14690 22876 14700 22932
rect 14756 22876 27804 22932
rect 27860 22876 27870 22932
rect 30874 22876 30884 22932
rect 30940 22876 31500 22932
rect 31556 22876 31566 22932
rect 34972 22876 35420 22932
rect 35476 22876 35486 22932
rect 37314 22876 37324 22932
rect 37380 22876 42028 22932
rect 42084 22876 42094 22932
rect 44034 22876 44044 22932
rect 44100 22876 45108 22932
rect 45164 22876 45174 22932
rect 34972 22820 35028 22876
rect 14578 22764 14588 22820
rect 14644 22764 35028 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 15250 22652 15260 22708
rect 15316 22652 22484 22708
rect 22540 22652 22550 22708
rect 41010 22652 41020 22708
rect 41076 22652 41468 22708
rect 41524 22652 41534 22708
rect 3434 22540 3444 22596
rect 3500 22540 5068 22596
rect 5124 22540 5134 22596
rect 27906 22540 27916 22596
rect 27972 22540 28476 22596
rect 28532 22540 30548 22596
rect 30604 22540 30614 22596
rect 40338 22540 40348 22596
rect 40404 22540 41244 22596
rect 41300 22540 44492 22596
rect 44548 22540 45724 22596
rect 45780 22540 46732 22596
rect 46788 22540 46798 22596
rect 12450 22428 12460 22484
rect 12516 22428 12852 22484
rect 27794 22428 27804 22484
rect 27860 22428 29316 22484
rect 29372 22428 29932 22484
rect 29988 22428 29998 22484
rect 34066 22428 34076 22484
rect 34132 22428 34636 22484
rect 34692 22428 35644 22484
rect 35700 22428 35710 22484
rect 38882 22428 38892 22484
rect 38948 22428 40908 22484
rect 40964 22428 40974 22484
rect 12796 22372 12852 22428
rect 5842 22316 5852 22372
rect 5908 22316 7868 22372
rect 7924 22316 8876 22372
rect 8932 22316 11228 22372
rect 11284 22316 11294 22372
rect 11554 22316 11564 22372
rect 11620 22316 11900 22372
rect 11956 22316 12348 22372
rect 12404 22316 12414 22372
rect 12786 22316 12796 22372
rect 12852 22316 14252 22372
rect 14308 22316 15596 22372
rect 15652 22316 15662 22372
rect 20850 22316 20860 22372
rect 20916 22316 21644 22372
rect 21700 22316 23884 22372
rect 23940 22316 23950 22372
rect 27906 22316 27916 22372
rect 27972 22316 29484 22372
rect 29540 22316 29550 22372
rect 33730 22316 33740 22372
rect 33796 22316 34860 22372
rect 34916 22316 35420 22372
rect 35476 22316 35486 22372
rect 40114 22316 40124 22372
rect 40180 22316 43988 22372
rect 44044 22316 44054 22372
rect 2370 22204 2380 22260
rect 2436 22204 3836 22260
rect 3892 22204 4676 22260
rect 4732 22204 5292 22260
rect 5348 22204 5358 22260
rect 10220 22204 12068 22260
rect 12124 22204 12134 22260
rect 26562 22204 26572 22260
rect 26628 22204 27636 22260
rect 27692 22204 27702 22260
rect 34290 22204 34300 22260
rect 34356 22204 37548 22260
rect 37604 22204 37614 22260
rect 43362 22204 43372 22260
rect 43428 22204 44156 22260
rect 44212 22204 44828 22260
rect 44884 22204 44894 22260
rect 10220 22148 10276 22204
rect 4162 22092 4172 22148
rect 4228 22092 4956 22148
rect 5012 22092 5022 22148
rect 10210 22092 10220 22148
rect 10276 22092 10286 22148
rect 12226 22092 12236 22148
rect 12292 22092 12572 22148
rect 12628 22092 14028 22148
rect 14084 22092 16044 22148
rect 16100 22092 20524 22148
rect 20580 22092 20590 22148
rect 28578 22092 28588 22148
rect 28644 22092 30156 22148
rect 30212 22092 30222 22148
rect 30538 22092 30548 22148
rect 30604 22092 39228 22148
rect 39284 22092 39294 22148
rect 12338 21980 12348 22036
rect 12404 21980 14364 22036
rect 14420 21980 14430 22036
rect 21858 21980 21868 22036
rect 21924 21980 36988 22036
rect 37044 21980 37054 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 13794 21868 13804 21924
rect 13860 21868 15148 21924
rect 15204 21868 17276 21924
rect 17332 21868 17342 21924
rect 23202 21868 23212 21924
rect 23268 21868 23660 21924
rect 23716 21868 25116 21924
rect 25172 21868 25182 21924
rect 25340 21868 25452 21924
rect 25508 21868 25518 21924
rect 30258 21868 30268 21924
rect 30324 21868 30604 21924
rect 30660 21868 30670 21924
rect 34962 21868 34972 21924
rect 35028 21868 37212 21924
rect 37268 21868 37278 21924
rect 25340 21812 25396 21868
rect 3042 21756 3052 21812
rect 3108 21756 3118 21812
rect 11386 21756 11396 21812
rect 11452 21756 12908 21812
rect 12964 21756 12974 21812
rect 17602 21756 17612 21812
rect 17668 21756 18844 21812
rect 18900 21756 18910 21812
rect 22474 21756 22484 21812
rect 22540 21756 22652 21812
rect 22708 21756 23996 21812
rect 24052 21756 25396 21812
rect 27458 21756 27468 21812
rect 27524 21756 27534 21812
rect 28130 21756 28140 21812
rect 28196 21756 29708 21812
rect 29764 21756 29774 21812
rect 29978 21756 29988 21812
rect 30044 21756 30940 21812
rect 30996 21756 31006 21812
rect 33394 21756 33404 21812
rect 33460 21756 33740 21812
rect 33796 21756 34412 21812
rect 34468 21756 34478 21812
rect 3052 21252 3108 21756
rect 27468 21700 27524 21756
rect 14578 21644 14588 21700
rect 14644 21644 16268 21700
rect 16324 21644 17500 21700
rect 17556 21644 17566 21700
rect 27468 21644 31276 21700
rect 31332 21644 31342 21700
rect 37986 21644 37996 21700
rect 38052 21644 38220 21700
rect 38276 21644 38286 21700
rect 42242 21644 42252 21700
rect 42308 21644 44604 21700
rect 44660 21644 44670 21700
rect 45490 21644 45500 21700
rect 45556 21644 46060 21700
rect 46116 21644 48860 21700
rect 48916 21644 48926 21700
rect 21746 21532 21756 21588
rect 21812 21532 22876 21588
rect 22932 21532 22942 21588
rect 25666 21532 25676 21588
rect 25732 21532 26964 21588
rect 27020 21532 30716 21588
rect 30772 21532 30782 21588
rect 31602 21532 31612 21588
rect 31668 21532 32956 21588
rect 33012 21532 33022 21588
rect 33842 21532 33852 21588
rect 33908 21532 36092 21588
rect 36148 21532 36428 21588
rect 36484 21532 36494 21588
rect 37426 21532 37436 21588
rect 37492 21532 38892 21588
rect 38948 21532 38958 21588
rect 41122 21532 41132 21588
rect 41188 21532 44884 21588
rect 44940 21532 44950 21588
rect 46162 21532 46172 21588
rect 46228 21532 47852 21588
rect 47908 21532 47918 21588
rect 4274 21420 4284 21476
rect 4340 21420 4844 21476
rect 4900 21420 5180 21476
rect 5236 21420 5246 21476
rect 11834 21420 11844 21476
rect 11900 21420 12348 21476
rect 12404 21420 12414 21476
rect 17042 21420 17052 21476
rect 17108 21420 23100 21476
rect 23156 21420 23166 21476
rect 31266 21420 31276 21476
rect 31332 21420 32396 21476
rect 32452 21420 32462 21476
rect 37538 21420 37548 21476
rect 37604 21420 37884 21476
rect 37940 21420 37950 21476
rect 38210 21420 38220 21476
rect 38276 21420 40460 21476
rect 40516 21420 40526 21476
rect 41290 21420 41300 21476
rect 41356 21420 42140 21476
rect 42196 21420 42206 21476
rect 42690 21420 42700 21476
rect 42756 21420 43820 21476
rect 43876 21420 47348 21476
rect 47404 21420 47414 21476
rect 47730 21420 47740 21476
rect 47796 21420 48524 21476
rect 48580 21420 48590 21476
rect 18610 21308 18620 21364
rect 18676 21308 19236 21364
rect 3052 21196 3276 21252
rect 3332 21196 3342 21252
rect 18498 21196 18508 21252
rect 18564 21196 18574 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 5618 21084 5628 21140
rect 5684 21084 7084 21140
rect 7140 21084 7150 21140
rect 3042 20972 3052 21028
rect 3108 20972 4284 21028
rect 4340 20972 4350 21028
rect 6458 20972 6468 21028
rect 6524 20972 6972 21028
rect 7028 20972 7700 21028
rect 7756 20972 7766 21028
rect 2594 20860 2604 20916
rect 2660 20860 3724 20916
rect 3780 20860 3790 20916
rect 12562 20860 12572 20916
rect 12628 20860 14028 20916
rect 14084 20860 17444 20916
rect 17500 20860 17510 20916
rect 18508 20804 18564 21196
rect 19180 21028 19236 21308
rect 29484 21308 29820 21364
rect 29876 21308 30492 21364
rect 30548 21308 31388 21364
rect 31444 21308 31454 21364
rect 34300 21308 35308 21364
rect 35364 21308 35374 21364
rect 35858 21308 35868 21364
rect 35924 21308 36092 21364
rect 36148 21308 36158 21364
rect 38770 21308 38780 21364
rect 38836 21308 40012 21364
rect 40068 21308 40078 21364
rect 41738 21308 41748 21364
rect 41804 21308 42364 21364
rect 42420 21308 42430 21364
rect 45266 21308 45276 21364
rect 45332 21308 48636 21364
rect 48692 21308 48860 21364
rect 48916 21308 48926 21364
rect 29484 21252 29540 21308
rect 34300 21252 34356 21308
rect 20178 21196 20188 21252
rect 20244 21196 20356 21252
rect 20412 21196 22428 21252
rect 22484 21196 22494 21252
rect 22642 21196 22652 21252
rect 22708 21196 22718 21252
rect 29474 21196 29484 21252
rect 29540 21196 29550 21252
rect 34290 21196 34300 21252
rect 34356 21196 34366 21252
rect 38882 21196 38892 21252
rect 38948 21196 39564 21252
rect 39620 21196 42588 21252
rect 42644 21196 42654 21252
rect 43978 21196 43988 21252
rect 44044 21196 45836 21252
rect 45892 21196 45902 21252
rect 22652 21140 22708 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 22082 21084 22092 21140
rect 22148 21084 22708 21140
rect 24770 21084 24780 21140
rect 24836 21084 32564 21140
rect 32620 21084 34188 21140
rect 34244 21084 34254 21140
rect 19180 20972 19272 21028
rect 19328 20972 20188 21028
rect 20244 20972 20254 21028
rect 24098 20972 24108 21028
rect 24164 20972 25228 21028
rect 25284 20972 25294 21028
rect 33618 20972 33628 21028
rect 33684 20972 34860 21028
rect 34916 20972 35532 21028
rect 35588 20972 35598 21028
rect 38612 20972 40908 21028
rect 40964 20972 40974 21028
rect 38612 20916 38668 20972
rect 23090 20860 23100 20916
rect 23156 20860 23772 20916
rect 23828 20860 25340 20916
rect 25396 20860 25406 20916
rect 30706 20860 30716 20916
rect 30772 20860 38668 20916
rect 24780 20804 24836 20860
rect 2370 20748 2380 20804
rect 2436 20748 3500 20804
rect 3556 20748 3566 20804
rect 7858 20748 7868 20804
rect 7924 20748 8092 20804
rect 8148 20748 8540 20804
rect 8596 20748 8606 20804
rect 9314 20748 9324 20804
rect 9380 20748 9660 20804
rect 9716 20748 12460 20804
rect 12516 20748 13356 20804
rect 13412 20748 14476 20804
rect 14532 20748 14924 20804
rect 14980 20748 14990 20804
rect 15922 20748 15932 20804
rect 15988 20748 18060 20804
rect 18116 20748 18126 20804
rect 18498 20748 18508 20804
rect 18564 20748 18574 20804
rect 23426 20748 23436 20804
rect 23492 20748 24444 20804
rect 24500 20748 24510 20804
rect 24770 20748 24780 20804
rect 24836 20748 24846 20804
rect 28690 20748 28700 20804
rect 28756 20748 29204 20804
rect 29260 20748 29270 20804
rect 32050 20748 32060 20804
rect 32116 20748 43148 20804
rect 43204 20748 43214 20804
rect 44258 20748 44268 20804
rect 44324 20748 45052 20804
rect 45108 20748 45118 20804
rect 47730 20748 47740 20804
rect 47796 20748 48972 20804
rect 49028 20748 49038 20804
rect 2706 20636 2716 20692
rect 2772 20636 4956 20692
rect 5012 20636 5022 20692
rect 22194 20636 22204 20692
rect 22260 20636 23548 20692
rect 23604 20636 23614 20692
rect 29586 20524 29596 20580
rect 29652 20524 35196 20580
rect 35252 20524 36372 20580
rect 36428 20524 36438 20580
rect 26852 20412 36988 20468
rect 37044 20412 38668 20468
rect 40898 20412 40908 20468
rect 40964 20412 41804 20468
rect 41860 20412 42700 20468
rect 42756 20412 42766 20468
rect 46834 20412 46844 20468
rect 46900 20412 49308 20468
rect 49364 20412 49374 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 26852 20356 26908 20412
rect 38108 20356 38164 20412
rect 38612 20356 38668 20412
rect 6626 20300 6636 20356
rect 6692 20300 7364 20356
rect 15318 20300 15328 20356
rect 15384 20300 16828 20356
rect 16884 20300 17948 20356
rect 18004 20300 18396 20356
rect 18452 20300 18462 20356
rect 22418 20300 22428 20356
rect 22484 20300 26908 20356
rect 29138 20300 29148 20356
rect 29204 20300 30044 20356
rect 30100 20300 33068 20356
rect 33124 20300 37548 20356
rect 37604 20300 37614 20356
rect 38098 20300 38108 20356
rect 38164 20300 38174 20356
rect 38612 20300 41356 20356
rect 41412 20300 41422 20356
rect 46610 20300 46620 20356
rect 46676 20300 48300 20356
rect 48356 20300 48366 20356
rect 7308 20244 7364 20300
rect 5898 20188 5908 20244
rect 5964 20188 6188 20244
rect 6244 20188 6254 20244
rect 6850 20188 6860 20244
rect 6916 20188 6926 20244
rect 7298 20188 7308 20244
rect 7364 20188 8820 20244
rect 8876 20188 8886 20244
rect 12562 20188 12572 20244
rect 12628 20188 14700 20244
rect 14756 20188 14766 20244
rect 30258 20188 30268 20244
rect 30324 20188 32060 20244
rect 32116 20188 32126 20244
rect 34346 20188 34356 20244
rect 34412 20188 36204 20244
rect 36260 20188 36270 20244
rect 41906 20188 41916 20244
rect 41972 20188 43652 20244
rect 46050 20188 46060 20244
rect 46116 20188 46956 20244
rect 47012 20188 47022 20244
rect 6860 20132 6916 20188
rect 43596 20132 43652 20188
rect 4946 20076 4956 20132
rect 5012 20076 6412 20132
rect 6468 20076 6916 20132
rect 12674 20076 12684 20132
rect 12740 20076 12750 20132
rect 13458 20076 13468 20132
rect 13524 20076 17612 20132
rect 17668 20076 19852 20132
rect 19908 20076 24052 20132
rect 24108 20076 24724 20132
rect 24882 20076 24892 20132
rect 24948 20076 27468 20132
rect 27524 20076 27534 20132
rect 28242 20076 28252 20132
rect 28308 20076 28812 20132
rect 28868 20076 28878 20132
rect 29474 20076 29484 20132
rect 29540 20076 33236 20132
rect 33292 20076 33302 20132
rect 33842 20076 33852 20132
rect 33908 20076 34748 20132
rect 34804 20076 34814 20132
rect 42354 20076 42364 20132
rect 42420 20076 42920 20132
rect 42976 20076 42986 20132
rect 43586 20076 43596 20132
rect 43652 20076 45332 20132
rect 45388 20076 45948 20132
rect 46004 20076 46014 20132
rect 3602 19964 3612 20020
rect 3668 19964 4732 20020
rect 4788 19964 4798 20020
rect 5394 19964 5404 20020
rect 5460 19964 5740 20020
rect 5796 19964 7756 20020
rect 7812 19964 7822 20020
rect 12684 19684 12740 20076
rect 24668 20020 24724 20076
rect 16706 19964 16716 20020
rect 16772 19964 16940 20020
rect 16996 19964 20412 20020
rect 20468 19964 20478 20020
rect 21018 19964 21028 20020
rect 21084 19964 21868 20020
rect 21924 19964 22876 20020
rect 22932 19964 22942 20020
rect 24668 19964 25228 20020
rect 25284 19964 25294 20020
rect 31042 19964 31052 20020
rect 31108 19964 31276 20020
rect 31332 19964 31342 20020
rect 31938 19964 31948 20020
rect 32004 19964 35140 20020
rect 35196 19964 35206 20020
rect 37650 19964 37660 20020
rect 37716 19964 38556 20020
rect 38612 19964 39004 20020
rect 39060 19964 39070 20020
rect 43698 19964 43708 20020
rect 43764 19964 44322 20020
rect 44378 19964 44388 20020
rect 47058 19964 47068 20020
rect 47124 19964 48636 20020
rect 48692 19964 48702 20020
rect 17602 19852 17612 19908
rect 17668 19852 18732 19908
rect 18788 19852 18798 19908
rect 18946 19852 18956 19908
rect 19012 19852 20188 19908
rect 20244 19852 21476 19908
rect 21532 19852 22540 19908
rect 22596 19852 22606 19908
rect 23482 19852 23492 19908
rect 23548 19852 29260 19908
rect 29316 19852 29326 19908
rect 30762 19852 30772 19908
rect 30828 19852 31612 19908
rect 31668 19852 31678 19908
rect 33954 19852 33964 19908
rect 34020 19852 35588 19908
rect 37874 19852 37884 19908
rect 37940 19852 38444 19908
rect 38500 19852 38510 19908
rect 39890 19852 39900 19908
rect 39956 19852 41356 19908
rect 41412 19852 42028 19908
rect 42084 19852 42094 19908
rect 42634 19852 42644 19908
rect 42700 19852 44996 19908
rect 45052 19852 45062 19908
rect 13010 19740 13020 19796
rect 13076 19740 14194 19796
rect 14250 19740 14260 19796
rect 19618 19740 19628 19796
rect 19684 19740 20076 19796
rect 20132 19740 20142 19796
rect 24434 19740 24444 19796
rect 24500 19740 25564 19796
rect 25620 19740 25630 19796
rect 29698 19740 29708 19796
rect 29764 19740 30380 19796
rect 30436 19740 34860 19796
rect 34916 19740 34926 19796
rect 30828 19684 30884 19740
rect 35532 19684 35588 19852
rect 38658 19740 38668 19796
rect 38724 19740 40124 19796
rect 40180 19740 40190 19796
rect 43474 19740 43484 19796
rect 43540 19740 46956 19796
rect 47012 19740 47022 19796
rect 12684 19628 16716 19684
rect 16772 19628 16782 19684
rect 28914 19628 28924 19684
rect 28980 19628 30156 19684
rect 30212 19628 30222 19684
rect 30818 19628 30828 19684
rect 30884 19628 30894 19684
rect 31378 19628 31388 19684
rect 31444 19628 32956 19684
rect 33012 19628 33022 19684
rect 35532 19628 44716 19684
rect 44772 19628 44782 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 12450 19516 12460 19572
rect 12516 19516 13916 19572
rect 13972 19516 13982 19572
rect 27570 19516 27580 19572
rect 27636 19516 28364 19572
rect 28420 19516 34636 19572
rect 34692 19516 34702 19572
rect 38882 19516 38892 19572
rect 38948 19516 39788 19572
rect 39844 19516 40684 19572
rect 40740 19516 40750 19572
rect 42910 19516 42920 19572
rect 42976 19516 42986 19572
rect 42924 19460 42980 19516
rect 2370 19404 2380 19460
rect 2436 19404 5292 19460
rect 5348 19404 5358 19460
rect 27346 19404 27356 19460
rect 27412 19404 28140 19460
rect 28196 19404 29596 19460
rect 29652 19404 29662 19460
rect 30146 19404 30156 19460
rect 30212 19404 32452 19460
rect 32508 19404 37100 19460
rect 37156 19404 37166 19460
rect 39890 19404 39900 19460
rect 39956 19404 40348 19460
rect 40404 19404 40414 19460
rect 42924 19404 43484 19460
rect 43540 19404 45444 19460
rect 45500 19404 49532 19460
rect 49588 19404 49598 19460
rect 4722 19292 4732 19348
rect 4788 19292 5628 19348
rect 5684 19292 5694 19348
rect 14578 19292 14588 19348
rect 14644 19292 16436 19348
rect 16492 19292 16502 19348
rect 28578 19292 28588 19348
rect 28644 19292 29484 19348
rect 29540 19292 29550 19348
rect 35746 19292 35756 19348
rect 35812 19292 36652 19348
rect 36708 19292 36718 19348
rect 48626 19292 48636 19348
rect 48692 19292 49084 19348
rect 49140 19292 49150 19348
rect 11890 19180 11900 19236
rect 11956 19180 13356 19236
rect 13412 19180 13422 19236
rect 15082 19180 15092 19236
rect 15148 19180 16268 19236
rect 16324 19180 16334 19236
rect 20850 19180 20860 19236
rect 20916 19180 21196 19236
rect 21252 19180 24892 19236
rect 24948 19180 24958 19236
rect 28242 19180 28252 19236
rect 28308 19180 29260 19236
rect 29316 19180 29326 19236
rect 31154 19180 31164 19236
rect 31220 19180 31388 19236
rect 31444 19180 31454 19236
rect 36530 19180 36540 19236
rect 36596 19180 37100 19236
rect 37156 19180 37166 19236
rect 46386 19180 46396 19236
rect 46452 19180 47292 19236
rect 47348 19180 49308 19236
rect 49364 19180 49374 19236
rect 31164 19124 31220 19180
rect 50200 19124 51000 19152
rect 13738 19068 13748 19124
rect 13804 19068 16604 19124
rect 16660 19068 16670 19124
rect 23202 19068 23212 19124
rect 23268 19068 23884 19124
rect 23940 19068 23950 19124
rect 28578 19068 28588 19124
rect 28644 19068 31220 19124
rect 49410 19068 49420 19124
rect 49476 19068 51000 19124
rect 50200 19040 51000 19068
rect 13514 18956 13524 19012
rect 13580 18956 15596 19012
rect 15652 18956 15662 19012
rect 3826 18844 3836 18900
rect 3892 18844 5068 18900
rect 5124 18844 5134 18900
rect 13906 18844 13916 18900
rect 13972 18844 16492 18900
rect 16548 18844 16558 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 20906 18732 20916 18788
rect 20972 18732 21980 18788
rect 22036 18732 22046 18788
rect 28018 18732 28028 18788
rect 28084 18732 29988 18788
rect 30044 18732 30054 18788
rect 35970 18732 35980 18788
rect 36036 18732 36652 18788
rect 36708 18732 36718 18788
rect 15810 18620 15820 18676
rect 15876 18620 15886 18676
rect 33898 18620 33908 18676
rect 33964 18620 35532 18676
rect 35588 18620 35598 18676
rect 35858 18620 35868 18676
rect 35924 18620 36484 18676
rect 36978 18620 36988 18676
rect 37044 18620 39900 18676
rect 39956 18620 39966 18676
rect 15820 18564 15876 18620
rect 3042 18508 3052 18564
rect 3108 18508 4284 18564
rect 4340 18508 4350 18564
rect 12796 18508 13916 18564
rect 13972 18508 13982 18564
rect 15820 18508 17500 18564
rect 17556 18508 20524 18564
rect 20580 18508 20590 18564
rect 22262 18508 22272 18564
rect 22328 18508 23212 18564
rect 23268 18508 23278 18564
rect 26338 18508 26348 18564
rect 26404 18508 27916 18564
rect 27972 18508 27982 18564
rect 1586 18396 1596 18452
rect 1652 18396 2044 18452
rect 2100 18396 4060 18452
rect 4116 18396 6524 18452
rect 6580 18396 6590 18452
rect 3490 18284 3500 18340
rect 3556 18284 4508 18340
rect 4564 18284 6076 18340
rect 6132 18284 6142 18340
rect 4386 18172 4396 18228
rect 4452 18172 5460 18228
rect 5516 18172 5526 18228
rect 5730 18172 5740 18228
rect 5796 18172 7084 18228
rect 7140 18172 7644 18228
rect 7700 18172 7710 18228
rect 6300 18116 6356 18172
rect 12796 18116 12852 18508
rect 36428 18452 36484 18620
rect 36866 18508 36876 18564
rect 36932 18508 37100 18564
rect 37156 18508 37660 18564
rect 37716 18508 38332 18564
rect 38388 18508 38398 18564
rect 13346 18396 13356 18452
rect 13412 18396 15036 18452
rect 15092 18396 15102 18452
rect 18946 18396 18956 18452
rect 19012 18396 20748 18452
rect 20804 18396 21868 18452
rect 21924 18396 21934 18452
rect 23426 18396 23436 18452
rect 23492 18396 24220 18452
rect 24276 18396 24286 18452
rect 27122 18396 27132 18452
rect 27188 18396 31948 18452
rect 32004 18396 32014 18452
rect 32834 18396 32844 18452
rect 32900 18396 33628 18452
rect 33684 18396 34524 18452
rect 34580 18396 34590 18452
rect 36418 18396 36428 18452
rect 36484 18396 36494 18452
rect 38770 18396 38780 18452
rect 38836 18396 39116 18452
rect 39172 18396 39182 18452
rect 40226 18396 40236 18452
rect 40292 18396 41244 18452
rect 41300 18396 41804 18452
rect 41860 18396 41870 18452
rect 46442 18396 46452 18452
rect 46508 18396 47516 18452
rect 47572 18396 47582 18452
rect 39116 18340 39172 18396
rect 18386 18284 18396 18340
rect 18452 18284 21532 18340
rect 21588 18284 22540 18340
rect 22596 18284 22606 18340
rect 24546 18284 24556 18340
rect 24612 18284 24892 18340
rect 24948 18284 27356 18340
rect 27412 18284 27422 18340
rect 27682 18284 27692 18340
rect 27748 18284 28924 18340
rect 28980 18284 28990 18340
rect 39116 18284 42364 18340
rect 42420 18284 42430 18340
rect 41804 18228 41860 18284
rect 41794 18172 41804 18228
rect 41860 18172 41870 18228
rect 42578 18172 42588 18228
rect 42644 18172 45612 18228
rect 45668 18172 45678 18228
rect 6290 18060 6300 18116
rect 6356 18060 6366 18116
rect 12786 18060 12796 18116
rect 12852 18060 12862 18116
rect 15530 18060 15540 18116
rect 15596 18060 15932 18116
rect 15988 18060 16716 18116
rect 16772 18060 17276 18116
rect 17332 18060 17342 18116
rect 37986 18060 37996 18116
rect 38052 18060 39564 18116
rect 39620 18060 41356 18116
rect 41412 18060 41422 18116
rect 43810 18060 43820 18116
rect 43876 18060 44044 18116
rect 44100 18060 44110 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 4834 17948 4844 18004
rect 4900 17948 6636 18004
rect 6692 17948 6702 18004
rect 11909 17948 11919 18004
rect 11975 17948 13580 18004
rect 13636 17948 15148 18004
rect 39890 17948 39900 18004
rect 39956 17948 43708 18004
rect 43764 17948 43774 18004
rect 15092 17892 15148 17948
rect 5170 17836 5180 17892
rect 5236 17836 5516 17892
rect 5572 17836 6972 17892
rect 7028 17836 7038 17892
rect 15092 17836 16156 17892
rect 16212 17836 16222 17892
rect 18050 17836 18060 17892
rect 18116 17836 18396 17892
rect 18452 17836 19348 17892
rect 19404 17836 24052 17892
rect 24108 17836 24118 17892
rect 32274 17836 32284 17892
rect 32340 17836 35028 17892
rect 35084 17836 35094 17892
rect 40394 17836 40404 17892
rect 40460 17836 48972 17892
rect 49028 17836 49038 17892
rect 5954 17724 5964 17780
rect 6020 17724 6524 17780
rect 6580 17724 6590 17780
rect 8306 17724 8316 17780
rect 8372 17724 8988 17780
rect 9044 17724 9054 17780
rect 11554 17724 11564 17780
rect 11620 17724 12236 17780
rect 12292 17724 12302 17780
rect 14802 17724 14812 17780
rect 14868 17724 15820 17780
rect 15876 17724 15886 17780
rect 21410 17724 21420 17780
rect 21476 17724 25228 17780
rect 25284 17724 26348 17780
rect 26404 17724 26414 17780
rect 33730 17724 33740 17780
rect 33796 17724 35420 17780
rect 35476 17724 35486 17780
rect 4274 17612 4284 17668
rect 4340 17612 5740 17668
rect 5796 17612 5806 17668
rect 8866 17612 8876 17668
rect 8932 17612 9548 17668
rect 9604 17612 9940 17668
rect 9996 17612 10006 17668
rect 11442 17612 11452 17668
rect 11508 17612 13860 17668
rect 13916 17612 16716 17668
rect 16772 17612 16782 17668
rect 17938 17612 17948 17668
rect 18004 17612 18844 17668
rect 18900 17612 18910 17668
rect 23090 17612 23100 17668
rect 23156 17612 23772 17668
rect 23828 17612 23838 17668
rect 24322 17612 24332 17668
rect 24388 17612 25452 17668
rect 25508 17612 25518 17668
rect 26786 17612 26796 17668
rect 26852 17612 27020 17668
rect 27076 17612 27086 17668
rect 31042 17612 31052 17668
rect 31108 17612 31948 17668
rect 32004 17612 33404 17668
rect 33460 17612 33470 17668
rect 34514 17612 34524 17668
rect 34580 17612 35308 17668
rect 35364 17612 35374 17668
rect 43810 17612 43820 17668
rect 43876 17612 45276 17668
rect 45332 17612 46620 17668
rect 46676 17612 46686 17668
rect 5394 17500 5404 17556
rect 5460 17500 5908 17556
rect 5964 17500 5974 17556
rect 12562 17500 12572 17556
rect 12628 17500 14812 17556
rect 14868 17500 16996 17556
rect 17052 17500 17062 17556
rect 20850 17500 20860 17556
rect 20916 17500 21980 17556
rect 22036 17500 22046 17556
rect 23650 17500 23660 17556
rect 23716 17500 24780 17556
rect 24836 17500 28588 17556
rect 28644 17500 28654 17556
rect 5170 17388 5180 17444
rect 5236 17388 9100 17444
rect 9156 17388 9166 17444
rect 11890 17388 11900 17444
rect 11956 17388 16156 17444
rect 16212 17388 16604 17444
rect 16660 17388 17612 17444
rect 17668 17388 17678 17444
rect 25330 17388 25340 17444
rect 25396 17388 25788 17444
rect 25844 17388 25854 17444
rect 26012 17388 27244 17444
rect 27300 17388 27310 17444
rect 34178 17388 34188 17444
rect 34244 17388 35980 17444
rect 36036 17388 36046 17444
rect 37874 17388 37884 17444
rect 37940 17388 41692 17444
rect 41748 17388 45948 17444
rect 46004 17388 46014 17444
rect 26012 17332 26068 17388
rect 6962 17276 6972 17332
rect 7028 17276 8596 17332
rect 23650 17276 23660 17332
rect 23716 17276 24612 17332
rect 24668 17276 26068 17332
rect 26620 17276 26630 17332
rect 26686 17276 27542 17332
rect 27598 17276 34412 17332
rect 34468 17276 34478 17332
rect 8540 17108 8596 17276
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 25554 17164 25564 17220
rect 25620 17164 27132 17220
rect 27188 17164 27692 17220
rect 27748 17164 27758 17220
rect 29036 17164 31164 17220
rect 31220 17164 31230 17220
rect 3938 17052 3948 17108
rect 4004 17052 4284 17108
rect 4340 17052 5852 17108
rect 5908 17052 6636 17108
rect 6692 17052 6702 17108
rect 8530 17052 8540 17108
rect 8596 17052 9324 17108
rect 9380 17052 9390 17108
rect 11218 17052 11228 17108
rect 11284 17052 12796 17108
rect 12852 17052 12862 17108
rect 21746 17052 21756 17108
rect 21812 17052 23100 17108
rect 23156 17052 23548 17108
rect 23604 17052 23614 17108
rect 24098 17052 24108 17108
rect 24164 17052 27020 17108
rect 27076 17052 27356 17108
rect 27412 17052 27422 17108
rect 24108 16996 24164 17052
rect 29036 16996 29092 17164
rect 30146 17052 30156 17108
rect 30212 17052 31612 17108
rect 31668 17052 31678 17108
rect 38994 17052 39004 17108
rect 39060 17052 39070 17108
rect 39004 16996 39060 17052
rect 5954 16940 5964 16996
rect 6020 16940 7420 16996
rect 7476 16940 7486 16996
rect 8698 16940 8708 16996
rect 8764 16940 9436 16996
rect 9492 16940 9502 16996
rect 15026 16940 15036 16996
rect 15092 16940 16380 16996
rect 16436 16940 16446 16996
rect 23426 16940 23436 16996
rect 23492 16940 24164 16996
rect 26796 16940 29092 16996
rect 30370 16940 30380 16996
rect 30436 16940 31276 16996
rect 31332 16940 31948 16996
rect 32004 16940 33236 16996
rect 33292 16940 33302 16996
rect 39004 16940 41076 16996
rect 41132 16940 41142 16996
rect 23436 16884 23492 16940
rect 26796 16884 26852 16940
rect 40124 16884 40180 16940
rect 4162 16828 4172 16884
rect 4228 16828 5068 16884
rect 5124 16828 5134 16884
rect 6122 16828 6132 16884
rect 6188 16828 10052 16884
rect 13682 16828 13692 16884
rect 13748 16828 14028 16884
rect 14084 16828 16044 16884
rect 16100 16828 16110 16884
rect 17938 16828 17948 16884
rect 18004 16828 19516 16884
rect 19572 16828 19582 16884
rect 22082 16828 22092 16884
rect 22148 16828 23492 16884
rect 26786 16828 26796 16884
rect 26852 16828 26862 16884
rect 26954 16828 26964 16884
rect 27020 16828 27916 16884
rect 27972 16828 27982 16884
rect 28914 16828 28924 16884
rect 28980 16828 29260 16884
rect 29316 16828 30044 16884
rect 30100 16828 30110 16884
rect 34402 16828 34412 16884
rect 34468 16828 37548 16884
rect 37604 16828 37614 16884
rect 40114 16828 40124 16884
rect 40180 16828 40190 16884
rect 41234 16828 41244 16884
rect 41300 16828 42476 16884
rect 42532 16828 42700 16884
rect 42756 16828 43484 16884
rect 43540 16828 43550 16884
rect 43708 16828 44268 16884
rect 44324 16828 44334 16884
rect 44538 16828 44548 16884
rect 44604 16828 45276 16884
rect 45332 16828 47068 16884
rect 47124 16828 47134 16884
rect 9996 16772 10052 16828
rect 43708 16772 43764 16828
rect 6738 16716 6748 16772
rect 6804 16716 8204 16772
rect 8260 16716 8270 16772
rect 9996 16716 11004 16772
rect 11060 16716 11070 16772
rect 22754 16716 22764 16772
rect 22820 16716 23324 16772
rect 23380 16716 23390 16772
rect 35746 16716 35756 16772
rect 35812 16716 36764 16772
rect 36820 16716 38556 16772
rect 38612 16716 39340 16772
rect 39396 16716 39406 16772
rect 40002 16716 40012 16772
rect 40068 16716 40236 16772
rect 40292 16716 40302 16772
rect 42252 16716 43764 16772
rect 7084 16660 7140 16716
rect 42252 16660 42308 16716
rect 7074 16604 7084 16660
rect 7140 16604 7150 16660
rect 9762 16604 9772 16660
rect 9828 16604 10444 16660
rect 10500 16604 10510 16660
rect 16650 16604 16660 16660
rect 16716 16604 18172 16660
rect 18228 16604 18844 16660
rect 18900 16604 18910 16660
rect 41804 16604 42084 16660
rect 42140 16604 42308 16660
rect 41804 16548 41860 16604
rect 41794 16492 41804 16548
rect 41860 16492 41870 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 18386 16380 18396 16436
rect 18452 16380 19068 16436
rect 19124 16380 19134 16436
rect 43250 16380 43260 16436
rect 43316 16380 44044 16436
rect 44100 16380 44940 16436
rect 44996 16380 45006 16436
rect 3378 16268 3388 16324
rect 3444 16268 4732 16324
rect 4788 16268 5404 16324
rect 5460 16268 5470 16324
rect 10882 16268 10892 16324
rect 10948 16268 11676 16324
rect 11732 16268 11742 16324
rect 24210 16268 24220 16324
rect 24276 16268 24286 16324
rect 30774 16268 30784 16324
rect 30840 16268 36204 16324
rect 36260 16268 36270 16324
rect 24220 16212 24276 16268
rect 19506 16156 19516 16212
rect 19572 16156 20132 16212
rect 20188 16156 20198 16212
rect 24220 16156 25508 16212
rect 25666 16156 25676 16212
rect 25732 16156 27916 16212
rect 27972 16156 27982 16212
rect 33226 16156 33236 16212
rect 33292 16156 36484 16212
rect 36540 16156 36988 16212
rect 37044 16156 37054 16212
rect 43698 16156 43708 16212
rect 43764 16156 44212 16212
rect 44268 16156 45724 16212
rect 45780 16156 45790 16212
rect 25452 16100 25508 16156
rect 2818 16044 2828 16100
rect 2884 16044 5292 16100
rect 5348 16044 5358 16100
rect 13458 16044 13468 16100
rect 13524 16044 13916 16100
rect 13972 16044 13982 16100
rect 17154 16044 17164 16100
rect 17220 16044 19964 16100
rect 20020 16044 20030 16100
rect 22194 16044 22204 16100
rect 22260 16044 22988 16100
rect 23044 16044 23054 16100
rect 23314 16044 23324 16100
rect 23380 16044 24220 16100
rect 24276 16044 24286 16100
rect 25452 16044 25564 16100
rect 25620 16044 25630 16100
rect 27794 16044 27804 16100
rect 27860 16044 28252 16100
rect 28308 16044 28700 16100
rect 28756 16044 30940 16100
rect 30996 16044 31006 16100
rect 37650 16044 37660 16100
rect 37716 16044 40236 16100
rect 40292 16044 40302 16100
rect 3154 15932 3164 15988
rect 3220 15932 4284 15988
rect 4340 15932 4620 15988
rect 4676 15932 6300 15988
rect 6356 15932 6366 15988
rect 24714 15932 24724 15988
rect 24780 15932 25116 15988
rect 25172 15932 25182 15988
rect 10994 15820 11004 15876
rect 11060 15820 13636 15876
rect 13692 15820 15932 15876
rect 15988 15820 15998 15876
rect 47170 15820 47180 15876
rect 47236 15820 48076 15876
rect 48132 15820 48142 15876
rect 3490 15708 3500 15764
rect 3556 15708 4620 15764
rect 4676 15708 4686 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 23874 15596 23884 15652
rect 23940 15596 24668 15652
rect 24724 15596 24734 15652
rect 29474 15596 29484 15652
rect 29540 15596 30604 15652
rect 30660 15596 31724 15652
rect 31780 15596 33124 15652
rect 33180 15596 33190 15652
rect 42354 15596 42364 15652
rect 42420 15596 43036 15652
rect 43092 15596 43102 15652
rect 20010 15484 20020 15540
rect 20076 15484 20300 15540
rect 20356 15484 20366 15540
rect 20850 15484 20860 15540
rect 20916 15484 22428 15540
rect 22484 15484 22494 15540
rect 22978 15484 22988 15540
rect 23044 15484 24500 15540
rect 24556 15484 24566 15540
rect 29250 15484 29260 15540
rect 29316 15484 30492 15540
rect 30548 15484 30558 15540
rect 39106 15484 39116 15540
rect 39172 15484 39900 15540
rect 39956 15484 39966 15540
rect 42466 15484 42476 15540
rect 42532 15484 42924 15540
rect 42980 15484 43372 15540
rect 43428 15484 43820 15540
rect 43876 15484 44716 15540
rect 44772 15484 47628 15540
rect 47684 15484 47694 15540
rect 22754 15372 22764 15428
rect 22820 15372 24332 15428
rect 24388 15372 24398 15428
rect 41794 15372 41804 15428
rect 41860 15372 43148 15428
rect 43204 15372 43214 15428
rect 2818 15260 2828 15316
rect 2884 15260 4620 15316
rect 4676 15260 4686 15316
rect 5170 15260 5180 15316
rect 5236 15260 6972 15316
rect 7028 15260 8036 15316
rect 8092 15260 8102 15316
rect 9762 15260 9772 15316
rect 9828 15260 11004 15316
rect 11060 15260 11070 15316
rect 19208 15260 19218 15316
rect 19274 15260 20524 15316
rect 20580 15260 21980 15316
rect 22036 15260 22046 15316
rect 22418 15260 22428 15316
rect 22484 15260 23212 15316
rect 23268 15260 23278 15316
rect 23874 15260 23884 15316
rect 23940 15260 26012 15316
rect 26068 15260 26236 15316
rect 26292 15260 26302 15316
rect 31938 15260 31948 15316
rect 32004 15260 33628 15316
rect 33684 15260 33694 15316
rect 34906 15260 34916 15316
rect 34972 15260 35756 15316
rect 35812 15260 36540 15316
rect 36596 15260 36606 15316
rect 42242 15260 42252 15316
rect 42308 15260 42700 15316
rect 42756 15260 42766 15316
rect 43474 15260 43484 15316
rect 43540 15260 46396 15316
rect 46452 15260 47348 15316
rect 47404 15260 47414 15316
rect 6402 15148 6412 15204
rect 6468 15148 6860 15204
rect 6916 15148 6926 15204
rect 14578 15148 14588 15204
rect 14644 15148 18060 15204
rect 18116 15148 18126 15204
rect 18610 15148 18620 15204
rect 18676 15148 19516 15204
rect 19572 15148 19582 15204
rect 23650 15148 23660 15204
rect 23716 15148 24892 15204
rect 24948 15148 24958 15204
rect 33730 15148 33740 15204
rect 33796 15148 34076 15204
rect 34132 15148 35084 15204
rect 35140 15148 35150 15204
rect 41626 15148 41636 15204
rect 41692 15148 42308 15204
rect 19292 15092 19348 15148
rect 9986 15036 9996 15092
rect 10052 15036 11228 15092
rect 11284 15036 11900 15092
rect 11956 15036 13468 15092
rect 13524 15036 13534 15092
rect 19282 15036 19292 15092
rect 19348 15036 19358 15092
rect 25442 15036 25452 15092
rect 25508 15036 26796 15092
rect 26852 15036 26862 15092
rect 34300 15036 34468 15092
rect 34524 15036 35196 15092
rect 35252 15036 37100 15092
rect 37156 15036 37166 15092
rect 38322 15036 38332 15092
rect 38388 15036 39228 15092
rect 39284 15036 39294 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 5954 14812 5964 14868
rect 6020 14812 6524 14868
rect 6580 14812 7084 14868
rect 7140 14812 9548 14868
rect 9604 14812 9614 14868
rect 31826 14812 31836 14868
rect 31892 14812 32620 14868
rect 32676 14812 32686 14868
rect 6066 14700 6076 14756
rect 6132 14700 6412 14756
rect 6468 14700 7196 14756
rect 7252 14700 7262 14756
rect 29922 14700 29932 14756
rect 29988 14700 30884 14756
rect 30940 14700 30950 14756
rect 7410 14588 7420 14644
rect 7476 14588 8540 14644
rect 8596 14588 8606 14644
rect 9874 14588 9884 14644
rect 9940 14588 10444 14644
rect 10500 14588 10510 14644
rect 12114 14588 12124 14644
rect 12180 14588 13132 14644
rect 13188 14588 13198 14644
rect 18946 14588 18956 14644
rect 19012 14588 19404 14644
rect 19460 14588 20636 14644
rect 20692 14588 20702 14644
rect 31714 14588 31724 14644
rect 31780 14588 33404 14644
rect 33460 14588 33470 14644
rect 12124 14532 12180 14588
rect 34300 14532 34356 15036
rect 42252 14980 42308 15148
rect 43596 15148 46732 15204
rect 46788 15148 46798 15204
rect 43596 15092 43652 15148
rect 42802 15036 42812 15092
rect 42868 15036 43652 15092
rect 42252 14924 42364 14980
rect 42420 14924 43036 14980
rect 43092 14924 43484 14980
rect 43540 14924 43550 14980
rect 47730 14924 47740 14980
rect 47796 14924 48860 14980
rect 48916 14924 48926 14980
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 50200 14868 51000 14896
rect 47282 14812 47292 14868
rect 47348 14812 47628 14868
rect 47684 14812 47694 14868
rect 48066 14812 48076 14868
rect 48132 14812 48636 14868
rect 48692 14812 49084 14868
rect 49140 14812 49150 14868
rect 49308 14812 51000 14868
rect 49308 14756 49364 14812
rect 50200 14784 51000 14812
rect 35522 14700 35532 14756
rect 35588 14700 37324 14756
rect 37380 14700 37390 14756
rect 40114 14700 40124 14756
rect 40180 14700 49364 14756
rect 35634 14588 35644 14644
rect 35700 14588 36988 14644
rect 37044 14588 37054 14644
rect 6290 14476 6300 14532
rect 6356 14476 6972 14532
rect 7028 14476 7038 14532
rect 7746 14476 7756 14532
rect 7812 14476 9996 14532
rect 10052 14476 10062 14532
rect 10210 14476 10220 14532
rect 10276 14476 12180 14532
rect 12450 14476 12460 14532
rect 12516 14476 13020 14532
rect 13076 14476 13804 14532
rect 13860 14476 13870 14532
rect 16482 14476 16492 14532
rect 16548 14476 17276 14532
rect 17332 14476 17342 14532
rect 17490 14476 17500 14532
rect 17556 14476 18396 14532
rect 18452 14476 18462 14532
rect 19058 14476 19068 14532
rect 19124 14476 21084 14532
rect 21140 14476 21150 14532
rect 29362 14476 29372 14532
rect 29428 14476 30044 14532
rect 30100 14476 31052 14532
rect 31108 14476 31118 14532
rect 31378 14476 31388 14532
rect 31444 14476 32284 14532
rect 32340 14476 32350 14532
rect 34290 14476 34300 14532
rect 34356 14476 34366 14532
rect 35970 14476 35980 14532
rect 36036 14476 37660 14532
rect 37716 14476 37726 14532
rect 38658 14476 38668 14532
rect 38724 14476 39956 14532
rect 40012 14476 40022 14532
rect 5170 14364 5180 14420
rect 5236 14364 5516 14420
rect 5572 14364 6748 14420
rect 6804 14364 6814 14420
rect 16146 14364 16156 14420
rect 16212 14364 16716 14420
rect 16772 14364 16940 14420
rect 16996 14364 17006 14420
rect 18106 14364 18116 14420
rect 18172 14364 23212 14420
rect 23268 14364 23278 14420
rect 44818 14364 44828 14420
rect 44884 14364 45183 14420
rect 45239 14364 45249 14420
rect 20178 14252 20188 14308
rect 20244 14252 21644 14308
rect 21700 14252 22540 14308
rect 22596 14252 23436 14308
rect 23492 14252 23502 14308
rect 39218 14252 39228 14308
rect 39284 14252 39900 14308
rect 39956 14252 39966 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 21074 14028 21084 14084
rect 21140 14028 23100 14084
rect 23156 14028 23166 14084
rect 38210 14028 38220 14084
rect 38276 14028 41468 14084
rect 41524 14028 41972 14084
rect 42028 14028 42038 14084
rect 17602 13916 17612 13972
rect 17668 13916 19068 13972
rect 19124 13916 19134 13972
rect 40226 13916 40236 13972
rect 40292 13916 41692 13972
rect 41748 13916 41758 13972
rect 16818 13804 16828 13860
rect 16884 13804 17836 13860
rect 17892 13804 17902 13860
rect 19506 13804 19516 13860
rect 19572 13804 20524 13860
rect 20580 13804 20590 13860
rect 5282 13692 5292 13748
rect 5348 13692 6412 13748
rect 6468 13692 7868 13748
rect 7924 13692 7934 13748
rect 9090 13692 9100 13748
rect 9156 13692 9660 13748
rect 9716 13692 9726 13748
rect 17938 13692 17948 13748
rect 18004 13692 18956 13748
rect 19012 13692 19022 13748
rect 19730 13692 19740 13748
rect 19796 13692 20188 13748
rect 20244 13692 20254 13748
rect 21746 13692 21756 13748
rect 21812 13692 24668 13748
rect 24724 13692 25340 13748
rect 25396 13692 25406 13748
rect 32610 13692 32620 13748
rect 32676 13692 33740 13748
rect 33796 13692 33806 13748
rect 44818 13692 44828 13748
rect 44884 13692 47852 13748
rect 47908 13692 47918 13748
rect 48290 13692 48300 13748
rect 48356 13692 48860 13748
rect 48916 13692 48926 13748
rect 21756 13636 21812 13692
rect 20290 13580 20300 13636
rect 20356 13580 21812 13636
rect 47852 13636 47908 13692
rect 47852 13580 49140 13636
rect 49196 13580 49206 13636
rect 7802 13468 7812 13524
rect 7868 13468 10220 13524
rect 10276 13468 10286 13524
rect 16314 13468 16324 13524
rect 16380 13468 17836 13524
rect 17892 13468 18620 13524
rect 18676 13468 18686 13524
rect 19394 13468 19404 13524
rect 19460 13468 19628 13524
rect 19684 13468 22428 13524
rect 22484 13468 22988 13524
rect 23044 13468 23054 13524
rect 24098 13468 24108 13524
rect 24164 13468 25900 13524
rect 25956 13468 25966 13524
rect 29922 13468 29932 13524
rect 29988 13468 30492 13524
rect 30548 13468 31724 13524
rect 31780 13468 31790 13524
rect 31938 13468 31948 13524
rect 32004 13468 32284 13524
rect 32340 13468 32350 13524
rect 33506 13468 33516 13524
rect 33572 13468 38500 13524
rect 38556 13468 38566 13524
rect 42578 13468 42588 13524
rect 42644 13468 43596 13524
rect 43652 13468 46452 13524
rect 46508 13468 46518 13524
rect 18106 13356 18116 13412
rect 18172 13356 18788 13412
rect 18844 13356 18854 13412
rect 23202 13356 23212 13412
rect 23268 13356 25228 13412
rect 25284 13356 26572 13412
rect 26628 13356 26638 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 8978 13244 8988 13300
rect 9044 13244 9884 13300
rect 9940 13244 9950 13300
rect 24742 13244 24780 13300
rect 24836 13244 24846 13300
rect 25890 13244 25900 13300
rect 25956 13244 26796 13300
rect 26852 13244 27468 13300
rect 27524 13244 28364 13300
rect 28420 13244 29484 13300
rect 29540 13244 31052 13300
rect 31108 13244 31118 13300
rect 2538 13132 2548 13188
rect 2604 13132 4396 13188
rect 4452 13132 5180 13188
rect 5236 13132 6076 13188
rect 6132 13132 6142 13188
rect 22642 13132 22652 13188
rect 22708 13132 38668 13188
rect 14242 13020 14252 13076
rect 14308 13020 18060 13076
rect 18116 13020 18126 13076
rect 25442 13020 25452 13076
rect 25508 13020 26684 13076
rect 26740 13020 26750 13076
rect 29698 13020 29708 13076
rect 29764 13020 30380 13076
rect 30436 13020 30446 13076
rect 37762 13020 37772 13076
rect 37828 13020 38108 13076
rect 38164 13020 38174 13076
rect 38612 12964 38668 13132
rect 38882 13020 38892 13076
rect 38948 13020 39396 13076
rect 39452 13020 39900 13076
rect 39956 13020 41244 13076
rect 41300 13020 41310 13076
rect 43922 13020 43932 13076
rect 43988 13020 44940 13076
rect 44996 13020 45006 13076
rect 3714 12908 3724 12964
rect 3780 12908 5740 12964
rect 5796 12908 5806 12964
rect 6962 12908 6972 12964
rect 7028 12908 7532 12964
rect 7588 12908 7598 12964
rect 18610 12908 18620 12964
rect 18676 12908 19068 12964
rect 19124 12908 19964 12964
rect 20020 12908 20030 12964
rect 28242 12908 28252 12964
rect 28308 12908 29260 12964
rect 29316 12908 29326 12964
rect 29586 12908 29596 12964
rect 29652 12908 30716 12964
rect 30772 12908 31500 12964
rect 31556 12908 31566 12964
rect 38612 12908 39564 12964
rect 39620 12908 40516 12964
rect 40572 12908 40582 12964
rect 41906 12908 41916 12964
rect 41972 12908 45500 12964
rect 45556 12908 45566 12964
rect 6290 12796 6300 12852
rect 6356 12796 6636 12852
rect 6692 12796 8092 12852
rect 8148 12796 8876 12852
rect 8932 12796 8942 12852
rect 33058 12796 33068 12852
rect 33124 12796 34300 12852
rect 34356 12796 34366 12852
rect 41346 12796 41356 12852
rect 41412 12796 42756 12852
rect 42812 12796 43820 12852
rect 43876 12796 43886 12852
rect 44258 12796 44268 12852
rect 44324 12796 47180 12852
rect 47236 12796 47246 12852
rect 44268 12740 44324 12796
rect 24742 12684 24780 12740
rect 24836 12684 24846 12740
rect 28354 12684 28364 12740
rect 28420 12684 28812 12740
rect 28868 12684 29372 12740
rect 29428 12684 31948 12740
rect 32004 12684 32014 12740
rect 41010 12684 41020 12740
rect 41076 12684 41692 12740
rect 41748 12684 44324 12740
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 2706 12348 2716 12404
rect 2772 12348 6412 12404
rect 6468 12348 8428 12404
rect 8484 12348 8494 12404
rect 12450 12348 12460 12404
rect 12516 12348 13188 12404
rect 13244 12348 13254 12404
rect 21914 12348 21924 12404
rect 21980 12348 22876 12404
rect 22932 12348 22942 12404
rect 29138 12348 29148 12404
rect 29204 12348 32060 12404
rect 32116 12348 32564 12404
rect 32620 12348 32630 12404
rect 1586 12236 1596 12292
rect 1652 12236 5180 12292
rect 5236 12236 5246 12292
rect 7532 12236 10220 12292
rect 10276 12236 10286 12292
rect 14466 12236 14476 12292
rect 14532 12236 18060 12292
rect 18116 12236 18126 12292
rect 18218 12236 18228 12292
rect 18284 12236 19180 12292
rect 19236 12236 19246 12292
rect 27570 12236 27580 12292
rect 27636 12236 30044 12292
rect 30100 12236 30110 12292
rect 42578 12236 42588 12292
rect 42644 12236 43260 12292
rect 43316 12236 43326 12292
rect 7532 12180 7588 12236
rect 4274 12124 4284 12180
rect 4340 12124 5068 12180
rect 5124 12124 5628 12180
rect 5684 12124 5694 12180
rect 7522 12124 7532 12180
rect 7588 12124 7598 12180
rect 8306 12124 8316 12180
rect 8372 12124 8708 12180
rect 10434 12124 10444 12180
rect 10500 12124 11676 12180
rect 11732 12124 11742 12180
rect 17826 12124 17836 12180
rect 17892 12124 18508 12180
rect 18564 12124 18574 12180
rect 25778 12124 25788 12180
rect 25844 12124 26684 12180
rect 26740 12124 27244 12180
rect 27300 12124 27310 12180
rect 31042 12124 31052 12180
rect 31108 12124 32956 12180
rect 33012 12124 33022 12180
rect 41906 12124 41916 12180
rect 41972 12124 43932 12180
rect 43988 12124 43998 12180
rect 8652 12068 8708 12124
rect 4834 12012 4844 12068
rect 4900 12012 7924 12068
rect 7980 12012 8428 12068
rect 8484 12012 8494 12068
rect 8642 12012 8652 12068
rect 8708 12012 11004 12068
rect 11060 12012 11070 12068
rect 14802 12012 14812 12068
rect 14868 12012 19740 12068
rect 19796 12012 19806 12068
rect 32610 12012 32620 12068
rect 32676 12012 33740 12068
rect 33796 12012 33806 12068
rect 41402 12012 41412 12068
rect 41468 12012 42140 12068
rect 42196 12012 42206 12068
rect 46722 12012 46732 12068
rect 46788 12012 47404 12068
rect 47460 12012 47470 12068
rect 4946 11900 4956 11956
rect 5012 11900 7420 11956
rect 7476 11900 9716 11956
rect 9772 11900 9782 11956
rect 5170 11788 5180 11844
rect 5236 11788 8540 11844
rect 8596 11788 8606 11844
rect 8764 11788 9548 11844
rect 9604 11788 9614 11844
rect 18106 11788 18116 11844
rect 18172 11788 21420 11844
rect 21476 11788 21486 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 8764 11732 8820 11788
rect 26236 11732 26292 11956
rect 26348 11900 26358 11956
rect 34300 11900 35644 11956
rect 35700 11900 35710 11956
rect 36530 11900 36540 11956
rect 36596 11900 39508 11956
rect 39564 11900 39574 11956
rect 42802 11900 42812 11956
rect 42868 11900 43372 11956
rect 43428 11900 44996 11956
rect 34300 11844 34356 11900
rect 44940 11844 44996 11900
rect 34290 11788 34300 11844
rect 34356 11788 34366 11844
rect 42354 11788 42364 11844
rect 42420 11788 42476 11844
rect 42532 11788 42542 11844
rect 43810 11788 43820 11844
rect 43876 11788 44604 11844
rect 44660 11788 44670 11844
rect 44930 11788 44940 11844
rect 44996 11788 46284 11844
rect 46340 11788 48412 11844
rect 48468 11788 48478 11844
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 6738 11676 6748 11732
rect 6804 11676 7868 11732
rect 7924 11676 7934 11732
rect 8418 11676 8428 11732
rect 8484 11676 8820 11732
rect 19282 11676 19292 11732
rect 19348 11676 20412 11732
rect 20468 11676 20478 11732
rect 24658 11676 24668 11732
rect 24724 11676 26292 11732
rect 41010 11676 41020 11732
rect 41076 11676 44716 11732
rect 44772 11676 46172 11732
rect 46228 11676 46238 11732
rect 11890 11564 11900 11620
rect 11956 11564 13916 11620
rect 13972 11564 14588 11620
rect 14644 11564 14654 11620
rect 18274 11564 18284 11620
rect 18340 11564 19740 11620
rect 19796 11564 19806 11620
rect 20738 11564 20748 11620
rect 20804 11564 21084 11620
rect 21140 11564 25340 11620
rect 25396 11564 25406 11620
rect 20748 11508 20804 11564
rect 12338 11452 12348 11508
rect 12404 11452 14252 11508
rect 14308 11452 14318 11508
rect 16314 11452 16324 11508
rect 16380 11452 16940 11508
rect 16996 11452 20804 11508
rect 25442 11452 25452 11508
rect 25508 11452 25676 11508
rect 25732 11452 26124 11508
rect 26180 11452 26190 11508
rect 28466 11452 28476 11508
rect 28532 11452 29596 11508
rect 29652 11452 29662 11508
rect 30930 11452 30940 11508
rect 30996 11452 31724 11508
rect 31780 11452 31790 11508
rect 35970 11452 35980 11508
rect 36036 11452 36046 11508
rect 37762 11452 37772 11508
rect 37828 11452 38220 11508
rect 38276 11452 38286 11508
rect 35980 11396 36036 11452
rect 2706 11340 2716 11396
rect 2772 11340 3948 11396
rect 4004 11340 4014 11396
rect 6290 11340 6300 11396
rect 6356 11340 7532 11396
rect 7588 11340 7598 11396
rect 11890 11340 11900 11396
rect 11956 11340 11966 11396
rect 13178 11340 13188 11396
rect 13244 11340 13804 11396
rect 13860 11340 14364 11396
rect 14420 11340 14430 11396
rect 19004 11340 19014 11396
rect 19070 11340 20412 11396
rect 20468 11340 20478 11396
rect 21970 11340 21980 11396
rect 22036 11340 25340 11396
rect 25396 11340 25406 11396
rect 30818 11340 30828 11396
rect 30884 11340 31836 11396
rect 31892 11340 31902 11396
rect 35980 11340 36204 11396
rect 36260 11340 36876 11396
rect 36932 11340 37996 11396
rect 38052 11340 38062 11396
rect 46610 11340 46620 11396
rect 46676 11340 47964 11396
rect 48020 11340 48030 11396
rect 11900 11284 11956 11340
rect 3378 11228 3388 11284
rect 3444 11228 4060 11284
rect 4116 11228 4126 11284
rect 8194 11228 8204 11284
rect 8260 11228 9212 11284
rect 9268 11228 10444 11284
rect 10500 11228 11956 11284
rect 12562 11228 12572 11284
rect 12628 11228 13524 11284
rect 13580 11228 13590 11284
rect 21858 11228 21868 11284
rect 21924 11228 22092 11284
rect 22148 11228 22158 11284
rect 31154 11228 31164 11284
rect 31220 11228 33628 11284
rect 33684 11228 34412 11284
rect 34468 11228 34478 11284
rect 7858 11116 7868 11172
rect 7924 11116 8876 11172
rect 8932 11116 8942 11172
rect 11218 11116 11228 11172
rect 11284 11116 11564 11172
rect 11620 11116 11900 11172
rect 11956 11116 11966 11172
rect 16650 11116 16660 11172
rect 16716 11116 17612 11172
rect 17668 11116 17678 11172
rect 37986 11116 37996 11172
rect 38052 11116 38668 11172
rect 38724 11116 38734 11172
rect 42438 11116 42476 11172
rect 42532 11116 42542 11172
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 24780 10892 34356 10948
rect 34412 10892 34422 10948
rect 24780 10836 24836 10892
rect 3154 10780 3164 10836
rect 3220 10780 4284 10836
rect 4340 10780 5404 10836
rect 5460 10780 5964 10836
rect 6020 10780 6030 10836
rect 8082 10780 8092 10836
rect 8148 10780 9324 10836
rect 9380 10780 9390 10836
rect 12562 10780 12572 10836
rect 12628 10780 12638 10836
rect 17266 10780 17276 10836
rect 17332 10780 19002 10836
rect 19058 10780 20338 10836
rect 20394 10780 21678 10836
rect 21734 10780 21744 10836
rect 24164 10780 24174 10836
rect 24230 10780 24780 10836
rect 24836 10780 24846 10836
rect 26562 10780 26572 10836
rect 26628 10780 27804 10836
rect 27860 10780 27870 10836
rect 5282 10668 5292 10724
rect 5348 10668 5628 10724
rect 5684 10668 6188 10724
rect 6244 10668 6254 10724
rect 11218 10668 11228 10724
rect 11284 10668 11788 10724
rect 11844 10668 11854 10724
rect 4050 10556 4060 10612
rect 4116 10556 4788 10612
rect 4844 10556 5852 10612
rect 5908 10556 5918 10612
rect 8418 10556 8428 10612
rect 8484 10556 9660 10612
rect 9716 10556 9726 10612
rect 6290 10332 6300 10388
rect 6356 10332 6692 10388
rect 6748 10332 6758 10388
rect 12572 10276 12628 10780
rect 17546 10668 17556 10724
rect 17612 10668 18620 10724
rect 18676 10668 18686 10724
rect 20514 10668 20524 10724
rect 20580 10668 20972 10724
rect 21028 10668 21532 10724
rect 21588 10668 21980 10724
rect 22036 10668 24332 10724
rect 24388 10668 24398 10724
rect 31826 10668 31836 10724
rect 31892 10668 33180 10724
rect 33236 10668 33246 10724
rect 35690 10668 35700 10724
rect 35756 10668 38892 10724
rect 38948 10668 39676 10724
rect 39732 10668 40012 10724
rect 40068 10668 40078 10724
rect 46834 10668 46844 10724
rect 46900 10668 48468 10724
rect 17938 10556 17948 10612
rect 18004 10556 18732 10612
rect 18788 10556 18798 10612
rect 19170 10556 19180 10612
rect 19236 10556 20636 10612
rect 20692 10556 20702 10612
rect 22866 10556 22876 10612
rect 22932 10556 24444 10612
rect 24500 10556 24510 10612
rect 25442 10556 25452 10612
rect 25508 10556 26348 10612
rect 26404 10556 26414 10612
rect 28130 10556 28140 10612
rect 28196 10556 29260 10612
rect 29316 10556 29326 10612
rect 14802 10444 14812 10500
rect 14868 10444 17724 10500
rect 17780 10444 17790 10500
rect 18050 10444 18060 10500
rect 18116 10444 19292 10500
rect 19348 10444 19358 10500
rect 20412 10444 21420 10500
rect 21476 10444 26516 10500
rect 26572 10444 26582 10500
rect 20412 10388 20468 10444
rect 32508 10388 32564 10668
rect 48412 10612 48468 10668
rect 50200 10612 51000 10640
rect 38210 10556 38220 10612
rect 38276 10556 41244 10612
rect 41300 10556 41310 10612
rect 42354 10556 42364 10612
rect 42420 10556 43708 10612
rect 43764 10556 43774 10612
rect 44370 10556 44380 10612
rect 44436 10556 47404 10612
rect 47460 10556 48244 10612
rect 48300 10556 48310 10612
rect 48412 10556 51000 10612
rect 50200 10528 51000 10556
rect 39330 10444 39340 10500
rect 39396 10444 40908 10500
rect 40964 10444 40974 10500
rect 44482 10444 44492 10500
rect 44548 10444 48524 10500
rect 48580 10444 48590 10500
rect 20402 10332 20412 10388
rect 20468 10332 20478 10388
rect 32498 10332 32508 10388
rect 32564 10332 32574 10388
rect 33618 10332 33628 10388
rect 33684 10332 35308 10388
rect 35364 10332 35374 10388
rect 38546 10332 38556 10388
rect 38612 10332 39228 10388
rect 39284 10332 39732 10388
rect 44706 10332 44716 10388
rect 44772 10332 46060 10388
rect 46116 10332 46126 10388
rect 47394 10332 47404 10388
rect 47460 10332 48972 10388
rect 49028 10332 49038 10388
rect 12226 10220 12236 10276
rect 12292 10220 12628 10276
rect 20178 10220 20188 10276
rect 20244 10220 23100 10276
rect 23156 10220 23166 10276
rect 38098 10220 38108 10276
rect 38164 10220 39340 10276
rect 39396 10220 39406 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 39676 10164 39732 10332
rect 18274 10108 18284 10164
rect 18340 10108 18956 10164
rect 19012 10108 19022 10164
rect 34346 10108 34356 10164
rect 34412 10108 35028 10164
rect 36978 10108 36988 10164
rect 37044 10108 38668 10164
rect 38724 10108 38734 10164
rect 39666 10108 39676 10164
rect 39732 10108 41020 10164
rect 41076 10108 41086 10164
rect 46162 10108 46172 10164
rect 46228 10108 48636 10164
rect 48692 10108 48702 10164
rect 34972 10052 35028 10108
rect 3714 9996 3724 10052
rect 3780 9996 5572 10052
rect 5628 9996 5638 10052
rect 34972 9996 35252 10052
rect 35308 9996 35318 10052
rect 35858 9996 35868 10052
rect 35924 9996 37156 10052
rect 37212 9996 37772 10052
rect 37828 9996 37838 10052
rect 42858 9996 42868 10052
rect 42924 9996 45500 10052
rect 45556 9996 45566 10052
rect 4722 9884 4732 9940
rect 4788 9884 6412 9940
rect 6468 9884 6478 9940
rect 10098 9884 10108 9940
rect 10164 9884 12348 9940
rect 12404 9884 12414 9940
rect 22642 9884 22652 9940
rect 22708 9884 23660 9940
rect 23716 9884 23726 9940
rect 35410 9884 35420 9940
rect 35476 9884 35980 9940
rect 36036 9884 38332 9940
rect 38388 9884 38398 9940
rect 40282 9884 40292 9940
rect 40348 9884 41916 9940
rect 41972 9884 41982 9940
rect 44146 9884 44156 9940
rect 44212 9884 44716 9940
rect 44772 9884 44782 9940
rect 2706 9772 2716 9828
rect 2772 9772 3612 9828
rect 3668 9772 3678 9828
rect 8392 9772 8402 9828
rect 8458 9772 10780 9828
rect 10836 9772 10846 9828
rect 16706 9772 16716 9828
rect 16772 9772 17724 9828
rect 17780 9772 17790 9828
rect 19282 9772 19292 9828
rect 19348 9772 21868 9828
rect 21924 9772 22092 9828
rect 22148 9772 22158 9828
rect 28242 9772 28252 9828
rect 28308 9772 29148 9828
rect 29204 9772 29214 9828
rect 41010 9772 41020 9828
rect 41076 9772 43316 9828
rect 43372 9772 43382 9828
rect 45602 9772 45612 9828
rect 45668 9772 46060 9828
rect 46116 9772 48188 9828
rect 48244 9772 49308 9828
rect 49364 9772 49374 9828
rect 6402 9660 6412 9716
rect 6468 9660 8092 9716
rect 8148 9660 8158 9716
rect 14802 9660 14812 9716
rect 14868 9660 19516 9716
rect 19572 9660 19582 9716
rect 20626 9660 20636 9716
rect 20692 9660 21308 9716
rect 21364 9660 21374 9716
rect 31602 9660 31612 9716
rect 31668 9660 33292 9716
rect 33348 9660 33358 9716
rect 40002 9660 40012 9716
rect 40068 9660 40852 9716
rect 40908 9660 44156 9716
rect 44212 9660 44222 9716
rect 17042 9548 17052 9604
rect 17108 9548 18060 9604
rect 18116 9548 18126 9604
rect 41570 9548 41580 9604
rect 41636 9548 42252 9604
rect 42308 9548 42318 9604
rect 42466 9548 42476 9604
rect 42532 9548 43260 9604
rect 43316 9548 44996 9604
rect 45052 9548 45062 9604
rect 20626 9436 20636 9492
rect 20692 9436 22316 9492
rect 22372 9436 22876 9492
rect 22932 9436 23324 9492
rect 23380 9436 23390 9492
rect 38994 9436 39004 9492
rect 39060 9436 42868 9492
rect 42924 9436 42934 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 5808 9212 5818 9268
rect 5874 9212 6580 9268
rect 6636 9212 7084 9268
rect 7140 9212 7150 9268
rect 15138 9212 15148 9268
rect 15204 9212 19404 9268
rect 19460 9212 19470 9268
rect 40114 9212 40124 9268
rect 40180 9212 41132 9268
rect 41188 9212 41198 9268
rect 18722 9100 18732 9156
rect 18788 9100 19908 9156
rect 19964 9100 19974 9156
rect 39788 9100 40572 9156
rect 40628 9100 43148 9156
rect 43204 9100 43214 9156
rect 43474 9100 43484 9156
rect 43540 9100 43820 9156
rect 43876 9100 44268 9156
rect 44324 9100 44334 9156
rect 39788 9044 39844 9100
rect 4890 8988 4900 9044
rect 4956 8988 5628 9044
rect 5684 8988 6076 9044
rect 6132 8988 6142 9044
rect 7410 8988 7420 9044
rect 7476 8988 7868 9044
rect 7924 8988 7934 9044
rect 11554 8988 11564 9044
rect 11620 8988 12796 9044
rect 12852 8988 12862 9044
rect 18050 8988 18060 9044
rect 18116 8988 19740 9044
rect 19796 8988 19806 9044
rect 28018 8988 28028 9044
rect 28084 8988 30604 9044
rect 30660 8988 30670 9044
rect 38770 8988 38780 9044
rect 38836 8988 39788 9044
rect 39844 8988 39854 9044
rect 40226 8988 40236 9044
rect 40292 8988 43988 9044
rect 44044 8988 44054 9044
rect 16706 8876 16716 8932
rect 16772 8876 18284 8932
rect 18340 8876 18350 8932
rect 24098 8876 24108 8932
rect 24164 8876 25116 8932
rect 25172 8876 26684 8932
rect 26740 8876 28924 8932
rect 28980 8876 28990 8932
rect 8642 8764 8652 8820
rect 8708 8764 10444 8820
rect 10500 8764 10510 8820
rect 24322 8764 24332 8820
rect 24388 8764 25452 8820
rect 25508 8764 25518 8820
rect 35634 8764 35644 8820
rect 35700 8764 35868 8820
rect 35924 8764 35934 8820
rect 44706 8764 44716 8820
rect 44772 8764 48636 8820
rect 48692 8764 48702 8820
rect 3378 8652 3388 8708
rect 3444 8652 3724 8708
rect 3780 8652 4284 8708
rect 4340 8652 4350 8708
rect 37538 8652 37548 8708
rect 37604 8652 39116 8708
rect 39172 8652 39182 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 14802 8540 14812 8596
rect 14868 8540 17612 8596
rect 17668 8540 17678 8596
rect 31892 8540 33180 8596
rect 33236 8540 33246 8596
rect 31892 8484 31948 8540
rect 3602 8428 3612 8484
rect 3668 8428 4732 8484
rect 4788 8428 4798 8484
rect 21858 8428 21868 8484
rect 21980 8428 21990 8484
rect 23314 8428 23324 8484
rect 23380 8428 25116 8484
rect 25172 8428 25182 8484
rect 25442 8428 25452 8484
rect 25508 8428 27132 8484
rect 27188 8428 28028 8484
rect 28084 8428 28094 8484
rect 31490 8428 31500 8484
rect 31556 8428 31948 8484
rect 2370 8316 2380 8372
rect 2436 8316 4956 8372
rect 5012 8316 5022 8372
rect 19394 8316 19404 8372
rect 19460 8316 20188 8372
rect 20244 8316 20254 8372
rect 32396 8260 32452 8540
rect 43810 8428 43820 8484
rect 43876 8428 48972 8484
rect 49028 8428 49038 8484
rect 43026 8316 43036 8372
rect 43092 8316 44828 8372
rect 44884 8316 44894 8372
rect 7746 8204 7756 8260
rect 7812 8204 10668 8260
rect 10724 8204 10734 8260
rect 12338 8204 12348 8260
rect 12404 8204 12414 8260
rect 16146 8204 16156 8260
rect 16212 8204 18620 8260
rect 18676 8204 21588 8260
rect 21644 8204 22316 8260
rect 22372 8204 26964 8260
rect 27020 8204 27030 8260
rect 32386 8204 32396 8260
rect 32452 8204 32462 8260
rect 34178 8204 34188 8260
rect 34244 8204 34748 8260
rect 34804 8204 34814 8260
rect 34906 8204 34916 8260
rect 34972 8204 35644 8260
rect 35700 8204 35710 8260
rect 37660 8204 38108 8260
rect 38164 8204 38174 8260
rect 38490 8204 38500 8260
rect 38556 8204 39004 8260
rect 39060 8204 39070 8260
rect 43362 8204 43372 8260
rect 43428 8204 43596 8260
rect 43652 8204 45276 8260
rect 45332 8204 48748 8260
rect 48804 8204 48814 8260
rect 12348 8148 12404 8204
rect 37660 8148 37716 8204
rect 10098 8092 10108 8148
rect 10164 8092 10892 8148
rect 10948 8092 10958 8148
rect 12348 8092 16044 8148
rect 16100 8092 16110 8148
rect 19842 8092 19852 8148
rect 19908 8092 20412 8148
rect 20468 8092 20860 8148
rect 20916 8092 20926 8148
rect 23986 8092 23996 8148
rect 24052 8092 25508 8148
rect 25564 8092 25574 8148
rect 33506 8092 33516 8148
rect 33572 8092 37716 8148
rect 38210 8092 38220 8148
rect 38276 8092 39788 8148
rect 39844 8092 39854 8148
rect 44594 8092 44604 8148
rect 44660 8092 45500 8148
rect 45556 8092 46284 8148
rect 46340 8092 46350 8148
rect 38556 8036 38612 8092
rect 3994 7980 4004 8036
rect 4060 7980 4284 8036
rect 4340 7980 4350 8036
rect 18386 7980 18396 8036
rect 18452 7980 20524 8036
rect 20580 7980 20590 8036
rect 38546 7980 38556 8036
rect 38612 7980 38622 8036
rect 44370 7980 44380 8036
rect 44436 7980 45052 8036
rect 45108 7980 45118 8036
rect 48850 7868 48860 7924
rect 48916 7868 49196 7924
rect 49252 7868 49262 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 45490 7756 45500 7812
rect 45556 7756 45724 7812
rect 45780 7756 46620 7812
rect 46676 7756 46686 7812
rect 1586 7644 1596 7700
rect 1652 7644 2268 7700
rect 2324 7644 3724 7700
rect 3780 7644 5852 7700
rect 5908 7644 7420 7700
rect 7476 7644 7486 7700
rect 9874 7644 9884 7700
rect 9940 7644 11228 7700
rect 11284 7644 11294 7700
rect 34178 7644 34188 7700
rect 34244 7644 38312 7700
rect 38368 7644 38378 7700
rect 8194 7532 8204 7588
rect 8260 7532 8652 7588
rect 8708 7532 8718 7588
rect 10434 7532 10444 7588
rect 10500 7532 11844 7588
rect 11900 7532 12292 7588
rect 12348 7532 13448 7588
rect 13504 7532 13514 7588
rect 20290 7532 20300 7588
rect 20356 7532 21084 7588
rect 21140 7532 21150 7588
rect 29250 7532 29260 7588
rect 29316 7532 31276 7588
rect 31332 7532 31612 7588
rect 31668 7532 31678 7588
rect 43698 7532 43708 7588
rect 43764 7532 45276 7588
rect 45332 7532 45342 7588
rect 8082 7420 8092 7476
rect 8148 7420 9660 7476
rect 9716 7420 9726 7476
rect 19730 7420 19740 7476
rect 19796 7420 20636 7476
rect 20692 7420 21756 7476
rect 21812 7420 21822 7476
rect 27458 7420 27468 7476
rect 27524 7420 28364 7476
rect 28420 7420 29484 7476
rect 29540 7420 29550 7476
rect 30706 7420 30716 7476
rect 30772 7420 31780 7476
rect 31836 7420 31846 7476
rect 34850 7420 34860 7476
rect 34916 7420 35420 7476
rect 35476 7420 36316 7476
rect 36372 7420 36382 7476
rect 36530 7420 36540 7476
rect 36596 7420 37044 7476
rect 37100 7420 37110 7476
rect 44482 7420 44492 7476
rect 44548 7420 44558 7476
rect 44492 7364 44548 7420
rect 10098 7308 10108 7364
rect 10164 7308 11116 7364
rect 11172 7308 11182 7364
rect 34234 7308 34244 7364
rect 34300 7308 38668 7364
rect 38724 7308 39172 7364
rect 39228 7308 43036 7364
rect 43092 7308 45724 7364
rect 45780 7308 45790 7364
rect 38612 7196 39900 7252
rect 39956 7196 41244 7252
rect 41300 7196 41310 7252
rect 44538 7196 44548 7252
rect 44604 7196 47292 7252
rect 47348 7196 47358 7252
rect 33170 7084 33180 7140
rect 33236 7084 34972 7140
rect 35028 7084 35038 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 38612 7028 38668 7196
rect 38882 7084 38892 7140
rect 38948 7084 39564 7140
rect 39620 7084 39630 7140
rect 7746 6972 7756 7028
rect 7812 6972 8092 7028
rect 8148 6972 8158 7028
rect 37650 6972 37660 7028
rect 37716 6972 38312 7028
rect 38368 6972 38668 7028
rect 4274 6860 4284 6916
rect 4340 6860 7084 6916
rect 7140 6860 10556 6916
rect 10612 6860 10622 6916
rect 37034 6860 37044 6916
rect 37100 6860 39228 6916
rect 39284 6860 43260 6916
rect 43316 6860 43326 6916
rect 4946 6748 4956 6804
rect 5012 6748 6300 6804
rect 6356 6748 6366 6804
rect 9762 6748 9772 6804
rect 9828 6748 10780 6804
rect 10836 6748 10846 6804
rect 11452 6748 12236 6804
rect 12292 6748 12302 6804
rect 13682 6748 13692 6804
rect 13748 6748 14140 6804
rect 14196 6748 14206 6804
rect 19394 6748 19404 6804
rect 19460 6748 20748 6804
rect 20804 6748 20814 6804
rect 25330 6748 25340 6804
rect 25396 6748 26460 6804
rect 26516 6748 28644 6804
rect 28700 6748 28710 6804
rect 28812 6748 29372 6804
rect 29428 6748 33404 6804
rect 33460 6748 33470 6804
rect 34962 6748 34972 6804
rect 35028 6748 36092 6804
rect 36148 6748 36158 6804
rect 39106 6748 39116 6804
rect 39172 6748 40460 6804
rect 40516 6748 40526 6804
rect 45490 6748 45500 6804
rect 45556 6748 46396 6804
rect 46452 6748 46462 6804
rect 2818 6636 2828 6692
rect 2884 6636 5740 6692
rect 5796 6636 5806 6692
rect 6066 6636 6076 6692
rect 6132 6636 6916 6692
rect 6972 6636 6982 6692
rect 7858 6636 7868 6692
rect 7924 6636 8428 6692
rect 8484 6636 8494 6692
rect 3826 6524 3836 6580
rect 3892 6524 5964 6580
rect 6020 6524 6030 6580
rect 11452 6468 11508 6748
rect 16706 6636 16716 6692
rect 16772 6636 17612 6692
rect 17668 6636 17678 6692
rect 19618 6636 19628 6692
rect 19684 6636 19852 6692
rect 19908 6636 20300 6692
rect 20356 6636 20366 6692
rect 23426 6636 23436 6692
rect 23492 6636 23884 6692
rect 23940 6636 23950 6692
rect 24322 6636 24332 6692
rect 24388 6636 25452 6692
rect 25508 6636 25518 6692
rect 26786 6636 26796 6692
rect 26852 6636 27468 6692
rect 27524 6636 27534 6692
rect 28812 6580 28868 6748
rect 29922 6636 29932 6692
rect 29988 6636 30492 6692
rect 30548 6636 30558 6692
rect 31826 6636 31836 6692
rect 31892 6636 32340 6692
rect 32396 6636 32406 6692
rect 32508 6636 32844 6692
rect 32900 6636 33292 6692
rect 33348 6636 35756 6692
rect 35812 6636 35822 6692
rect 37538 6636 37548 6692
rect 37604 6636 38556 6692
rect 38612 6636 38622 6692
rect 39330 6636 39340 6692
rect 39396 6636 40348 6692
rect 40404 6636 40414 6692
rect 41234 6636 41244 6692
rect 41300 6636 47068 6692
rect 47124 6636 48300 6692
rect 48356 6636 49308 6692
rect 49364 6636 49374 6692
rect 32508 6580 32564 6636
rect 17154 6524 17164 6580
rect 17220 6524 18116 6580
rect 18172 6524 20412 6580
rect 20468 6524 20478 6580
rect 27010 6524 27020 6580
rect 27076 6524 28868 6580
rect 30146 6524 30156 6580
rect 30212 6524 30716 6580
rect 30772 6524 30782 6580
rect 31892 6524 32564 6580
rect 38098 6524 38108 6580
rect 38164 6524 41356 6580
rect 41412 6524 41422 6580
rect 44594 6524 44604 6580
rect 44660 6524 46620 6580
rect 46676 6524 47908 6580
rect 31892 6468 31948 6524
rect 47852 6468 47908 6524
rect 3602 6412 3612 6468
rect 3668 6412 5628 6468
rect 5684 6412 5694 6468
rect 11442 6412 11452 6468
rect 11508 6412 11518 6468
rect 16034 6412 16044 6468
rect 16100 6412 21196 6468
rect 21252 6412 21262 6468
rect 21522 6412 21532 6468
rect 21588 6412 22932 6468
rect 22988 6412 22998 6468
rect 25386 6412 25396 6468
rect 25452 6412 31948 6468
rect 37426 6412 37436 6468
rect 37492 6412 39004 6468
rect 39060 6412 39070 6468
rect 45490 6412 45500 6468
rect 45556 6412 46116 6468
rect 46172 6412 46182 6468
rect 47842 6412 47852 6468
rect 47908 6412 47918 6468
rect 4956 5908 5012 6412
rect 50200 6356 51000 6384
rect 6290 6300 6300 6356
rect 6356 6300 6860 6356
rect 6916 6300 7532 6356
rect 7588 6300 7980 6356
rect 8036 6300 8046 6356
rect 8418 6300 8428 6356
rect 8484 6300 9548 6356
rect 9604 6300 9996 6356
rect 10052 6300 10062 6356
rect 16594 6300 16604 6356
rect 16660 6300 19068 6356
rect 19124 6300 19134 6356
rect 46946 6300 46956 6356
rect 47012 6300 51000 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50200 6272 51000 6300
rect 5730 6188 5740 6244
rect 5796 6188 6412 6244
rect 6468 6188 6478 6244
rect 42578 6188 42588 6244
rect 42644 6188 44100 6244
rect 44156 6188 44166 6244
rect 45378 6188 45388 6244
rect 45444 6188 45836 6244
rect 45892 6188 49196 6244
rect 49252 6188 49262 6244
rect 5618 6076 5628 6132
rect 5684 6076 6580 6132
rect 6636 6076 8540 6132
rect 8596 6076 9436 6132
rect 9492 6076 9502 6132
rect 16930 6076 16940 6132
rect 16996 6076 17500 6132
rect 17556 6076 17566 6132
rect 18330 6076 18340 6132
rect 18396 6076 20076 6132
rect 20132 6076 24556 6132
rect 24612 6076 25396 6132
rect 25452 6076 25462 6132
rect 25834 6076 25844 6132
rect 25900 6076 26516 6132
rect 26572 6076 26582 6132
rect 29586 6076 29596 6132
rect 29652 6076 30380 6132
rect 30436 6076 30446 6132
rect 43362 6076 43372 6132
rect 43428 6076 44660 6132
rect 47142 6076 47180 6132
rect 47236 6076 47246 6132
rect 47730 6076 47740 6132
rect 47796 6076 48412 6132
rect 48468 6076 48478 6132
rect 44604 6020 44660 6076
rect 4946 5852 4956 5908
rect 5012 5852 5022 5908
rect 6962 5852 6972 5908
rect 7028 5852 8092 5908
rect 8148 5852 8158 5908
rect 8372 5796 8428 6020
rect 8484 5964 8988 6020
rect 9044 5964 10220 6020
rect 10276 5964 10286 6020
rect 19394 5964 19404 6020
rect 19460 5964 23772 6020
rect 23828 5964 23838 6020
rect 39218 5964 39228 6020
rect 39284 5964 39900 6020
rect 39956 5964 39966 6020
rect 43698 5964 43708 6020
rect 43764 5964 44380 6020
rect 44436 5964 44446 6020
rect 44594 5964 44604 6020
rect 44660 5964 45164 6020
rect 45220 5964 45836 6020
rect 45892 5964 45902 6020
rect 9426 5852 9436 5908
rect 9492 5852 9772 5908
rect 9828 5852 10332 5908
rect 10388 5852 10398 5908
rect 15922 5852 15932 5908
rect 15988 5852 16492 5908
rect 16548 5852 16558 5908
rect 19058 5852 19068 5908
rect 19124 5852 22186 5908
rect 22242 5852 22252 5908
rect 27906 5852 27916 5908
rect 27972 5852 29260 5908
rect 29316 5852 29326 5908
rect 30258 5852 30268 5908
rect 30324 5852 31612 5908
rect 31668 5852 31678 5908
rect 33394 5852 33404 5908
rect 33460 5852 34188 5908
rect 34244 5852 34748 5908
rect 34804 5852 34814 5908
rect 43474 5852 43484 5908
rect 43540 5852 44492 5908
rect 44548 5852 44828 5908
rect 44884 5852 44894 5908
rect 47506 5852 47516 5908
rect 47572 5852 49084 5908
rect 49140 5852 49150 5908
rect 4610 5740 4620 5796
rect 4676 5740 6076 5796
rect 6132 5740 7140 5796
rect 7196 5740 7206 5796
rect 7298 5740 7308 5796
rect 7364 5740 7532 5796
rect 7588 5740 8428 5796
rect 32050 5740 32060 5796
rect 32116 5740 34300 5796
rect 34356 5740 34366 5796
rect 3042 5628 3052 5684
rect 3108 5628 4396 5684
rect 4452 5628 4462 5684
rect 7690 5628 7700 5684
rect 7756 5628 8428 5684
rect 8484 5628 8494 5684
rect 16818 5628 16828 5684
rect 16884 5628 17500 5684
rect 17556 5628 17836 5684
rect 17892 5628 17902 5684
rect 19058 5628 19068 5684
rect 19124 5628 20300 5684
rect 20356 5628 20366 5684
rect 38546 5628 38556 5684
rect 38612 5628 39452 5684
rect 39508 5628 41356 5684
rect 41412 5628 41422 5684
rect 41570 5628 41580 5684
rect 41636 5628 41646 5684
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 16258 5404 16268 5460
rect 16324 5404 16604 5460
rect 16660 5404 16670 5460
rect 31378 5404 31388 5460
rect 31444 5404 31724 5460
rect 31780 5404 31790 5460
rect 41580 5348 41636 5628
rect 46274 5516 46284 5572
rect 46340 5516 46956 5572
rect 47012 5516 47022 5572
rect 44034 5404 44044 5460
rect 44100 5404 44940 5460
rect 44996 5404 45006 5460
rect 7858 5292 7868 5348
rect 7924 5292 8876 5348
rect 8932 5292 9212 5348
rect 9268 5292 9996 5348
rect 10052 5292 10062 5348
rect 16370 5292 16380 5348
rect 16436 5292 16716 5348
rect 16772 5292 16782 5348
rect 41580 5292 41916 5348
rect 41972 5292 41982 5348
rect 45602 5292 45612 5348
rect 45668 5292 48412 5348
rect 48468 5292 48478 5348
rect 4946 5180 4956 5236
rect 5012 5180 5740 5236
rect 5796 5180 5806 5236
rect 7970 5180 7980 5236
rect 8036 5180 8652 5236
rect 8708 5180 8718 5236
rect 15362 5180 15372 5236
rect 15428 5180 17500 5236
rect 17556 5180 17566 5236
rect 20178 5180 20188 5236
rect 20244 5180 20636 5236
rect 20692 5180 28196 5236
rect 28252 5180 28262 5236
rect 28466 5180 28476 5236
rect 28532 5180 30716 5236
rect 30772 5180 30782 5236
rect 35634 5180 35644 5236
rect 35700 5180 37156 5236
rect 37212 5180 37222 5236
rect 38098 5180 38108 5236
rect 38164 5180 38892 5236
rect 38948 5180 38958 5236
rect 39330 5180 39340 5236
rect 39396 5180 43484 5236
rect 43540 5180 43550 5236
rect 44930 5180 44940 5236
rect 44996 5180 45388 5236
rect 45444 5180 45724 5236
rect 45780 5180 45790 5236
rect 46610 5180 46620 5236
rect 46676 5180 47964 5236
rect 48020 5180 48030 5236
rect 48178 5180 48188 5236
rect 48244 5180 49196 5236
rect 49252 5180 49262 5236
rect 7858 5068 7868 5124
rect 7924 5068 8540 5124
rect 8596 5068 8606 5124
rect 14018 5068 14028 5124
rect 14084 5068 16940 5124
rect 16996 5068 17006 5124
rect 17266 5068 17276 5124
rect 17332 5068 18508 5124
rect 18564 5068 18574 5124
rect 18946 5068 18956 5124
rect 19012 5068 19404 5124
rect 19460 5068 19470 5124
rect 20738 5068 20748 5124
rect 20804 5068 20814 5124
rect 23090 5068 23100 5124
rect 23156 5068 23772 5124
rect 23828 5068 23838 5124
rect 24434 5068 24444 5124
rect 24500 5068 25564 5124
rect 25620 5068 25630 5124
rect 26338 5068 26348 5124
rect 26404 5068 26908 5124
rect 26964 5068 27132 5124
rect 27188 5068 27468 5124
rect 27524 5068 29484 5124
rect 29540 5068 30492 5124
rect 30548 5068 31164 5124
rect 31220 5068 33628 5124
rect 33684 5068 35868 5124
rect 35924 5068 35934 5124
rect 38434 5068 38444 5124
rect 38500 5068 39452 5124
rect 39508 5068 39518 5124
rect 41234 5068 41244 5124
rect 41300 5068 47068 5124
rect 47124 5068 47134 5124
rect 47282 5068 47292 5124
rect 47348 5068 47628 5124
rect 47684 5068 48300 5124
rect 48356 5068 48366 5124
rect 20748 5012 20804 5068
rect 18722 4956 18732 5012
rect 18788 4956 20804 5012
rect 27906 4956 27916 5012
rect 27972 4956 29036 5012
rect 29092 4956 29102 5012
rect 32498 4956 32508 5012
rect 32564 4956 33964 5012
rect 34020 4956 34030 5012
rect 44706 4956 44716 5012
rect 44772 4956 48524 5012
rect 48580 4956 48590 5012
rect 15334 4844 15372 4900
rect 15428 4844 15438 4900
rect 17714 4844 17724 4900
rect 17780 4844 20188 4900
rect 20244 4844 20254 4900
rect 28186 4844 28196 4900
rect 28252 4844 28812 4900
rect 28868 4844 28878 4900
rect 31490 4844 31500 4900
rect 31556 4844 35084 4900
rect 35140 4844 35150 4900
rect 38994 4844 39004 4900
rect 39060 4844 43036 4900
rect 43092 4844 43102 4900
rect 44146 4844 44156 4900
rect 44212 4844 49140 4900
rect 49196 4844 49206 4900
rect 42354 4732 42364 4788
rect 42420 4732 45500 4788
rect 45556 4732 45566 4788
rect 46722 4732 46732 4788
rect 46788 4732 47180 4788
rect 47236 4732 47246 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 22922 4620 22932 4676
rect 22988 4620 23604 4676
rect 23660 4620 25396 4676
rect 25452 4620 25462 4676
rect 38210 4620 38220 4676
rect 38276 4620 39788 4676
rect 39844 4620 39854 4676
rect 14354 4508 14364 4564
rect 14420 4508 22186 4564
rect 22242 4508 22252 4564
rect 22530 4508 22540 4564
rect 22596 4508 26142 4564
rect 26198 4508 26208 4564
rect 15698 4396 15708 4452
rect 15764 4396 22858 4452
rect 22914 4396 22924 4452
rect 23762 4396 23772 4452
rect 23828 4396 25228 4452
rect 25284 4396 25788 4452
rect 25844 4396 25854 4452
rect 39218 4396 39228 4452
rect 39284 4396 42028 4452
rect 42084 4396 42094 4452
rect 6962 4284 6972 4340
rect 7028 4284 8316 4340
rect 8372 4284 8382 4340
rect 15026 4284 15036 4340
rect 15092 4284 18508 4340
rect 18564 4284 18574 4340
rect 25890 4284 25900 4340
rect 25956 4284 33180 4340
rect 33236 4284 33246 4340
rect 36754 4284 36764 4340
rect 36820 4284 40124 4340
rect 40180 4284 40190 4340
rect 16482 4172 16492 4228
rect 16548 4172 17444 4228
rect 17500 4172 18396 4228
rect 18452 4172 18462 4228
rect 37874 4172 37884 4228
rect 37940 4172 39116 4228
rect 39172 4172 39182 4228
rect 46834 4172 46844 4228
rect 46900 4172 48972 4228
rect 49028 4172 49038 4228
rect 34636 4060 43820 4116
rect 43876 4060 43886 4116
rect 34636 4004 34692 4060
rect 34626 3948 34636 4004
rect 34692 3948 34702 4004
rect 43922 3948 43932 4004
rect 43988 3948 45948 4004
rect 46004 3948 46014 4004
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 45798 3836 45836 3892
rect 45892 3836 45902 3892
rect 41794 3724 41804 3780
rect 41860 3724 42700 3780
rect 42756 3724 42766 3780
rect 46498 3724 46508 3780
rect 46564 3724 48300 3780
rect 48356 3724 48366 3780
rect 14690 3612 14700 3668
rect 14756 3612 17724 3668
rect 17780 3612 17790 3668
rect 17938 3612 17948 3668
rect 18004 3612 19628 3668
rect 19684 3612 20300 3668
rect 20356 3612 20366 3668
rect 20850 3612 20860 3668
rect 20916 3612 22092 3668
rect 22148 3612 22158 3668
rect 22418 3612 22428 3668
rect 22484 3612 24780 3668
rect 24836 3612 24846 3668
rect 29474 3612 29484 3668
rect 29540 3612 30604 3668
rect 30660 3612 30670 3668
rect 33394 3612 33404 3668
rect 33460 3612 36988 3668
rect 37044 3612 37054 3668
rect 37986 3612 37996 3668
rect 38052 3612 47628 3668
rect 47684 3612 47694 3668
rect 28802 3500 28812 3556
rect 28868 3500 29148 3556
rect 29204 3500 29214 3556
rect 29586 3500 29596 3556
rect 29652 3500 30156 3556
rect 30212 3500 30222 3556
rect 31602 3500 31612 3556
rect 31668 3500 32396 3556
rect 32452 3500 32462 3556
rect 35074 3500 35084 3556
rect 35140 3500 38668 3556
rect 38724 3500 38734 3556
rect 43754 3500 43764 3556
rect 43820 3500 47964 3556
rect 48020 3500 48030 3556
rect 1138 3388 1148 3444
rect 1204 3388 1764 3444
rect 1820 3388 1830 3444
rect 4722 3388 4732 3444
rect 4788 3388 5572 3444
rect 5628 3388 5638 3444
rect 20122 3388 20132 3444
rect 20188 3388 22652 3444
rect 22708 3388 22718 3444
rect 27738 3388 27748 3444
rect 27804 3388 29820 3444
rect 29876 3388 29886 3444
rect 36978 3388 36988 3444
rect 37044 3388 40572 3444
rect 40628 3388 40638 3444
rect 44258 3388 44268 3444
rect 44324 3388 44334 3444
rect 45154 3388 45164 3444
rect 45220 3388 45230 3444
rect 45322 3388 45332 3444
rect 45388 3388 46732 3444
rect 46788 3388 46798 3444
rect 44268 3332 44324 3388
rect 45164 3332 45220 3388
rect 44268 3276 46620 3332
rect 46676 3276 46686 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50200 2100 51000 2128
rect 44706 2044 44716 2100
rect 44772 2044 51000 2100
rect 50200 2016 51000 2044
<< via3 >>
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 43708 47404 43764 47460
rect 47628 47180 47684 47236
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 31164 46956 31220 47012
rect 43708 46956 43764 47012
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 31164 45948 31220 46004
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 42812 44380 42868 44436
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 40908 43484 40964 43540
rect 45948 43260 46004 43316
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 42812 43036 42868 43092
rect 12236 42700 12292 42756
rect 12236 42476 12292 42532
rect 40908 42476 40964 42532
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 34524 41692 34580 41748
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 27692 40796 27748 40852
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 21980 40684 22036 40740
rect 34524 40572 34580 40628
rect 34972 40572 35028 40628
rect 21980 40012 22036 40068
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 27692 39900 27748 39956
rect 33740 39564 33796 39620
rect 9212 39228 9268 39284
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 20188 39004 20244 39060
rect 47180 39004 47236 39060
rect 33740 38556 33796 38612
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 44940 38332 44996 38388
rect 45164 37996 45220 38052
rect 12236 37772 12292 37828
rect 33964 37772 34020 37828
rect 45164 37772 45220 37828
rect 9212 37660 9268 37716
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 34860 37548 34916 37604
rect 47180 37548 47236 37604
rect 44940 37212 44996 37268
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35644 36988 35700 37044
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 33964 36428 34020 36484
rect 45164 36428 45220 36484
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 34860 35756 34916 35812
rect 41468 35756 41524 35812
rect 47292 35756 47348 35812
rect 20188 35532 20244 35588
rect 22876 35308 22932 35364
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 41468 35196 41524 35252
rect 17724 34860 17780 34916
rect 18620 34524 18676 34580
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 18060 34412 18116 34468
rect 18508 34188 18564 34244
rect 20524 33964 20580 34020
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 18060 33628 18116 33684
rect 35644 33516 35700 33572
rect 47292 33516 47348 33572
rect 18620 33404 18676 33460
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 11900 32732 11956 32788
rect 38220 32396 38276 32452
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19180 32060 19236 32116
rect 34300 32060 34356 32116
rect 17836 31948 17892 32004
rect 21644 31836 21700 31892
rect 22876 31724 22932 31780
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 47180 31276 47236 31332
rect 38108 31164 38164 31220
rect 21644 30716 21700 30772
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 17724 30492 17780 30548
rect 17836 30268 17892 30324
rect 20524 30268 20580 30324
rect 26796 30268 26852 30324
rect 19180 30044 19236 30100
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 38220 29484 38276 29540
rect 11900 29036 11956 29092
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 36988 28588 37044 28644
rect 26796 28364 26852 28420
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 47628 28028 47684 28084
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 34300 26796 34356 26852
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 38108 26572 38164 26628
rect 5180 26236 5236 26292
rect 38668 26236 38724 26292
rect 18508 25900 18564 25956
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 37772 25452 37828 25508
rect 38668 25228 38724 25284
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 34860 24220 34916 24276
rect 37772 24108 37828 24164
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 34972 23436 35028 23492
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 36988 20412 37044 20468
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 45948 20076 46004 20132
rect 33964 19852 34020 19908
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 5180 15260 5236 15316
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 24780 13244 24836 13300
rect 5180 13132 5236 13188
rect 24780 12684 24836 12740
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 8428 12012 8484 12068
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 42476 11788 42532 11844
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 8428 11676 8484 11732
rect 21868 11228 21924 11284
rect 42476 11116 42532 11172
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 21868 9772 21924 9828
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 21868 8428 21924 8484
rect 38108 8204 38164 8260
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 38108 6524 38164 6580
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 45836 6188 45892 6244
rect 47180 6076 47236 6132
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 15372 5180 15428 5236
rect 15372 4844 15428 4900
rect 47180 4732 47236 4788
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 45836 3836 45892 3892
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 47852 4768 47884
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 19808 47068 20128 47884
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 35168 47852 35488 47884
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 19808 45500 20128 47012
rect 31164 47012 31220 47022
rect 31164 46004 31220 46956
rect 31164 45938 31220 45948
rect 35168 46284 35488 47796
rect 43708 47460 43764 47470
rect 43708 47012 43764 47404
rect 43708 46946 43764 46956
rect 47628 47236 47684 47246
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 12236 42756 12292 42766
rect 12236 42532 12292 42700
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 9212 39284 9268 39294
rect 9212 37716 9268 39228
rect 12236 37828 12292 42476
rect 12236 37762 12292 37772
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 42812 44436 42868 44446
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 34524 41748 34580 41758
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 27692 40852 27748 40862
rect 19808 39228 20128 40740
rect 21980 40740 22036 40750
rect 21980 40068 22036 40684
rect 21980 40002 22036 40012
rect 27692 39956 27748 40796
rect 34524 40628 34580 41692
rect 35168 41580 35488 43092
rect 40908 43540 40964 43550
rect 40908 42532 40964 43484
rect 42812 43092 42868 44380
rect 42812 43026 42868 43036
rect 45948 43316 46004 43326
rect 40908 42466 40964 42476
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 34524 40562 34580 40572
rect 34972 40628 35028 40638
rect 27692 39890 27748 39900
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 9212 37650 9268 37660
rect 19808 37660 20128 39172
rect 33740 39620 33796 39630
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 17724 34916 17780 34926
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 11900 32788 11956 32798
rect 11900 29092 11956 32732
rect 17724 30548 17780 34860
rect 18620 34580 18676 34590
rect 18060 34468 18116 34478
rect 18060 33684 18116 34412
rect 18060 33618 18116 33628
rect 18508 34244 18564 34254
rect 17724 30482 17780 30492
rect 17836 32004 17892 32014
rect 17836 30324 17892 31948
rect 17836 30258 17892 30268
rect 11900 29026 11956 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 5180 26292 5236 26302
rect 5180 15316 5236 26236
rect 18508 25956 18564 34188
rect 18620 33460 18676 34524
rect 18620 33394 18676 33404
rect 19808 34524 20128 36036
rect 20188 39060 20244 39070
rect 20188 35588 20244 39004
rect 33740 38612 33796 39564
rect 33740 38546 33796 38556
rect 20188 35522 20244 35532
rect 33964 37828 34020 37838
rect 33964 36484 34020 37772
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 22876 35364 22932 35374
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19180 32116 19236 32126
rect 19180 30100 19236 32060
rect 19180 30034 19236 30044
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 18508 25890 18564 25900
rect 19808 29820 20128 31332
rect 20524 34020 20580 34030
rect 20524 30324 20580 33964
rect 21644 31892 21700 31902
rect 21644 30772 21700 31836
rect 22876 31780 22932 35308
rect 22876 31714 22932 31724
rect 21644 30706 21700 30716
rect 20524 30258 20580 30268
rect 26796 30324 26852 30334
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 26796 28420 26852 30268
rect 26796 28354 26852 28364
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 5180 13188 5236 15260
rect 5180 13122 5236 13132
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 33964 19908 34020 36428
rect 34860 37604 34916 37614
rect 34860 35812 34916 37548
rect 34300 32116 34356 32126
rect 34300 26852 34356 32060
rect 34300 26786 34356 26796
rect 34860 24276 34916 35756
rect 34860 24210 34916 24220
rect 34972 23492 35028 40572
rect 34972 23426 35028 23436
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 44940 38388 44996 38398
rect 44940 37268 44996 38332
rect 44940 37202 44996 37212
rect 45164 38052 45220 38062
rect 45164 37828 45220 37996
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35644 37044 35700 37054
rect 35644 33572 35700 36988
rect 45164 36484 45220 37772
rect 45164 36418 45220 36428
rect 41468 35812 41524 35822
rect 41468 35252 41524 35756
rect 41468 35186 41524 35196
rect 35644 33506 35700 33516
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 38220 32452 38276 32462
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 38108 31220 38164 31230
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 33964 19842 34020 19852
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 35168 19628 35488 21140
rect 36988 28644 37044 28654
rect 36988 20468 37044 28588
rect 38108 26628 38164 31164
rect 38220 29540 38276 32396
rect 38220 29474 38276 29484
rect 38108 26562 38164 26572
rect 38668 26292 38724 26302
rect 37772 25508 37828 25518
rect 37772 24164 37828 25452
rect 38668 25284 38724 26236
rect 38668 25218 38724 25228
rect 37772 24098 37828 24108
rect 36988 20402 37044 20412
rect 45948 20132 46004 43260
rect 47180 39060 47236 39070
rect 47180 37604 47236 39004
rect 47180 31332 47236 37548
rect 47292 35812 47348 35822
rect 47292 33572 47348 35756
rect 47292 33506 47348 33516
rect 47180 31266 47236 31276
rect 47628 28084 47684 47180
rect 47628 28018 47684 28028
rect 45948 20066 46004 20076
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 24780 13300 24836 13310
rect 24780 12740 24836 13244
rect 24780 12674 24836 12684
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 8428 12068 8484 12078
rect 8428 11732 8484 12012
rect 8428 11666 8484 11676
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 19808 11004 20128 12516
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 21868 11284 21924 11294
rect 21868 9828 21924 11228
rect 21868 8484 21924 9772
rect 21868 8418 21924 8428
rect 35168 10220 35488 11732
rect 42476 11844 42532 11854
rect 42476 11172 42532 11788
rect 42476 11106 42532 11116
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 15372 5236 15428 5246
rect 15372 4900 15428 5180
rect 15372 4834 15428 4844
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 38108 8260 38164 8270
rect 38108 6580 38164 8204
rect 38108 6514 38164 6524
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 45836 6244 45892 6254
rect 45836 3892 45892 6188
rect 47180 6132 47236 6142
rect 47180 4788 47236 6076
rect 47180 4722 47236 4732
rect 45836 3826 45892 3836
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1271_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751534193
transform 1 0 21168 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1272_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751914308
transform -1 0 23296 0 1 4704
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1273_
timestamp 1751534193
transform -1 0 14448 0 -1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1274_
timestamp 1751914308
transform -1 0 23968 0 -1 4704
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1275_
timestamp 1751534193
transform -1 0 15792 0 -1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1276_
timestamp 1751914308
transform -1 0 23296 0 -1 6272
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1277_
timestamp 1751534193
transform -1 0 19152 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1278_
timestamp 1751914308
transform 1 0 25088 0 -1 4704
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1279_
timestamp 1751534193
transform -1 0 22512 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_4  _1280_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753277880
transform -1 0 44464 0 1 20384
box -86 -86 1990 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _1281_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751905124
transform -1 0 30912 0 1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1282_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751889808
transform 1 0 27104 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1283_
timestamp 1751889808
transform -1 0 35616 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _1284_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1752345181
transform 1 0 31472 0 -1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_4  _1285_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753432499
transform 1 0 31472 0 1 18816
box -86 -86 2214 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1286_
timestamp 1751889808
transform 1 0 29456 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1287_
timestamp 1751889808
transform 1 0 26768 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1288_
timestamp 1751534193
transform -1 0 29008 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _1289_
timestamp 1751905124
transform -1 0 33936 0 1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _1290_
timestamp 1752345181
transform 1 0 30800 0 -1 21952
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_4  _1291_
timestamp 1753432499
transform -1 0 32816 0 1 20384
box -86 -86 2214 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1292_
timestamp 1751889808
transform 1 0 34608 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1293_
timestamp 1751889808
transform -1 0 31472 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _1294_
timestamp 1751905124
transform 1 0 30352 0 1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _1295_
timestamp 1752345181
transform -1 0 32144 0 -1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1296_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753371985
transform 1 0 29792 0 -1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1297_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753277515
transform 1 0 31472 0 1 9408
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1298_
timestamp 1753277515
transform 1 0 32256 0 1 7840
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1299_
timestamp 1751534193
transform 1 0 41328 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1300_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753272495
transform 1 0 33040 0 1 9408
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1301_
timestamp 1751534193
transform 1 0 33824 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1302_
timestamp 1751534193
transform 1 0 7504 0 1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _1303_
timestamp 1752345181
transform 1 0 11424 0 -1 12544
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1304_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1752061876
transform -1 0 11200 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1305_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532043
transform 1 0 7840 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1306_
timestamp 1751532043
transform -1 0 7952 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1307_
timestamp 1751532043
transform 1 0 6048 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1308_
timestamp 1751532043
transform 1 0 5824 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1309_
timestamp 1751532043
transform -1 0 9072 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1310_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753960525
transform -1 0 6832 0 1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1311_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751740063
transform 1 0 5824 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1312_
timestamp 1751740063
transform 1 0 6496 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1313_
timestamp 1751532043
transform -1 0 9968 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1314_
timestamp 1753960525
transform 1 0 6384 0 1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1315_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751531619
transform 1 0 6720 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1316_
timestamp 1751531619
transform -1 0 7840 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1317_
timestamp 1751889808
transform 1 0 9184 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1318_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753182340
transform 1 0 10416 0 1 7840
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1319_
timestamp 1751889808
transform 1 0 6160 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1320_
timestamp 1753182340
transform 1 0 5488 0 1 9408
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _1321_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753891287
transform 1 0 7168 0 1 9408
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1322_
timestamp 1751534193
transform 1 0 8512 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1323_
timestamp 1751534193
transform -1 0 7504 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1324_
timestamp 1751740063
transform -1 0 4256 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1325_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751889408
transform 1 0 5488 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1326_
timestamp 1751740063
transform 1 0 6720 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1327_
timestamp 1753182340
transform 1 0 5488 0 1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1328_
timestamp 1751534193
transform -1 0 2912 0 1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1329_
timestamp 1751534193
transform -1 0 8288 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1330_
timestamp 1751534193
transform 1 0 8288 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1331_
timestamp 1751534193
transform -1 0 10080 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1332_
timestamp 1753277515
transform 1 0 6048 0 -1 31360
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1333_
timestamp 1751740063
transform 1 0 6944 0 -1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _1334_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753172561
transform -1 0 5264 0 1 29792
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1335_
timestamp 1753960525
transform 1 0 4816 0 -1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1336_
timestamp 1751531619
transform -1 0 5264 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1337_
timestamp 1751740063
transform 1 0 3024 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1338_
timestamp 1751532043
transform 1 0 7056 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1339_
timestamp 1751534193
transform -1 0 7504 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1340_
timestamp 1751740063
transform 1 0 2688 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1341_
timestamp 1751889808
transform 1 0 5152 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1342_
timestamp 1753371985
transform -1 0 6608 0 1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1343_
timestamp 1753277515
transform -1 0 4032 0 -1 28224
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1344_
timestamp 1751740063
transform 1 0 1680 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1345_
timestamp 1751532043
transform 1 0 4592 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1346_
timestamp 1753182340
transform 1 0 5488 0 1 26656
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1347_
timestamp 1751740063
transform -1 0 7504 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1348_
timestamp 1751889408
transform -1 0 5152 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1349_
timestamp 1753182340
transform -1 0 6720 0 1 25088
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1350_
timestamp 1751534193
transform 1 0 5936 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1351_
timestamp 1751534193
transform -1 0 5264 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1352_
timestamp 1751889408
transform -1 0 5264 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1353_
timestamp 1751740063
transform 1 0 3696 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1354_
timestamp 1753182340
transform 1 0 3360 0 -1 23520
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1355_
timestamp 1751534193
transform -1 0 2800 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1356_
timestamp 1753277515
transform 1 0 2688 0 -1 25088
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1357_
timestamp 1751740063
transform 1 0 2576 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1358_
timestamp 1751889408
transform 1 0 2128 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1359_
timestamp 1751740063
transform -1 0 3248 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1360_
timestamp 1751889408
transform -1 0 5264 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1361_
timestamp 1753182340
transform 1 0 3248 0 1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1362_
timestamp 1751534193
transform -1 0 2464 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1363_
timestamp 1751740063
transform 1 0 3248 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1364_
timestamp 1751889408
transform 1 0 2912 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1365_
timestamp 1751889408
transform 1 0 4816 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1366_
timestamp 1751889408
transform 1 0 5264 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1367_
timestamp 1753182340
transform 1 0 4592 0 -1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1368_
timestamp 1751534193
transform -1 0 2464 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _1369_
timestamp 1753172561
transform 1 0 5488 0 1 23520
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1370_
timestamp 1753277515
transform -1 0 7728 0 -1 21952
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1371_
timestamp 1751740063
transform 1 0 5600 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1372_
timestamp 1753182340
transform -1 0 7504 0 -1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1373_
timestamp 1751534193
transform 1 0 7280 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1374_
timestamp 1753371985
transform 1 0 7504 0 -1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1375_
timestamp 1753182340
transform 1 0 6496 0 -1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1376_
timestamp 1751534193
transform 1 0 7728 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1377_
timestamp 1751534193
transform -1 0 5264 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1378_
timestamp 1751740063
transform -1 0 6272 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1379_
timestamp 1751889408
transform -1 0 6048 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1380_
timestamp 1753182340
transform -1 0 5264 0 -1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1381_
timestamp 1751534193
transform -1 0 3136 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1382_
timestamp 1751740063
transform 1 0 3696 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1383_
timestamp 1751889408
transform 1 0 5600 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1384_
timestamp 1751889408
transform -1 0 6496 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1385_
timestamp 1753182340
transform 1 0 4592 0 -1 17248
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1386_
timestamp 1751534193
transform -1 0 2912 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1387_
timestamp 1751740063
transform 1 0 2912 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1388_
timestamp 1751889408
transform 1 0 4480 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1389_
timestamp 1753182340
transform 1 0 4368 0 -1 15680
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1390_
timestamp 1751534193
transform -1 0 2912 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _1391_
timestamp 1753172561
transform 1 0 6272 0 -1 17248
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1392_
timestamp 1751740063
transform -1 0 9632 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1393_
timestamp 1751740063
transform -1 0 8848 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1394_
timestamp 1751889408
transform 1 0 8176 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1395_
timestamp 1751534193
transform 1 0 9408 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1396_
timestamp 1751740063
transform 1 0 5824 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1397_
timestamp 1751889808
transform 1 0 6944 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1398_
timestamp 1753371985
transform 1 0 6608 0 1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1399_
timestamp 1751740063
transform -1 0 6608 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1400_
timestamp 1753182340
transform -1 0 7840 0 -1 14112
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1401_
timestamp 1751534193
transform -1 0 7616 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1402_
timestamp 1753182340
transform 1 0 5488 0 1 12544
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1403_
timestamp 1751534193
transform -1 0 3808 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1404_
timestamp 1751534193
transform 1 0 7840 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1405_
timestamp 1751740063
transform 1 0 8400 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1406_
timestamp 1751889408
transform -1 0 8400 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1407_
timestamp 1753182340
transform 1 0 9408 0 -1 14112
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1408_
timestamp 1751534193
transform -1 0 9184 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1409_
timestamp 1751740063
transform -1 0 12656 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1410_
timestamp 1751889408
transform 1 0 12656 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1411_
timestamp 1753182340
transform 1 0 11648 0 1 12544
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1412_
timestamp 1751534193
transform -1 0 11872 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1413_
timestamp 1751740063
transform -1 0 14896 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1414_
timestamp 1751889408
transform -1 0 14112 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1415_
timestamp 1753182340
transform 1 0 11760 0 1 10976
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1416_
timestamp 1751534193
transform 1 0 12432 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1417_
timestamp 1751740063
transform 1 0 11760 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1418_
timestamp 1751889408
transform 1 0 7392 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1419_
timestamp 1753182340
transform -1 0 10640 0 -1 10976
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1420_
timestamp 1751534193
transform -1 0 8512 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1421_
timestamp 1751534193
transform -1 0 4480 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1422_
timestamp 1751740063
transform -1 0 5264 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1423_
timestamp 1751889408
transform -1 0 5376 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1424_
timestamp 1753182340
transform -1 0 4928 0 1 10976
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1425_
timestamp 1751534193
transform -1 0 2800 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1426_
timestamp 1751740063
transform 1 0 2912 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1427_
timestamp 1751889408
transform -1 0 6160 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1428_
timestamp 1753182340
transform -1 0 4592 0 1 9408
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1429_
timestamp 1751534193
transform -1 0 2800 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1430_
timestamp 1751532043
transform 1 0 4704 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _1431_
timestamp 1753172561
transform 1 0 5488 0 1 10976
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1432_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753441877
transform -1 0 6272 0 -1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1433_
timestamp 1753371985
transform 1 0 4144 0 1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1434_
timestamp 1753371985
transform 1 0 3024 0 1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1435_
timestamp 1751532043
transform -1 0 7168 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1436_
timestamp 1753182340
transform 1 0 5488 0 1 7840
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1437_
timestamp 1751534193
transform 1 0 6496 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1438_
timestamp 1753182340
transform 1 0 5488 0 1 6272
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1439_
timestamp 1751534193
transform -1 0 2912 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1440_
timestamp 1751534193
transform 1 0 5824 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1441_
timestamp 1751740063
transform 1 0 4480 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1442_
timestamp 1751889408
transform 1 0 6048 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1443_
timestamp 1753182340
transform 1 0 4816 0 -1 6272
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1444_
timestamp 1751534193
transform -1 0 4816 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1445_
timestamp 1751534193
transform 1 0 9968 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1446_
timestamp 1751740063
transform 1 0 7392 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1447_
timestamp 1753960525
transform 1 0 6832 0 -1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1448_
timestamp 1751740063
transform -1 0 8960 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1449_
timestamp 1751534193
transform -1 0 10080 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1450_
timestamp 1751532043
transform -1 0 7840 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _1451_
timestamp 1752345181
transform 1 0 7280 0 1 6272
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1452_
timestamp 1753960525
transform 1 0 7952 0 -1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1453_
timestamp 1753371985
transform 1 0 7840 0 -1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _1454_
timestamp 1753891287
transform 1 0 8512 0 1 6272
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1455_
timestamp 1751531619
transform 1 0 9856 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1456_
timestamp 1751740063
transform 1 0 9520 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1457_
timestamp 1753182340
transform 1 0 10304 0 -1 7840
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1458_
timestamp 1751534193
transform 1 0 11088 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1459_
timestamp 1752061876
transform 1 0 10640 0 1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1460_
timestamp 1751534193
transform -1 0 39648 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1461_
timestamp 1751534193
transform -1 0 16576 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1462_
timestamp 1751534193
transform 1 0 32032 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1463_
timestamp 1751534193
transform -1 0 30464 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1464_
timestamp 1752061876
transform -1 0 32032 0 -1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1465_
timestamp 1751532043
transform 1 0 33376 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1466_
timestamp 1751532043
transform -1 0 39536 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _1467_
timestamp 1753172561
transform -1 0 38416 0 1 28224
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1468_
timestamp 1753182340
transform 1 0 33824 0 1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1469_
timestamp 1751889408
transform -1 0 28224 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1470_
timestamp 1751534193
transform 1 0 15232 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1471_
timestamp 1751532043
transform 1 0 41104 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1472_
timestamp 1751534193
transform -1 0 42336 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1473_
timestamp 1751534193
transform -1 0 25760 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1474_
timestamp 1751534193
transform 1 0 23072 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1475_
timestamp 1751740063
transform -1 0 24528 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1476_
timestamp 1751534193
transform -1 0 20944 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1477_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753868718
transform 1 0 15568 0 -1 21952
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1478_
timestamp 1751534193
transform -1 0 16576 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1479_
timestamp 1751534193
transform -1 0 21840 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1480_
timestamp 1753868718
transform -1 0 13104 0 1 21952
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1481_
timestamp 1751534193
transform -1 0 10304 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1482_
timestamp 1751534193
transform -1 0 14672 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1483_
timestamp 1753868718
transform -1 0 14560 0 1 21952
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1484_
timestamp 1751534193
transform 1 0 13328 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1485_
timestamp 1751534193
transform -1 0 14000 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1486_
timestamp 1753868718
transform -1 0 12768 0 -1 23520
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1487_
timestamp 1751534193
transform -1 0 10976 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1488_
timestamp 1751534193
transform -1 0 38304 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1489_
timestamp 1751534193
transform 1 0 29120 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1490_
timestamp 1753868718
transform -1 0 22400 0 1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1491_
timestamp 1751534193
transform 1 0 21392 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1492_
timestamp 1752061876
transform 1 0 30912 0 1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1493_
timestamp 1751889408
transform -1 0 28448 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1494_
timestamp 1751534193
transform -1 0 9184 0 -1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1495_
timestamp 1751534193
transform -1 0 44352 0 1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1496_
timestamp 1751534193
transform -1 0 33600 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1497_
timestamp 1751740063
transform -1 0 10304 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1498_
timestamp 1753868718
transform -1 0 11200 0 1 32928
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1499_
timestamp 1751534193
transform -1 0 9184 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1500_
timestamp 1753868718
transform -1 0 10640 0 -1 36064
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1501_
timestamp 1751534193
transform -1 0 9184 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1502_
timestamp 1753868718
transform -1 0 10640 0 -1 34496
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1503_
timestamp 1751534193
transform -1 0 6272 0 1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1504_
timestamp 1753868718
transform -1 0 11872 0 -1 34496
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1505_
timestamp 1751534193
transform -1 0 6720 0 1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1506_
timestamp 1751534193
transform 1 0 24416 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1507_
timestamp 1751534193
transform 1 0 37520 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1508_
timestamp 1751740063
transform -1 0 39760 0 -1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1509_
timestamp 1751889408
transform -1 0 39424 0 1 3136
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1510_
timestamp 1753182340
transform 1 0 37296 0 1 4704
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1511_
timestamp 1751534193
transform 1 0 39760 0 -1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1512_
timestamp 1751532043
transform -1 0 37408 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1513_
timestamp 1753277515
transform 1 0 37296 0 -1 7840
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1514_
timestamp 1751534193
transform -1 0 38304 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1515_
timestamp 1751534193
transform 1 0 42112 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1516_
timestamp 1751889808
transform 1 0 39536 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1517_
timestamp 1751531619
transform -1 0 40208 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1518_
timestamp 1753371985
transform 1 0 38304 0 -1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1519_
timestamp 1751889408
transform 1 0 37408 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1520_
timestamp 1753960525
transform 1 0 37632 0 1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1521_
timestamp 1751740063
transform 1 0 37184 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1522_
timestamp 1751889408
transform 1 0 38752 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1523_
timestamp 1753182340
transform 1 0 38864 0 1 9408
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1524_
timestamp 1751534193
transform -1 0 37632 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1525_
timestamp 1751740063
transform -1 0 41552 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1526_
timestamp 1751889408
transform 1 0 38304 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1527_
timestamp 1753182340
transform -1 0 39872 0 -1 10976
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1528_
timestamp 1751534193
transform 1 0 39760 0 -1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1529_
timestamp 1751889808
transform 1 0 38976 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _1530_
timestamp 1753172561
transform -1 0 38864 0 1 9408
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1531_
timestamp 1751889408
transform 1 0 35728 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1532_
timestamp 1751889408
transform -1 0 36624 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1533_
timestamp 1751534193
transform 1 0 35952 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1534_
timestamp 1751532043
transform 1 0 35280 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1535_
timestamp 1751740063
transform 1 0 35728 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1536_
timestamp 1751534193
transform 1 0 24192 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1537_
timestamp 1753441877
transform -1 0 35728 0 1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1538_
timestamp 1751740063
transform 1 0 34496 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1539_
timestamp 1751889408
transform -1 0 35168 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1540_
timestamp 1751889808
transform 1 0 35168 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1541_
timestamp 1751531619
transform -1 0 36736 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1542_
timestamp 1751740063
transform 1 0 34496 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1543_
timestamp 1751534193
transform -1 0 24864 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1544_
timestamp 1751534193
transform 1 0 25424 0 -1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1545_
timestamp 1751534193
transform 1 0 28896 0 -1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1546_
timestamp 1751740063
transform 1 0 33712 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1547_
timestamp 1751889408
transform -1 0 33712 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1548_
timestamp 1753182340
transform 1 0 31472 0 -1 6272
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1549_
timestamp 1751534193
transform -1 0 31472 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1550_
timestamp 1751534193
transform -1 0 35728 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1551_
timestamp 1751889408
transform -1 0 32928 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1552_
timestamp 1751534193
transform -1 0 31920 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1553_
timestamp 1751534193
transform 1 0 22400 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1554_
timestamp 1751534193
transform 1 0 22512 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1555_
timestamp 1751889408
transform 1 0 45920 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1556_
timestamp 1751534193
transform -1 0 43680 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1557_
timestamp 1751534193
transform 1 0 48272 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1558_
timestamp 1751889808
transform 1 0 42224 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1559_
timestamp 1752061876
transform 1 0 43232 0 -1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1560_
timestamp 1751534193
transform 1 0 48608 0 -1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1561_
timestamp 1751889408
transform -1 0 43904 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1562_
timestamp 1753960525
transform -1 0 41216 0 1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1563_
timestamp 1751534193
transform 1 0 41888 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1564_
timestamp 1751740063
transform -1 0 45136 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1565_
timestamp 1753868718
transform -1 0 45024 0 -1 9408
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1566_
timestamp 1753960525
transform -1 0 40432 0 -1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1567_
timestamp 1751534193
transform 1 0 39872 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1568_
timestamp 1751534193
transform 1 0 48608 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1569_
timestamp 1751534193
transform -1 0 47040 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1570_
timestamp 1753868718
transform -1 0 43904 0 1 6272
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1571_
timestamp 1751534193
transform -1 0 43120 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1572_
timestamp 1753868718
transform -1 0 45136 0 -1 6272
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1573_
timestamp 1751534193
transform -1 0 42672 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1574_
timestamp 1753868718
transform -1 0 44800 0 1 3136
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1575_
timestamp 1751534193
transform 1 0 47936 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1576_
timestamp 1751534193
transform 1 0 43344 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1577_
timestamp 1751534193
transform 1 0 48496 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1578_
timestamp 1753868718
transform -1 0 45920 0 1 6272
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1579_
timestamp 1751534193
transform 1 0 48608 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1580_
timestamp 1753868718
transform -1 0 46368 0 1 3136
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1581_
timestamp 1751534193
transform 1 0 48608 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1582_
timestamp 1753868718
transform 1 0 47712 0 1 4704
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1583_
timestamp 1751534193
transform 1 0 48608 0 -1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1584_
timestamp 1753868718
transform -1 0 45584 0 -1 7840
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1585_
timestamp 1751534193
transform 1 0 47376 0 -1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1586_
timestamp 1753868718
transform 1 0 45024 0 1 7840
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1587_
timestamp 1751534193
transform 1 0 48608 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1588_
timestamp 1751740063
transform -1 0 32032 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1589_
timestamp 1751889408
transform -1 0 32368 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1590_
timestamp 1753182340
transform -1 0 31584 0 -1 7840
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1591_
timestamp 1751534193
transform -1 0 30912 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1592_
timestamp 1751740063
transform 1 0 29680 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1593_
timestamp 1751889408
transform 1 0 30464 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1594_
timestamp 1753182340
transform 1 0 30128 0 -1 6272
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1595_
timestamp 1751534193
transform -1 0 29680 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1596_
timestamp 1751740063
transform 1 0 30016 0 1 3136
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1597_
timestamp 1751889408
transform -1 0 28784 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1598_
timestamp 1753182340
transform -1 0 30016 0 1 3136
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1599_
timestamp 1751534193
transform -1 0 28000 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1600_
timestamp 1751534193
transform -1 0 24192 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1601_
timestamp 1751740063
transform 1 0 20160 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1602_
timestamp 1751889408
transform -1 0 18032 0 -1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1603_
timestamp 1753182340
transform -1 0 19264 0 -1 4704
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1604_
timestamp 1751534193
transform -1 0 15120 0 -1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1605_
timestamp 1751740063
transform 1 0 15456 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1606_
timestamp 1751889408
transform 1 0 16240 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1607_
timestamp 1753182340
transform 1 0 15792 0 -1 4704
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1608_
timestamp 1751534193
transform -1 0 15456 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1609_
timestamp 1751740063
transform -1 0 18032 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1610_
timestamp 1751889408
transform 1 0 17584 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1611_
timestamp 1753182340
transform 1 0 16352 0 1 6272
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1612_
timestamp 1751534193
transform 1 0 17248 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1613_
timestamp 1751740063
transform -1 0 21392 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1614_
timestamp 1751889408
transform -1 0 20160 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1615_
timestamp 1753182340
transform 1 0 18816 0 1 6272
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1616_
timestamp 1751534193
transform 1 0 20160 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1617_
timestamp 1751889408
transform 1 0 20048 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1618_
timestamp 1751534193
transform 1 0 21168 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1619_
timestamp 1751534193
transform 1 0 27216 0 -1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1620_
timestamp 1751740063
transform -1 0 32256 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1621_
timestamp 1751889408
transform -1 0 33712 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1622_
timestamp 1753182340
transform 1 0 30912 0 -1 15680
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1623_
timestamp 1751534193
transform 1 0 32256 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1624_
timestamp 1751740063
transform 1 0 29008 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1625_
timestamp 1751889408
transform 1 0 30352 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1626_
timestamp 1753182340
transform 1 0 29120 0 1 14112
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1627_
timestamp 1751534193
transform -1 0 29680 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1628_
timestamp 1751740063
transform -1 0 31024 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1629_
timestamp 1751889408
transform 1 0 31472 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1630_
timestamp 1753182340
transform -1 0 30240 0 1 12544
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1631_
timestamp 1751534193
transform -1 0 28336 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1632_
timestamp 1751740063
transform 1 0 27888 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1633_
timestamp 1751889408
transform 1 0 28560 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1634_
timestamp 1753182340
transform -1 0 30240 0 1 10976
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1635_
timestamp 1751534193
transform -1 0 28224 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1636_
timestamp 1751534193
transform 1 0 25088 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1637_
timestamp 1751740063
transform -1 0 28784 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1638_
timestamp 1751889408
transform 1 0 29008 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1639_
timestamp 1753182340
transform -1 0 28336 0 1 7840
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1640_
timestamp 1751534193
transform -1 0 27664 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1641_
timestamp 1751740063
transform -1 0 28112 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1642_
timestamp 1751889408
transform 1 0 28112 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1643_
timestamp 1753182340
transform -1 0 27328 0 1 6272
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1644_
timestamp 1751534193
transform -1 0 26656 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1645_
timestamp 1751740063
transform 1 0 24864 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1646_
timestamp 1751889408
transform 1 0 24976 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1647_
timestamp 1753182340
transform -1 0 24864 0 1 6272
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1648_
timestamp 1751534193
transform -1 0 23520 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1649_
timestamp 1751889408
transform -1 0 24752 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1650_
timestamp 1751534193
transform 1 0 24192 0 -1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1651_
timestamp 1751740063
transform 1 0 32032 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1652_
timestamp 1751889408
transform -1 0 27664 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1653_
timestamp 1751534193
transform -1 0 18816 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1654_
timestamp 1751534193
transform -1 0 30800 0 -1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1655_
timestamp 1751740063
transform -1 0 21504 0 -1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1656_
timestamp 1751534193
transform -1 0 19936 0 -1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1657_
timestamp 1753868718
transform -1 0 15456 0 1 34496
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1658_
timestamp 1751534193
transform 1 0 14560 0 1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1659_
timestamp 1753868718
transform 1 0 16240 0 1 36064
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1660_
timestamp 1751534193
transform 1 0 18816 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1661_
timestamp 1753868718
transform -1 0 13104 0 1 36064
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1662_
timestamp 1751534193
transform -1 0 11872 0 1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1663_
timestamp 1753868718
transform -1 0 12992 0 -1 36064
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1664_
timestamp 1751534193
transform 1 0 11872 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1665_
timestamp 1751534193
transform 1 0 18144 0 1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1666_
timestamp 1751534193
transform -1 0 19488 0 1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1667_
timestamp 1753868718
transform -1 0 20720 0 1 39200
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1668_
timestamp 1751534193
transform -1 0 20048 0 1 40768
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1669_
timestamp 1751534193
transform -1 0 37520 0 1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1670_
timestamp 1753868718
transform -1 0 20720 0 -1 43904
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1671_
timestamp 1751534193
transform -1 0 20048 0 -1 47040
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1672_
timestamp 1751534193
transform -1 0 38640 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1673_
timestamp 1753868718
transform -1 0 20720 0 1 43904
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1674_
timestamp 1751534193
transform -1 0 19488 0 1 43904
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1675_
timestamp 1751534193
transform -1 0 40320 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1676_
timestamp 1753868718
transform -1 0 20832 0 -1 42336
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1677_
timestamp 1751534193
transform -1 0 19488 0 -1 43904
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1678_
timestamp 1751889408
transform 1 0 31136 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1679_
timestamp 1753182340
transform 1 0 33824 0 -1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1680_
timestamp 1751889408
transform -1 0 30912 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1681_
timestamp 1751534193
transform -1 0 15680 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1682_
timestamp 1751740063
transform -1 0 15008 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1683_
timestamp 1753868718
transform 1 0 13552 0 -1 26656
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1684_
timestamp 1751534193
transform 1 0 14784 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1685_
timestamp 1753868718
transform -1 0 13104 0 1 23520
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1686_
timestamp 1751534193
transform 1 0 12208 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1687_
timestamp 1753868718
transform -1 0 12544 0 1 25088
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1688_
timestamp 1751534193
transform -1 0 10080 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1689_
timestamp 1753868718
transform -1 0 11200 0 -1 25088
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1690_
timestamp 1751534193
transform -1 0 9184 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1691_
timestamp 1751534193
transform -1 0 37520 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1692_
timestamp 1751889408
transform -1 0 28112 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1693_
timestamp 1751534193
transform 1 0 25312 0 -1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1694_
timestamp 1751740063
transform -1 0 24976 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1695_
timestamp 1751534193
transform 1 0 24192 0 -1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1696_
timestamp 1753868718
transform 1 0 25984 0 -1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1697_
timestamp 1751534193
transform 1 0 26768 0 -1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1698_
timestamp 1751534193
transform -1 0 37520 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1699_
timestamp 1753868718
transform -1 0 26320 0 -1 31360
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1700_
timestamp 1751534193
transform -1 0 24864 0 -1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1701_
timestamp 1751534193
transform -1 0 35392 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1702_
timestamp 1753868718
transform 1 0 25088 0 -1 26656
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1703_
timestamp 1751534193
transform 1 0 26992 0 1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1704_
timestamp 1751534193
transform 1 0 35392 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1705_
timestamp 1753868718
transform -1 0 26768 0 1 28224
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1706_
timestamp 1751534193
transform 1 0 26768 0 1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1707_
timestamp 1751534193
transform -1 0 25760 0 -1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1708_
timestamp 1751534193
transform -1 0 24192 0 -1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1709_
timestamp 1753868718
transform -1 0 23968 0 1 31360
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1710_
timestamp 1751534193
transform -1 0 22176 0 1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1711_
timestamp 1753868718
transform -1 0 23408 0 1 32928
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1712_
timestamp 1751534193
transform 1 0 22736 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1713_
timestamp 1753868718
transform 1 0 24304 0 1 34496
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1714_
timestamp 1751534193
transform 1 0 25088 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1715_
timestamp 1753868718
transform 1 0 24976 0 1 31360
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1716_
timestamp 1751534193
transform 1 0 26208 0 1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1717_
timestamp 1751534193
transform -1 0 41440 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1718_
timestamp 1751740063
transform 1 0 46144 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1719_
timestamp 1751889408
transform 1 0 47712 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1720_
timestamp 1753182340
transform 1 0 46928 0 -1 12544
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1721_
timestamp 1751534193
transform 1 0 48608 0 -1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1722_
timestamp 1751740063
transform -1 0 48272 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1723_
timestamp 1751889408
transform 1 0 48608 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1724_
timestamp 1753182340
transform 1 0 47040 0 -1 14112
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1725_
timestamp 1751534193
transform 1 0 47712 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1726_
timestamp 1753277515
transform -1 0 46256 0 1 14112
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1727_
timestamp 1751740063
transform -1 0 44464 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1728_
timestamp 1753371985
transform 1 0 44688 0 1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1729_
timestamp 1751740063
transform 1 0 41440 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1730_
timestamp 1751740063
transform -1 0 32368 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1731_
timestamp 1751889408
transform 1 0 32928 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1732_
timestamp 1753182340
transform 1 0 30352 0 1 10976
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1733_
timestamp 1751534193
transform -1 0 30912 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1734_
timestamp 1751534193
transform -1 0 27776 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1735_
timestamp 1751534193
transform -1 0 34608 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1736_
timestamp 1751740063
transform -1 0 34160 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1737_
timestamp 1751889408
transform 1 0 34160 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1738_
timestamp 1753182340
transform 1 0 34048 0 1 12544
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1739_
timestamp 1751534193
transform -1 0 33040 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1740_
timestamp 1751740063
transform 1 0 33600 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1741_
timestamp 1751889408
transform 1 0 33936 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1742_
timestamp 1753182340
transform 1 0 33488 0 -1 14112
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1743_
timestamp 1751534193
transform -1 0 32704 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1744_
timestamp 1751740063
transform -1 0 37632 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1745_
timestamp 1751889408
transform -1 0 35504 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1746_
timestamp 1753182340
transform 1 0 35056 0 1 14112
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1747_
timestamp 1751534193
transform 1 0 37632 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1748_
timestamp 1751740063
transform -1 0 36288 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1749_
timestamp 1751889408
transform 1 0 36288 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1750_
timestamp 1753182340
transform 1 0 34944 0 1 15680
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1751_
timestamp 1751534193
transform 1 0 35616 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1752_
timestamp 1751534193
transform 1 0 37520 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1753_
timestamp 1751740063
transform -1 0 39088 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1754_
timestamp 1751889408
transform 1 0 39088 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1755_
timestamp 1753182340
transform 1 0 38192 0 -1 15680
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1756_
timestamp 1751534193
transform 1 0 39872 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1757_
timestamp 1751740063
transform -1 0 39872 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1758_
timestamp 1751889408
transform 1 0 39424 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1759_
timestamp 1753182340
transform -1 0 39536 0 1 14112
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1760_
timestamp 1751534193
transform 1 0 39872 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1761_
timestamp 1751534193
transform 1 0 39536 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1762_
timestamp 1751889408
transform -1 0 39088 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1763_
timestamp 1751534193
transform -1 0 27104 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1764_
timestamp 1751532043
transform 1 0 35168 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1765_
timestamp 1753182340
transform -1 0 35168 0 1 28224
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1766_
timestamp 1751889408
transform -1 0 29120 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1767_
timestamp 1751740063
transform 1 0 27888 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1768_
timestamp 1753868718
transform -1 0 29120 0 -1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1769_
timestamp 1751534193
transform -1 0 26432 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1770_
timestamp 1753868718
transform 1 0 29008 0 1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1771_
timestamp 1751534193
transform -1 0 28112 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1772_
timestamp 1753182340
transform 1 0 35056 0 1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1773_
timestamp 1751889408
transform 1 0 33040 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1774_
timestamp 1751534193
transform 1 0 35392 0 1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1775_
timestamp 1751740063
transform 1 0 34496 0 1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1776_
timestamp 1751534193
transform -1 0 35280 0 -1 40768
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1777_
timestamp 1753868718
transform 1 0 36624 0 -1 39200
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1778_
timestamp 1751534193
transform 1 0 37968 0 -1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1779_
timestamp 1753868718
transform 1 0 36288 0 -1 40768
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1780_
timestamp 1751534193
transform 1 0 39648 0 -1 42336
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1781_
timestamp 1753868718
transform 1 0 35392 0 1 37632
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1782_
timestamp 1751534193
transform 1 0 36848 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1783_
timestamp 1753868718
transform 1 0 36848 0 1 39200
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1784_
timestamp 1751534193
transform 1 0 38752 0 1 42336
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1785_
timestamp 1751534193
transform -1 0 37632 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1786_
timestamp 1751534193
transform 1 0 38080 0 1 42336
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1787_
timestamp 1751534193
transform 1 0 40096 0 1 40768
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1788_
timestamp 1753868718
transform -1 0 38528 0 -1 45472
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1789_
timestamp 1751534193
transform 1 0 37296 0 1 47040
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1790_
timestamp 1753868718
transform 1 0 36064 0 -1 45472
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1791_
timestamp 1751534193
transform 1 0 38528 0 -1 45472
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1792_
timestamp 1753868718
transform 1 0 36848 0 1 42336
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1793_
timestamp 1751534193
transform 1 0 37632 0 1 43904
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1794_
timestamp 1753868718
transform -1 0 36624 0 -1 42336
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1795_
timestamp 1751534193
transform 1 0 35952 0 1 42336
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1796_
timestamp 1751889408
transform -1 0 29232 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1797_
timestamp 1751534193
transform -1 0 29120 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1798_
timestamp 1751740063
transform 1 0 28448 0 -1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1799_
timestamp 1751534193
transform 1 0 29232 0 -1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1800_
timestamp 1753868718
transform 1 0 28672 0 -1 34496
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1801_
timestamp 1751534193
transform 1 0 29904 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1802_
timestamp 1753868718
transform 1 0 29120 0 -1 36064
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1803_
timestamp 1751534193
transform 1 0 30128 0 -1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1804_
timestamp 1753868718
transform -1 0 27888 0 -1 36064
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1805_
timestamp 1751534193
transform 1 0 26880 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1806_
timestamp 1753868718
transform -1 0 28560 0 1 36064
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1807_
timestamp 1751534193
transform -1 0 26208 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1808_
timestamp 1751534193
transform 1 0 29568 0 -1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1809_
timestamp 1751534193
transform 1 0 28896 0 -1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1810_
timestamp 1753868718
transform 1 0 32928 0 -1 40768
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1811_
timestamp 1751534193
transform 1 0 33712 0 -1 42336
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1812_
timestamp 1753868718
transform 1 0 31472 0 -1 39200
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1813_
timestamp 1751534193
transform 1 0 32928 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1814_
timestamp 1753868718
transform -1 0 29456 0 -1 43904
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1815_
timestamp 1751534193
transform -1 0 27776 0 1 45472
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1816_
timestamp 1753868718
transform -1 0 28448 0 1 42336
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1817_
timestamp 1751534193
transform -1 0 25872 0 1 42336
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1818_
timestamp 1751531619
transform -1 0 35616 0 1 3136
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1819_
timestamp 1751740063
transform -1 0 43120 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _1820_
timestamp 1751914308
transform -1 0 43232 0 -1 10976
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1821_
timestamp 1751889408
transform -1 0 42336 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1822_
timestamp 1751534193
transform -1 0 41888 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1823_
timestamp 1751531619
transform -1 0 22400 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1824_
timestamp 1751532043
transform 1 0 20720 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1825_
timestamp 1751534193
transform -1 0 38976 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1826_
timestamp 1751889408
transform -1 0 33712 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1827_
timestamp 1751534193
transform -1 0 33376 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1828_
timestamp 1751740063
transform 1 0 33488 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1829_
timestamp 1751534193
transform -1 0 32704 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1830_
timestamp 1753868718
transform -1 0 32704 0 -1 23520
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1831_
timestamp 1751534193
transform 1 0 32928 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1832_
timestamp 1753868718
transform -1 0 26768 0 -1 23520
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1833_
timestamp 1751534193
transform -1 0 24864 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1834_
timestamp 1753868718
transform 1 0 25872 0 1 23520
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1835_
timestamp 1751534193
transform -1 0 26992 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1836_
timestamp 1753868718
transform -1 0 30352 0 -1 23520
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1837_
timestamp 1751534193
transform -1 0 29120 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1838_
timestamp 1753868718
transform -1 0 35168 0 1 21952
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1839_
timestamp 1751534193
transform 1 0 33936 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1840_
timestamp 1753868718
transform 1 0 35168 0 1 21952
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1841_
timestamp 1751534193
transform 1 0 36848 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1842_
timestamp 1751889408
transform 1 0 34944 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1843_
timestamp 1751534193
transform -1 0 39200 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1844_
timestamp 1752061876
transform 1 0 47264 0 -1 29792
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1845_
timestamp 1751532043
transform 1 0 44688 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1846_
timestamp 1751532043
transform -1 0 46368 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1847_
timestamp 1753960525
transform 1 0 44800 0 -1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1848_
timestamp 1751889408
transform 1 0 45696 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1849_
timestamp 1751889408
transform 1 0 48608 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1850_
timestamp 1751740063
transform 1 0 45024 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1851_
timestamp 1751889808
transform 1 0 42448 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1852_
timestamp 1751534193
transform -1 0 46816 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1853_
timestamp 1753182340
transform -1 0 47040 0 -1 21952
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1854_
timestamp 1751534193
transform -1 0 46480 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1855_
timestamp 1751740063
transform -1 0 47264 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1856_
timestamp 1751889408
transform -1 0 49392 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1857_
timestamp 1753182340
transform 1 0 47824 0 1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1858_
timestamp 1751534193
transform -1 0 47488 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1859_
timestamp 1751740063
transform -1 0 48272 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1860_
timestamp 1751889408
transform 1 0 48048 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1861_
timestamp 1753182340
transform 1 0 46816 0 1 23520
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1862_
timestamp 1751534193
transform 1 0 48608 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1863_
timestamp 1751889808
transform 1 0 47712 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1864_
timestamp 1753371985
transform -1 0 48272 0 -1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1865_
timestamp 1751889408
transform 1 0 48608 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1866_
timestamp 1751534193
transform -1 0 49280 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1867_
timestamp 1751889408
transform 1 0 48608 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _1868_
timestamp 1753172561
transform 1 0 46816 0 -1 25088
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1869_
timestamp 1753371985
transform 1 0 45248 0 1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1870_
timestamp 1751532043
transform -1 0 44464 0 1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1871_
timestamp 1751532043
transform 1 0 46256 0 -1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1872_
timestamp 1751532043
transform 1 0 44688 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_2  _1873_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753579406
transform -1 0 46256 0 1 40768
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1874_
timestamp 1751532043
transform -1 0 45136 0 1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1875_
timestamp 1751532043
transform -1 0 42784 0 -1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1876_
timestamp 1753868718
transform 1 0 44464 0 -1 43904
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1877_
timestamp 1751532043
transform 1 0 47936 0 1 47040
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1878_
timestamp 1751531619
transform -1 0 45472 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1879_
timestamp 1751532043
transform 1 0 41328 0 -1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1880_
timestamp 1751532043
transform 1 0 41776 0 -1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1881_
timestamp 1753868718
transform 1 0 42112 0 1 40768
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1882_
timestamp 1751889808
transform 1 0 42336 0 -1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1883_
timestamp 1753277515
transform 1 0 40768 0 -1 42336
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1884_
timestamp 1753277515
transform 1 0 40768 0 1 42336
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1885_
timestamp 1751889408
transform 1 0 42336 0 1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1886_
timestamp 1751532043
transform 1 0 40768 0 -1 43904
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1887_
timestamp 1751534193
transform -1 0 40544 0 -1 43904
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _1888_
timestamp 1752061876
transform 1 0 39648 0 1 42336
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1889_
timestamp 1753272495
transform 1 0 41216 0 -1 43904
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1890_
timestamp 1753960525
transform 1 0 43232 0 1 42336
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1891_
timestamp 1751532043
transform 1 0 42784 0 1 47040
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1892_
timestamp 1751532043
transform 1 0 42896 0 -1 43904
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1893_
timestamp 1753868718
transform 1 0 45584 0 -1 45472
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1894_
timestamp 1753371985
transform 1 0 43344 0 -1 43904
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1895_
timestamp 1751889808
transform 1 0 45696 0 -1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1896_
timestamp 1753868718
transform 1 0 45024 0 -1 40768
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1897_
timestamp 1751532043
transform 1 0 44912 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1898_
timestamp 1751532043
transform -1 0 45472 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1899_
timestamp 1751534193
transform -1 0 49280 0 1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1900_
timestamp 1751532043
transform 1 0 45920 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1901_
timestamp 1751532043
transform 1 0 42896 0 -1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1902_
timestamp 1751531619
transform -1 0 42560 0 -1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1903_
timestamp 1751532043
transform -1 0 40544 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1904_
timestamp 1751532043
transform 1 0 41776 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _1905_
timestamp 1751905124
transform 1 0 36848 0 1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1906_
timestamp 1753272495
transform 1 0 38304 0 -1 34496
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1907_
timestamp 1753272495
transform 1 0 40432 0 1 32928
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1908_
timestamp 1751532043
transform 1 0 42448 0 -1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1909_
timestamp 1751532043
transform -1 0 44128 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1910_
timestamp 1753868718
transform 1 0 42448 0 1 32928
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1911_
timestamp 1753441877
transform 1 0 42560 0 -1 32928
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1912_
timestamp 1751532043
transform -1 0 46368 0 1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1913_
timestamp 1751532043
transform 1 0 47712 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_2  _1914_
timestamp 1753579406
transform -1 0 45584 0 -1 32928
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1915_
timestamp 1753868718
transform -1 0 45920 0 1 32928
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _1916_
timestamp 1753272495
transform 1 0 44464 0 -1 34496
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1917_
timestamp 1753441877
transform 1 0 45136 0 -1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1918_
timestamp 1753182340
transform -1 0 46032 0 1 42336
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _1919_
timestamp 1753172561
transform -1 0 44688 0 -1 42336
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1920_
timestamp 1751532043
transform 1 0 45136 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1921_
timestamp 1751532043
transform -1 0 42672 0 -1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1922_
timestamp 1751532043
transform -1 0 45136 0 1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1923_
timestamp 1753868718
transform -1 0 45024 0 -1 40768
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _1924_
timestamp 1753371985
transform 1 0 42672 0 -1 40768
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _1925_
timestamp 1753172561
transform -1 0 46816 0 1 39200
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1926_
timestamp 1751532043
transform -1 0 42000 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1927_
timestamp 1751740063
transform 1 0 40768 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1928_
timestamp 1751532043
transform 1 0 40992 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_4  _1929_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753869255
transform -1 0 42560 0 1 20384
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1930_
timestamp 1751534193
transform 1 0 32032 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1931_
timestamp 1751740063
transform 1 0 43344 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1932_
timestamp 1751740063
transform 1 0 43568 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _1933_
timestamp 1751905124
transform 1 0 42784 0 -1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1934_
timestamp 1753441877
transform 1 0 43904 0 -1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1935_
timestamp 1751534193
transform -1 0 33264 0 1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1936_
timestamp 1751531619
transform -1 0 33712 0 -1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _1937_
timestamp 1753441877
transform 1 0 46816 0 1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1938_
timestamp 1751740063
transform -1 0 42896 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1939_
timestamp 1751531619
transform 1 0 47600 0 -1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1940_
timestamp 1751534193
transform 1 0 48608 0 -1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1941_
timestamp 1751531619
transform 1 0 46928 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _1942_
timestamp 1753868718
transform 1 0 46928 0 -1 39200
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1943_
timestamp 1751534193
transform 1 0 48608 0 -1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1944_
timestamp 1751534193
transform -1 0 46368 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1945_
timestamp 1751534193
transform 1 0 32032 0 -1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1946_
timestamp 1753277515
transform 1 0 33152 0 -1 37632
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _1947_
timestamp 1751889808
transform -1 0 35392 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1948_
timestamp 1751534193
transform 1 0 35952 0 -1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1949_
timestamp 1751534193
transform -1 0 46928 0 -1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1950_
timestamp 1751534193
transform -1 0 32032 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1951_
timestamp 1751534193
transform 1 0 37296 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1952_
timestamp 1753960525
transform 1 0 33264 0 -1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _1953_
timestamp 1753172561
transform -1 0 34608 0 1 34496
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1954_
timestamp 1751531619
transform 1 0 35056 0 1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1955_
timestamp 1751740063
transform -1 0 36624 0 1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1956_
timestamp 1751534193
transform 1 0 48608 0 -1 42336
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _1957_
timestamp 1751532043
transform 1 0 42560 0 1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1958_
timestamp 1751740063
transform -1 0 42448 0 -1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1959_
timestamp 1751889408
transform -1 0 41664 0 -1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1960_
timestamp 1753182340
transform 1 0 40768 0 -1 36064
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1961_
timestamp 1751534193
transform -1 0 39424 0 1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1962_
timestamp 1751740063
transform 1 0 39760 0 -1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1963_
timestamp 1753182340
transform -1 0 42560 0 1 34496
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1964_
timestamp 1751534193
transform 1 0 43232 0 1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1965_
timestamp 1753182340
transform 1 0 40768 0 -1 37632
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1966_
timestamp 1751534193
transform 1 0 42000 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1967_
timestamp 1751534193
transform 1 0 43792 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1968_
timestamp 1751889408
transform 1 0 45584 0 1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1969_
timestamp 1751740063
transform -1 0 49392 0 -1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1970_
timestamp 1753182340
transform 1 0 46368 0 -1 37632
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1971_
timestamp 1751534193
transform 1 0 47600 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1972_
timestamp 1753277515
transform 1 0 46032 0 -1 34496
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1973_
timestamp 1751740063
transform -1 0 48048 0 -1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1974_
timestamp 1753960525
transform -1 0 45808 0 1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _1975_
timestamp 1753172561
transform 1 0 45696 0 -1 36064
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1976_
timestamp 1751531619
transform 1 0 44688 0 1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1977_
timestamp 1751740063
transform -1 0 44352 0 1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1978_
timestamp 1751889408
transform 1 0 44688 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1979_
timestamp 1751740063
transform -1 0 44352 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1980_
timestamp 1753182340
transform -1 0 45136 0 -1 39200
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1981_
timestamp 1751534193
transform 1 0 48608 0 -1 43904
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1982_
timestamp 1753277515
transform -1 0 43568 0 1 37632
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1983_
timestamp 1751740063
transform 1 0 41104 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1984_
timestamp 1751534193
transform -1 0 46368 0 -1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1985_
timestamp 1751534193
transform 1 0 43120 0 1 43904
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1986_
timestamp 1753182340
transform 1 0 42672 0 1 39200
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1987_
timestamp 1753277515
transform 1 0 42560 0 1 45472
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1988_
timestamp 1751740063
transform -1 0 47040 0 1 47040
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1989_
timestamp 1751889408
transform -1 0 43120 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _1990_
timestamp 1753277515
transform 1 0 40768 0 -1 45472
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1991_
timestamp 1751740063
transform -1 0 42112 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _1992_
timestamp 1753960525
transform -1 0 42112 0 -1 47040
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _1993_
timestamp 1753172561
transform 1 0 40992 0 1 45472
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _1994_
timestamp 1751531619
transform -1 0 40992 0 1 45472
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1995_
timestamp 1751740063
transform 1 0 39760 0 -1 47040
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _1996_
timestamp 1751889408
transform -1 0 46256 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _1997_
timestamp 1751740063
transform -1 0 47040 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _1998_
timestamp 1753182340
transform 1 0 45136 0 1 45472
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1999_
timestamp 1751534193
transform 1 0 48608 0 -1 47040
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2000_
timestamp 1751740063
transform 1 0 47152 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2001_
timestamp 1751889408
transform 1 0 48608 0 -1 45472
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2002_
timestamp 1753182340
transform 1 0 47152 0 -1 45472
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2003_
timestamp 1751534193
transform -1 0 44464 0 1 43904
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2004_
timestamp 1753277515
transform 1 0 46816 0 -1 40768
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2005_
timestamp 1751740063
transform 1 0 47376 0 -1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2006_
timestamp 1753371985
transform 1 0 47936 0 1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2007_
timestamp 1751740063
transform -1 0 49392 0 -1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2008_
timestamp 1751532043
transform 1 0 44912 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2009_
timestamp 1751532043
transform 1 0 44016 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2010_
timestamp 1753277515
transform 1 0 42448 0 1 25088
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2011_
timestamp 1753441877
transform 1 0 44128 0 -1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2012_
timestamp 1753441877
transform 1 0 44688 0 1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2013_
timestamp 1753277515
transform 1 0 44688 0 1 21952
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _2014_
timestamp 1751914308
transform -1 0 44912 0 -1 23520
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2015_
timestamp 1751534193
transform -1 0 43680 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2016_
timestamp 1751532043
transform 1 0 26208 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _2017_
timestamp 1752061876
transform 1 0 22400 0 -1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2018_
timestamp 1751534193
transform -1 0 23184 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2019_
timestamp 1751534193
transform -1 0 22512 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2020_
timestamp 1751534193
transform 1 0 22736 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2021_
timestamp 1751532043
transform -1 0 24864 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _2022_
timestamp 1751905124
transform -1 0 22400 0 -1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2023_
timestamp 1751534193
transform 1 0 23072 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2024_
timestamp 1753441877
transform 1 0 27104 0 -1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2025_
timestamp 1753371985
transform 1 0 25984 0 -1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2026_
timestamp 1751532043
transform 1 0 25312 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2027_
timestamp 1753441877
transform -1 0 27104 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2028_
timestamp 1753371985
transform 1 0 24864 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2029_
timestamp 1751532043
transform 1 0 24304 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2030_
timestamp 1751531619
transform 1 0 22736 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2031_
timestamp 1751534193
transform 1 0 23744 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2032_
timestamp 1751534193
transform 1 0 24192 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2033_
timestamp 1753371985
transform 1 0 23744 0 -1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2034_
timestamp 1751889408
transform 1 0 24192 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2035_
timestamp 1751534193
transform 1 0 25088 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2036_
timestamp 1751532043
transform -1 0 20944 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2037_
timestamp 1751534193
transform 1 0 18368 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2038_
timestamp 1753441877
transform -1 0 22400 0 1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2039_
timestamp 1753371985
transform 1 0 21168 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2040_
timestamp 1751532043
transform 1 0 19936 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2041_
timestamp 1751534193
transform 1 0 23520 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2042_
timestamp 1751534193
transform -1 0 21840 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2043_
timestamp 1753441877
transform -1 0 20944 0 1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2044_
timestamp 1753371985
transform 1 0 18704 0 1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2045_
timestamp 1751532043
transform 1 0 16464 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2046_
timestamp 1751534193
transform -1 0 19488 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2047_
timestamp 1753441877
transform -1 0 19712 0 -1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2048_
timestamp 1753371985
transform 1 0 17584 0 -1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2049_
timestamp 1751532043
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2050_
timestamp 1753441877
transform 1 0 18704 0 -1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2051_
timestamp 1753371985
transform 1 0 17248 0 -1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2052_
timestamp 1751532043
transform -1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2053_
timestamp 1751534193
transform -1 0 20832 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2054_
timestamp 1753441877
transform 1 0 17696 0 -1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2055_
timestamp 1753371985
transform 1 0 17248 0 1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2056_
timestamp 1751532043
transform -1 0 16912 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2057_
timestamp 1751534193
transform -1 0 20384 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2058_
timestamp 1753441877
transform 1 0 18368 0 1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2059_
timestamp 1753371985
transform 1 0 17248 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2060_
timestamp 1751532043
transform 1 0 17920 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2061_
timestamp 1751534193
transform -1 0 20160 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2062_
timestamp 1753441877
transform 1 0 18368 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2063_
timestamp 1753371985
transform -1 0 20608 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2064_
timestamp 1751532043
transform 1 0 19712 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2065_
timestamp 1753441877
transform -1 0 19488 0 1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2066_
timestamp 1753371985
transform -1 0 18592 0 -1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2067_
timestamp 1751532043
transform 1 0 18368 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2068_
timestamp 1751534193
transform 1 0 16912 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2069_
timestamp 1753441877
transform 1 0 18592 0 -1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2070_
timestamp 1753371985
transform 1 0 18592 0 -1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2071_
timestamp 1751532043
transform -1 0 22176 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2072_
timestamp 1751534193
transform -1 0 21392 0 -1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2073_
timestamp 1753441877
transform -1 0 20832 0 -1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2074_
timestamp 1753371985
transform 1 0 18704 0 1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2075_
timestamp 1751532043
transform 1 0 26320 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2076_
timestamp 1753441877
transform -1 0 22288 0 1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2077_
timestamp 1753371985
transform 1 0 19824 0 1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2078_
timestamp 1751532043
transform 1 0 26096 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2079_
timestamp 1753441877
transform 1 0 21280 0 -1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2080_
timestamp 1753371985
transform -1 0 23520 0 -1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2081_
timestamp 1751532043
transform 1 0 26544 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2082_
timestamp 1753441877
transform -1 0 24640 0 -1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2083_
timestamp 1753371985
transform 1 0 22512 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2084_
timestamp 1753182340
transform -1 0 18592 0 1 9408
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2085_
timestamp 1751889408
transform 1 0 17584 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2086_
timestamp 1753182340
transform -1 0 26320 0 -1 10976
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2087_
timestamp 1751889408
transform -1 0 22288 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2088_
timestamp 1751889408
transform 1 0 21392 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2089_
timestamp 1753182340
transform 1 0 16464 0 1 14112
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2090_
timestamp 1751889408
transform -1 0 18704 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2091_
timestamp 1753182340
transform 1 0 23072 0 -1 15680
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _2092_
timestamp 1753891287
transform 1 0 22736 0 -1 14112
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2093_
timestamp 1753960525
transform 1 0 23184 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2094_
timestamp 1753441877
transform 1 0 25088 0 -1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2095_
timestamp 1753371985
transform 1 0 23632 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2096_
timestamp 1751889408
transform -1 0 33040 0 1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2097_
timestamp 1751534193
transform -1 0 16800 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2098_
timestamp 1751532043
transform 1 0 17248 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2099_
timestamp 1751532043
transform 1 0 11984 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _2100_
timestamp 1751905124
transform -1 0 15456 0 1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2101_
timestamp 1753272495
transform 1 0 11984 0 -1 20384
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2102_
timestamp 1753441877
transform 1 0 13776 0 1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2103_
timestamp 1751532043
transform 1 0 13328 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2104_
timestamp 1751889808
transform 1 0 13216 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2105_
timestamp 1751889808
transform 1 0 12320 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2106_
timestamp 1751532043
transform -1 0 20944 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2107_
timestamp 1753868718
transform -1 0 16128 0 1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2108_
timestamp 1753960525
transform 1 0 16128 0 1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2109_
timestamp 1751889808
transform 1 0 17248 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _2110_
timestamp 1752345181
transform 1 0 17248 0 -1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2111_
timestamp 1751531619
transform -1 0 19264 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2112_
timestamp 1753868718
transform 1 0 18256 0 -1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2113_
timestamp 1751534193
transform 1 0 19264 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2114_
timestamp 1753277515
transform 1 0 18256 0 1 20384
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2115_
timestamp 1751889808
transform 1 0 18480 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2116_
timestamp 1751534193
transform 1 0 19264 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2117_
timestamp 1751534193
transform -1 0 18032 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2118_
timestamp 1751889408
transform -1 0 17024 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2119_
timestamp 1753277515
transform -1 0 12992 0 -1 18816
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2120_
timestamp 1751740063
transform -1 0 11984 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2121_
timestamp 1751889408
transform 1 0 13328 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2122_
timestamp 1751740063
transform 1 0 10976 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2123_
timestamp 1751889408
transform 1 0 16464 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2124_
timestamp 1753182340
transform 1 0 11760 0 1 17248
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2125_
timestamp 1751534193
transform -1 0 12096 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2126_
timestamp 1753277515
transform 1 0 13776 0 1 15680
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2127_
timestamp 1751740063
transform -1 0 16912 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2128_
timestamp 1753371985
transform 1 0 14560 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2129_
timestamp 1751740063
transform -1 0 16464 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2130_
timestamp 1751532043
transform -1 0 47264 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2131_
timestamp 1751532043
transform 1 0 8624 0 1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2132_
timestamp 1751534193
transform -1 0 10080 0 -1 43904
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2133_
timestamp 1751532043
transform 1 0 10864 0 1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_2  _2134_
timestamp 1753579406
transform 1 0 9408 0 -1 40768
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2135_
timestamp 1751532043
transform 1 0 21168 0 1 47040
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2136_
timestamp 1751889808
transform -1 0 18032 0 -1 45472
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2137_
timestamp 1751532043
transform 1 0 17584 0 1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2138_
timestamp 1751532043
transform -1 0 17024 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2139_
timestamp 1753868718
transform -1 0 17584 0 1 37632
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2140_
timestamp 1751889808
transform -1 0 17024 0 -1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _2141_
timestamp 1751905124
transform 1 0 12208 0 -1 42336
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2142_
timestamp 1753277515
transform 1 0 11536 0 1 40768
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2143_
timestamp 1751531619
transform 1 0 14336 0 -1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2144_
timestamp 1753441877
transform 1 0 15344 0 1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2145_
timestamp 1751532043
transform -1 0 10976 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2146_
timestamp 1751532043
transform 1 0 13328 0 1 43904
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2147_
timestamp 1751532043
transform 1 0 13776 0 1 43904
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2148_
timestamp 1753868718
transform 1 0 13440 0 -1 42336
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _2149_
timestamp 1753891287
transform 1 0 13328 0 1 40768
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2150_
timestamp 1751740063
transform 1 0 14896 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2151_
timestamp 1753441877
transform 1 0 16464 0 1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2152_
timestamp 1751532043
transform -1 0 17024 0 -1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2153_
timestamp 1753868718
transform -1 0 18368 0 1 43904
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2154_
timestamp 1753441877
transform 1 0 16688 0 1 40768
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2155_
timestamp 1751532043
transform -1 0 17696 0 -1 47040
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2156_
timestamp 1751531619
transform 1 0 18032 0 -1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2157_
timestamp 1751532043
transform 1 0 21168 0 1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2158_
timestamp 1751889808
transform 1 0 17248 0 -1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2159_
timestamp 1751534193
transform -1 0 17136 0 1 43904
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2160_
timestamp 1751532043
transform 1 0 10416 0 1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2161_
timestamp 1753868718
transform 1 0 15456 0 -1 42336
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2162_
timestamp 1753960525
transform 1 0 18480 0 -1 42336
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2163_
timestamp 1751889808
transform -1 0 9184 0 -1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2164_
timestamp 1751532043
transform 1 0 8400 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2165_
timestamp 1751532043
transform -1 0 9856 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_2  _2166_
timestamp 1753579406
transform 1 0 8512 0 1 37632
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2167_
timestamp 1751889808
transform 1 0 10080 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2168_
timestamp 1751889408
transform -1 0 9184 0 -1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2169_
timestamp 1751531619
transform -1 0 11536 0 -1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2170_
timestamp 1753441877
transform 1 0 10640 0 1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2171_
timestamp 1753272495
transform 1 0 9408 0 -1 39200
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2172_
timestamp 1753868718
transform 1 0 9072 0 1 39200
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2173_
timestamp 1751889808
transform 1 0 8512 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _2174_
timestamp 1753172561
transform -1 0 17024 0 -1 40768
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2175_
timestamp 1751531619
transform 1 0 9632 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2176_
timestamp 1751534193
transform -1 0 16240 0 -1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2177_
timestamp 1751532043
transform -1 0 14896 0 -1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2178_
timestamp 1753371985
transform 1 0 14896 0 -1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _2179_
timestamp 1752345181
transform 1 0 10976 0 -1 40768
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2180_
timestamp 1753182340
transform -1 0 15120 0 1 39200
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _2181_
timestamp 1753172561
transform 1 0 12768 0 -1 40768
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2182_
timestamp 1753182340
transform 1 0 12320 0 -1 39200
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2183_
timestamp 1753868718
transform 1 0 17248 0 -1 42336
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2184_
timestamp 1751740063
transform -1 0 16688 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2185_
timestamp 1753868718
transform 1 0 11872 0 1 39200
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2186_
timestamp 1751531619
transform 1 0 17248 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2187_
timestamp 1751531619
transform 1 0 17248 0 -1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2188_
timestamp 1751534193
transform -1 0 12096 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2189_
timestamp 1753277515
transform -1 0 18816 0 -1 37632
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2190_
timestamp 1751889808
transform 1 0 12320 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2191_
timestamp 1751534193
transform 1 0 13216 0 -1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2192_
timestamp 1751534193
transform 1 0 18928 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _2193_
timestamp 1753172561
transform 1 0 21168 0 1 37632
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2194_
timestamp 1753960525
transform -1 0 20944 0 1 37632
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2195_
timestamp 1751531619
transform -1 0 20720 0 -1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2196_
timestamp 1751740063
transform 1 0 18144 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2197_
timestamp 1751534193
transform -1 0 12208 0 -1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2198_
timestamp 1751740063
transform 1 0 10304 0 -1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2199_
timestamp 1751889408
transform -1 0 13104 0 -1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2200_
timestamp 1753182340
transform 1 0 10976 0 -1 42336
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2201_
timestamp 1751534193
transform -1 0 10416 0 -1 42336
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2202_
timestamp 1753182340
transform -1 0 13104 0 1 42336
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2203_
timestamp 1751740063
transform -1 0 13104 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2204_
timestamp 1753182340
transform 1 0 11088 0 -1 43904
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2205_
timestamp 1751534193
transform -1 0 9520 0 1 43904
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2206_
timestamp 1751889408
transform 1 0 13216 0 -1 47040
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2207_
timestamp 1751740063
transform 1 0 10864 0 1 45472
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2208_
timestamp 1753182340
transform -1 0 12880 0 1 45472
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2209_
timestamp 1751534193
transform -1 0 11872 0 1 47040
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2210_
timestamp 1753277515
transform 1 0 13104 0 1 47040
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2211_
timestamp 1751740063
transform -1 0 15456 0 1 47040
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _2212_
timestamp 1752345181
transform -1 0 14336 0 -1 45472
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2213_
timestamp 1753277515
transform -1 0 14896 0 1 45472
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2214_
timestamp 1751740063
transform 1 0 15120 0 -1 45472
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2215_
timestamp 1751740063
transform -1 0 15120 0 -1 45472
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2216_
timestamp 1753277515
transform 1 0 13328 0 1 42336
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2217_
timestamp 1751740063
transform -1 0 16464 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2218_
timestamp 1751889408
transform -1 0 14000 0 -1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2219_
timestamp 1753277515
transform -1 0 8512 0 1 42336
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2220_
timestamp 1751740063
transform -1 0 8064 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2221_
timestamp 1751889408
transform -1 0 7504 0 -1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2222_
timestamp 1751889408
transform -1 0 6720 0 -1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2223_
timestamp 1751740063
transform -1 0 8288 0 -1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2224_
timestamp 1753182340
transform -1 0 7504 0 1 39200
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2225_
timestamp 1751534193
transform -1 0 5936 0 -1 42336
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2226_
timestamp 1753277515
transform -1 0 7840 0 -1 39200
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2227_
timestamp 1751740063
transform -1 0 6272 0 1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2228_
timestamp 1753371985
transform 1 0 7504 0 1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2229_
timestamp 1751740063
transform 1 0 5824 0 -1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2230_
timestamp 1753277515
transform -1 0 23744 0 1 23520
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2231_
timestamp 1751889808
transform -1 0 24528 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2232_
timestamp 1751534193
transform -1 0 23184 0 1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2233_
timestamp 1751889408
transform 1 0 31584 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2234_
timestamp 1751534193
transform 1 0 32368 0 1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2235_
timestamp 1751740063
transform -1 0 32816 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2236_
timestamp 1753868718
transform -1 0 34160 0 -1 32928
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2237_
timestamp 1751534193
transform -1 0 31360 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2238_
timestamp 1751534193
transform -1 0 38192 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2239_
timestamp 1753868718
transform -1 0 32592 0 -1 31360
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2240_
timestamp 1751534193
transform 1 0 31584 0 -1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2241_
timestamp 1751534193
transform -1 0 38752 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2242_
timestamp 1753868718
transform 1 0 33488 0 -1 31360
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2243_
timestamp 1751534193
transform 1 0 34608 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2244_
timestamp 1751534193
transform -1 0 37856 0 1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2245_
timestamp 1753868718
transform 1 0 34160 0 -1 32928
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2246_
timestamp 1751534193
transform -1 0 34496 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2247_
timestamp 1751532043
transform 1 0 10080 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2248_
timestamp 1751532043
transform 1 0 10080 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_2  _2249_
timestamp 1753579406
transform -1 0 12096 0 1 26656
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2250_
timestamp 1751532043
transform -1 0 13552 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2251_
timestamp 1751889808
transform 1 0 12320 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2252_
timestamp 1751534193
transform 1 0 10976 0 -1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2253_
timestamp 1751532043
transform 1 0 13888 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2254_
timestamp 1751532043
transform 1 0 13328 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2255_
timestamp 1751532043
transform 1 0 12208 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_2  _2256_
timestamp 1753579406
transform -1 0 15120 0 -1 31360
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2257_
timestamp 1751534193
transform -1 0 12320 0 -1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2258_
timestamp 1751532043
transform -1 0 15232 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2259_
timestamp 1751532043
transform -1 0 15904 0 1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2260_
timestamp 1751531619
transform -1 0 15680 0 1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2261_
timestamp 1751532043
transform -1 0 19488 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2262_
timestamp 1751889808
transform 1 0 20048 0 -1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2263_
timestamp 1751532043
transform -1 0 22736 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2264_
timestamp 1751532043
transform -1 0 25200 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2265_
timestamp 1751889808
transform 1 0 22736 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2266_
timestamp 1751532043
transform 1 0 18928 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2267_
timestamp 1753868718
transform 1 0 20160 0 -1 31360
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _2268_
timestamp 1751905124
transform -1 0 23184 0 -1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2269_
timestamp 1753277515
transform 1 0 21728 0 1 26656
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2270_
timestamp 1751531619
transform -1 0 23744 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2271_
timestamp 1753441877
transform -1 0 22736 0 -1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2272_
timestamp 1751532043
transform -1 0 21952 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2273_
timestamp 1751532043
transform -1 0 21616 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2274_
timestamp 1751532043
transform 1 0 22400 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2275_
timestamp 1753868718
transform 1 0 21168 0 1 28224
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _2276_
timestamp 1753891287
transform 1 0 21392 0 -1 28224
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2277_
timestamp 1753868718
transform 1 0 21168 0 1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2278_
timestamp 1751532043
transform 1 0 17472 0 1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2279_
timestamp 1753868718
transform 1 0 19488 0 1 32928
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2280_
timestamp 1753441877
transform -1 0 22288 0 1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2281_
timestamp 1753868718
transform 1 0 13776 0 1 31360
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2282_
timestamp 1753868718
transform -1 0 15568 0 1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2283_
timestamp 1751532043
transform 1 0 11760 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2284_
timestamp 1753868718
transform 1 0 13328 0 1 26656
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2285_
timestamp 1753441877
transform 1 0 14672 0 -1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2286_
timestamp 1751531619
transform -1 0 20944 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2287_
timestamp 1751740063
transform 1 0 15792 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2288_
timestamp 1751534193
transform -1 0 19712 0 1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_2  _2289_
timestamp 1753579406
transform 1 0 17248 0 -1 32928
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2290_
timestamp 1751889408
transform 1 0 15792 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2291_
timestamp 1751889408
transform -1 0 15456 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2292_
timestamp 1753868718
transform -1 0 13552 0 -1 31360
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2293_
timestamp 1751889808
transform 1 0 19376 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2294_
timestamp 1753182340
transform -1 0 22848 0 -1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2295_
timestamp 1751534193
transform 1 0 20832 0 -1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2296_
timestamp 1751532043
transform -1 0 15904 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2297_
timestamp 1753868718
transform -1 0 16352 0 -1 31360
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2298_
timestamp 1753441877
transform 1 0 15568 0 1 29792
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2299_
timestamp 1751740063
transform -1 0 21616 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2300_
timestamp 1751889408
transform 1 0 22848 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2301_
timestamp 1751740063
transform 1 0 10640 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2302_
timestamp 1753960525
transform 1 0 14672 0 1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2303_
timestamp 1753441877
transform 1 0 15456 0 1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2304_
timestamp 1753441877
transform -1 0 18032 0 1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2305_
timestamp 1751534193
transform 1 0 17248 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2306_
timestamp 1753277515
transform 1 0 17248 0 -1 31360
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2307_
timestamp 1751889808
transform 1 0 18816 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2308_
timestamp 1751534193
transform -1 0 17024 0 -1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2309_
timestamp 1751534193
transform 1 0 17360 0 1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _2310_
timestamp 1753172561
transform 1 0 20496 0 -1 34496
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2311_
timestamp 1753960525
transform -1 0 21728 0 -1 36064
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2312_
timestamp 1751531619
transform 1 0 19824 0 -1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2313_
timestamp 1751740063
transform 1 0 19600 0 -1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2314_
timestamp 1751534193
transform -1 0 17360 0 1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2315_
timestamp 1751740063
transform -1 0 20160 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2316_
timestamp 1751889408
transform -1 0 20720 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2317_
timestamp 1753182340
transform 1 0 18480 0 1 26656
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2318_
timestamp 1751534193
transform 1 0 19936 0 1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2319_
timestamp 1753182340
transform -1 0 21392 0 -1 28224
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2320_
timestamp 1751740063
transform -1 0 19376 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2321_
timestamp 1753182340
transform 1 0 17248 0 -1 28224
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2322_
timestamp 1751534193
transform 1 0 17920 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2323_
timestamp 1751889408
transform -1 0 19600 0 -1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2324_
timestamp 1751740063
transform -1 0 18816 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2325_
timestamp 1753182340
transform 1 0 16800 0 1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2326_
timestamp 1751534193
transform 1 0 18032 0 1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2327_
timestamp 1753277515
transform -1 0 18816 0 -1 34496
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2328_
timestamp 1751740063
transform 1 0 16240 0 -1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _2329_
timestamp 1752345181
transform -1 0 20048 0 -1 32928
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2330_
timestamp 1753277515
transform -1 0 14896 0 1 32928
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2331_
timestamp 1751740063
transform 1 0 12320 0 1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2332_
timestamp 1751740063
transform -1 0 13776 0 -1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2333_
timestamp 1753277515
transform -1 0 12320 0 1 31360
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2334_
timestamp 1751740063
transform -1 0 12096 0 1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2335_
timestamp 1751889408
transform -1 0 13104 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2336_
timestamp 1753277515
transform -1 0 11760 0 -1 29792
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2337_
timestamp 1751740063
transform -1 0 10192 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2338_
timestamp 1751889408
transform 1 0 11424 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2339_
timestamp 1751889408
transform -1 0 11984 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2340_
timestamp 1751740063
transform -1 0 12768 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2341_
timestamp 1753182340
transform -1 0 12992 0 -1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2342_
timestamp 1751534193
transform 1 0 13328 0 1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2343_
timestamp 1753277515
transform -1 0 9184 0 -1 28224
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2344_
timestamp 1751740063
transform -1 0 8736 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2345_
timestamp 1753371985
transform -1 0 10528 0 -1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2346_
timestamp 1751740063
transform -1 0 8848 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2347_
timestamp 1751532043
transform -1 0 21168 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2348_
timestamp 1753371985
transform 1 0 17360 0 -1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2349_
timestamp 1753960525
transform -1 0 17920 0 1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2350_
timestamp 1751889808
transform 1 0 18032 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2351_
timestamp 1751534193
transform 1 0 18928 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2352_
timestamp 1751532043
transform 1 0 24752 0 1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2353_
timestamp 1751532043
transform 1 0 25200 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2354_
timestamp 1751889808
transform 1 0 29008 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2355_
timestamp 1751532043
transform 1 0 23744 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2356_
timestamp 1751889808
transform 1 0 28448 0 -1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2357_
timestamp 1753277515
transform 1 0 26880 0 -1 40768
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2358_
timestamp 1751889408
transform 1 0 29792 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2359_
timestamp 1751532043
transform -1 0 31584 0 1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2360_
timestamp 1751532043
transform 1 0 30800 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2361_
timestamp 1753868718
transform 1 0 29120 0 1 37632
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2362_
timestamp 1751889808
transform 1 0 30352 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2363_
timestamp 1751531619
transform 1 0 30352 0 1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2364_
timestamp 1751532043
transform -1 0 26880 0 -1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2365_
timestamp 1753868718
transform -1 0 28672 0 1 40768
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2366_
timestamp 1753960525
transform 1 0 27552 0 1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2367_
timestamp 1753441877
transform -1 0 30352 0 1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2368_
timestamp 1753868718
transform -1 0 30576 0 -1 42336
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2369_
timestamp 1751889808
transform 1 0 29792 0 1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2370_
timestamp 1751532043
transform 1 0 23072 0 1 47040
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2371_
timestamp 1751889808
transform 1 0 29008 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2372_
timestamp 1751532043
transform 1 0 27776 0 1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2373_
timestamp 1753868718
transform 1 0 27552 0 1 43904
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2374_
timestamp 1753960525
transform 1 0 29680 0 -1 43904
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2375_
timestamp 1751532043
transform 1 0 32928 0 -1 47040
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2376_
timestamp 1751889808
transform 1 0 32480 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2377_
timestamp 1751889808
transform 1 0 29008 0 1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2378_
timestamp 1751532043
transform -1 0 31248 0 1 43904
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2379_
timestamp 1753868718
transform 1 0 31248 0 1 43904
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2380_
timestamp 1753960525
transform 1 0 32928 0 -1 43904
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2381_
timestamp 1751889808
transform 1 0 31472 0 -1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2382_
timestamp 1751532043
transform 1 0 36064 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2383_
timestamp 1751740063
transform -1 0 37632 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2384_
timestamp 1751532043
transform -1 0 34944 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2385_
timestamp 1753868718
transform -1 0 35504 0 -1 43904
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2386_
timestamp 1751740063
transform -1 0 35952 0 1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2387_
timestamp 1751532043
transform 1 0 36064 0 1 43904
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _2388_
timestamp 1753272495
transform -1 0 35168 0 1 42336
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2389_
timestamp 1753960525
transform -1 0 33152 0 1 42336
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2390_
timestamp 1751534193
transform -1 0 28896 0 -1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2391_
timestamp 1751532043
transform 1 0 31584 0 1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2392_
timestamp 1751531619
transform -1 0 31920 0 1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2393_
timestamp 1753371985
transform 1 0 30240 0 -1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _2394_
timestamp 1753172561
transform 1 0 30800 0 -1 40768
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2395_
timestamp 1753182340
transform -1 0 30576 0 -1 40768
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2396_
timestamp 1751531619
transform 1 0 30016 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2397_
timestamp 1751531619
transform -1 0 36288 0 -1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2398_
timestamp 1751531619
transform 1 0 30576 0 -1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _2399_
timestamp 1753172561
transform -1 0 32368 0 -1 43904
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2400_
timestamp 1753182340
transform -1 0 32032 0 1 42336
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2401_
timestamp 1751531619
transform 1 0 30800 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2402_
timestamp 1751889808
transform 1 0 31584 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2403_
timestamp 1753441877
transform -1 0 33040 0 1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2404_
timestamp 1751531619
transform -1 0 23184 0 1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2405_
timestamp 1751534193
transform -1 0 21504 0 -1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2406_
timestamp 1753277515
transform 1 0 25872 0 -1 37632
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2407_
timestamp 1751889808
transform 1 0 26432 0 -1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2408_
timestamp 1751534193
transform 1 0 27216 0 -1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2409_
timestamp 1751534193
transform 1 0 25760 0 -1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _2410_
timestamp 1753172561
transform 1 0 23856 0 1 37632
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _2411_
timestamp 1753960525
transform -1 0 24304 0 1 36064
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2412_
timestamp 1751531619
transform -1 0 23856 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2413_
timestamp 1751740063
transform -1 0 23408 0 -1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2414_
timestamp 1751534193
transform 1 0 25088 0 -1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2415_
timestamp 1751740063
transform -1 0 24416 0 -1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2416_
timestamp 1751889408
transform 1 0 24416 0 1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2417_
timestamp 1753182340
transform -1 0 26320 0 -1 40768
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2418_
timestamp 1751534193
transform -1 0 25872 0 1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2419_
timestamp 1753182340
transform -1 0 24864 0 -1 40768
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2420_
timestamp 1751740063
transform 1 0 21840 0 -1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2421_
timestamp 1753182340
transform -1 0 23744 0 1 40768
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2422_
timestamp 1751534193
transform 1 0 23744 0 1 40768
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2423_
timestamp 1751889408
transform -1 0 22848 0 -1 42336
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2424_
timestamp 1751740063
transform -1 0 24864 0 -1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2425_
timestamp 1753182340
transform 1 0 21280 0 -1 43904
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2426_
timestamp 1751534193
transform -1 0 22064 0 -1 42336
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2427_
timestamp 1753277515
transform -1 0 24080 0 -1 43904
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2428_
timestamp 1751740063
transform -1 0 23296 0 1 45472
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _2429_
timestamp 1752345181
transform -1 0 25312 0 1 43904
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2430_
timestamp 1753277515
transform -1 0 24752 0 -1 47040
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2431_
timestamp 1751740063
transform -1 0 23072 0 1 47040
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2432_
timestamp 1751740063
transform 1 0 25088 0 -1 45472
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2433_
timestamp 1753277515
transform -1 0 26656 0 -1 47040
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2434_
timestamp 1751740063
transform -1 0 25200 0 1 47040
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2435_
timestamp 1751889408
transform 1 0 26096 0 1 47040
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2436_
timestamp 1753277515
transform 1 0 28224 0 1 47040
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2437_
timestamp 1751740063
transform 1 0 29008 0 1 45472
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2438_
timestamp 1751889408
transform 1 0 30352 0 -1 47040
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2439_
timestamp 1751889408
transform 1 0 31696 0 -1 45472
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2440_
timestamp 1751740063
transform -1 0 31920 0 -1 47040
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2441_
timestamp 1753182340
transform 1 0 30464 0 -1 45472
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2442_
timestamp 1751534193
transform 1 0 30800 0 1 47040
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2443_
timestamp 1753277515
transform 1 0 33376 0 1 43904
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2444_
timestamp 1751740063
transform -1 0 36624 0 1 47040
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2445_
timestamp 1753371985
transform 1 0 34944 0 1 43904
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2446_
timestamp 1751740063
transform 1 0 32032 0 1 47040
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2447_
timestamp 1753277515
transform -1 0 32480 0 -1 25088
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2448_
timestamp 1751889808
transform 1 0 28000 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2449_
timestamp 1751534193
transform 1 0 29680 0 1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2450_
timestamp 1751740063
transform -1 0 39088 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2451_
timestamp 1751889408
transform -1 0 40880 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2452_
timestamp 1753182340
transform 1 0 39312 0 -1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2453_
timestamp 1751534193
transform 1 0 39648 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2454_
timestamp 1751740063
transform 1 0 40768 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2455_
timestamp 1751889408
transform 1 0 41552 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2456_
timestamp 1753182340
transform 1 0 41328 0 1 17248
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2457_
timestamp 1751534193
transform -1 0 40544 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2458_
timestamp 1751889408
transform -1 0 42672 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2459_
timestamp 1751889808
transform 1 0 42672 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2460_
timestamp 1751531619
transform -1 0 43344 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2461_
timestamp 1751740063
transform 1 0 41776 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2462_
timestamp 1751889408
transform 1 0 44016 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2463_
timestamp 1751889808
transform -1 0 43344 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2464_
timestamp 1751531619
transform 1 0 46256 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2465_
timestamp 1751740063
transform -1 0 47376 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2466_
timestamp 1751531619
transform 1 0 45024 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2467_
timestamp 1751889808
transform 1 0 45024 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2468_
timestamp 1751889408
transform 1 0 45808 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2469_
timestamp 1751889408
transform 1 0 45920 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2470_
timestamp 1751534193
transform 1 0 47488 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2471_
timestamp 1753277515
transform 1 0 44352 0 -1 18816
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2472_
timestamp 1751889408
transform 1 0 42336 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2473_
timestamp 1751534193
transform -1 0 43232 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _2474_
timestamp 1751531619
transform -1 0 39088 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2475_
timestamp 1751889808
transform 1 0 36736 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2476_
timestamp 1751889808
transform 1 0 37856 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _2477_
timestamp 1753182340
transform -1 0 38752 0 -1 28224
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _2478_
timestamp 1753441877
transform 1 0 38752 0 -1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2479_
timestamp 1751889408
transform 1 0 38864 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2480_
timestamp 1751534193
transform 1 0 39872 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2481_
timestamp 1751534193
transform -1 0 33936 0 1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2482_
timestamp 1751889808
transform -1 0 32928 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2483_
timestamp 1751532043
transform 1 0 26992 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2484_
timestamp 1751534193
transform -1 0 35168 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2485_
timestamp 1753371985
transform 1 0 27440 0 1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2486_
timestamp 1751889408
transform -1 0 28672 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2487_
timestamp 1751534193
transform 1 0 29008 0 1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2488_
timestamp 1751889808
transform -1 0 32144 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2489_
timestamp 1751532043
transform -1 0 31472 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2490_
timestamp 1753371985
transform 1 0 31472 0 -1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2491_
timestamp 1751889408
transform -1 0 31360 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2492_
timestamp 1751534193
transform -1 0 29792 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2493_
timestamp 1751889808
transform 1 0 33040 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2494_
timestamp 1751532043
transform 1 0 34048 0 -1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2495_
timestamp 1753371985
transform 1 0 33936 0 1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2496_
timestamp 1751889408
transform 1 0 35056 0 1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2497_
timestamp 1751534193
transform 1 0 35840 0 1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _2498_
timestamp 1751889808
transform 1 0 33936 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2499_
timestamp 1751532043
transform -1 0 33936 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _2500_
timestamp 1753371985
transform 1 0 33824 0 -1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2501_
timestamp 1751889408
transform 1 0 34720 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2502_
timestamp 1751534193
transform 1 0 35504 0 1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _2503_
timestamp 1751532043
transform -1 0 12432 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _2504_
timestamp 1753277515
transform 1 0 12432 0 -1 7840
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2505_
timestamp 1751889408
transform 1 0 33712 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2506_
timestamp 1751534193
transform -1 0 39088 0 1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2507_
timestamp 1751740063
transform 1 0 41664 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2508_
timestamp 1751534193
transform -1 0 42672 0 -1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2509_
timestamp 1753868718
transform 1 0 37184 0 1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2510_
timestamp 1751534193
transform 1 0 39648 0 1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2511_
timestamp 1753868718
transform 1 0 38752 0 -1 31360
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2512_
timestamp 1751534193
transform -1 0 39312 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2513_
timestamp 1753868718
transform 1 0 40768 0 -1 31360
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2514_
timestamp 1751534193
transform -1 0 40544 0 -1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2515_
timestamp 1753868718
transform 1 0 39312 0 -1 32928
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2516_
timestamp 1751534193
transform 1 0 40768 0 -1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2517_
timestamp 1751534193
transform 1 0 42224 0 1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2518_
timestamp 1751534193
transform 1 0 42896 0 1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2519_
timestamp 1753868718
transform 1 0 42448 0 1 28224
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2520_
timestamp 1751534193
transform 1 0 43232 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2521_
timestamp 1753868718
transform 1 0 44240 0 -1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2522_
timestamp 1751534193
transform 1 0 45472 0 -1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2523_
timestamp 1753868718
transform 1 0 44688 0 1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2524_
timestamp 1751534193
transform 1 0 45808 0 -1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2525_
timestamp 1753868718
transform 1 0 43120 0 1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2526_
timestamp 1751534193
transform -1 0 44240 0 1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2527_
timestamp 1751889408
transform 1 0 32816 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2528_
timestamp 1751740063
transform -1 0 35392 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2529_
timestamp 1753868718
transform 1 0 33376 0 -1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2530_
timestamp 1751534193
transform 1 0 36176 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2531_
timestamp 1753868718
transform 1 0 32928 0 -1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2532_
timestamp 1751534193
transform 1 0 35392 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _2533_
timestamp 1751889408
transform -1 0 29792 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2534_
timestamp 1751740063
transform 1 0 27664 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2535_
timestamp 1753868718
transform -1 0 28672 0 1 21952
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2536_
timestamp 1751534193
transform -1 0 26656 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2537_
timestamp 1753868718
transform -1 0 30240 0 1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2538_
timestamp 1751534193
transform -1 0 28784 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _2539_
timestamp 1751740063
transform 1 0 38080 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2540_
timestamp 1753868718
transform 1 0 39312 0 -1 25088
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2541_
timestamp 1751534193
transform 1 0 41104 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2542_
timestamp 1753868718
transform 1 0 37968 0 1 25088
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2543_
timestamp 1751534193
transform 1 0 39648 0 1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2544_
timestamp 1753868718
transform 1 0 38192 0 1 23520
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2545_
timestamp 1751534193
transform 1 0 38976 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _2546_
timestamp 1753868718
transform 1 0 39200 0 -1 26656
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2547_
timestamp 1751534193
transform 1 0 40432 0 1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2548_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751632746
transform 1 0 1904 0 -1 29792
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2549_
timestamp 1751632746
transform 1 0 1568 0 -1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2550_
timestamp 1751632746
transform -1 0 9408 0 1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2551_
timestamp 1751632746
transform -1 0 5152 0 -1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2552_
timestamp 1751632746
transform 1 0 4032 0 -1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2553_
timestamp 1751632746
transform 1 0 1568 0 1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2554_
timestamp 1751632746
transform -1 0 8176 0 -1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2555_
timestamp 1751632746
transform 1 0 1568 0 1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2556_
timestamp 1751632746
transform -1 0 4592 0 1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2557_
timestamp 1751632746
transform 1 0 1568 0 -1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2558_
timestamp 1751632746
transform 1 0 1568 0 -1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2559_
timestamp 1751632746
transform 1 0 5824 0 1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2560_
timestamp 1751632746
transform 1 0 6608 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2561_
timestamp 1751632746
transform 1 0 1568 0 1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2562_
timestamp 1751632746
transform 1 0 1568 0 -1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2563_
timestamp 1751632746
transform 1 0 1568 0 1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2564_
timestamp 1751632746
transform -1 0 11312 0 1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2565_
timestamp 1751632746
transform 1 0 7728 0 1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2566_
timestamp 1751632746
transform 1 0 2576 0 -1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2567_
timestamp 1751632746
transform 1 0 8400 0 1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2568_
timestamp 1751632746
transform 1 0 11088 0 -1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2569_
timestamp 1751632746
transform -1 0 14000 0 -1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2570_
timestamp 1751632746
transform 1 0 8512 0 1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2571_
timestamp 1751632746
transform 1 0 1568 0 -1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2572_
timestamp 1751632746
transform 1 0 1568 0 -1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2573_
timestamp 1751632746
transform 1 0 1568 0 -1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2574_
timestamp 1751632746
transform 1 0 1568 0 -1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2575_
timestamp 1751632746
transform 1 0 2240 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2576_
timestamp 1751632746
transform 1 0 6160 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2577_
timestamp 1751632746
transform 1 0 7392 0 1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2578_
timestamp 1751632746
transform -1 0 13104 0 1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2579_
timestamp 1751632746
transform -1 0 13664 0 -1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2580_
timestamp 1751632746
transform 1 0 14896 0 1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2581_
timestamp 1751632746
transform 1 0 8848 0 1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2582_
timestamp 1751632746
transform 1 0 12432 0 -1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2583_
timestamp 1751632746
transform 1 0 9296 0 1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2584_
timestamp 1751632746
transform -1 0 23744 0 -1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2585_
timestamp 1751632746
transform 1 0 6944 0 1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2586_
timestamp 1751632746
transform 1 0 7280 0 1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2587_
timestamp 1751632746
transform 1 0 5488 0 -1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2588_
timestamp 1751632746
transform 1 0 5152 0 -1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2589_
timestamp 1751632746
transform 1 0 35952 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2590_
timestamp 1751632746
transform -1 0 41328 0 1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2591_
timestamp 1751632746
transform 1 0 36176 0 -1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2592_
timestamp 1751632746
transform -1 0 40992 0 1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2593_
timestamp 1751632746
transform 1 0 35952 0 -1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2594_
timestamp 1751632746
transform -1 0 36176 0 -1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2595_
timestamp 1751632746
transform -1 0 35952 0 1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2596_
timestamp 1751632746
transform 1 0 30464 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2597_
timestamp 1751632746
transform -1 0 35952 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2598_
timestamp 1751632746
transform 1 0 40768 0 -1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2599_
timestamp 1751632746
transform 1 0 40320 0 1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2600_
timestamp 1751632746
transform 1 0 40880 0 -1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2601_
timestamp 1751632746
transform 1 0 41328 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2602_
timestamp 1751632746
transform -1 0 47376 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2603_
timestamp 1751632746
transform -1 0 47712 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2604_
timestamp 1751632746
transform -1 0 48384 0 -1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2605_
timestamp 1751632746
transform -1 0 49392 0 1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2606_
timestamp 1751632746
transform -1 0 49392 0 1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2607_
timestamp 1751632746
transform -1 0 48272 0 1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2608_
timestamp 1751632746
transform 1 0 29232 0 1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2609_
timestamp 1751632746
transform 1 0 27104 0 -1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2610_
timestamp 1751632746
transform 1 0 26880 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2611_
timestamp 1751632746
transform 1 0 16912 0 1 3136
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2612_
timestamp 1751632746
transform 1 0 14000 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2613_
timestamp 1751632746
transform 1 0 14000 0 -1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2614_
timestamp 1751632746
transform 1 0 17584 0 -1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2615_
timestamp 1751632746
transform 1 0 19600 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2616_
timestamp 1751632746
transform 1 0 30912 0 1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2617_
timestamp 1751632746
transform 1 0 27776 0 -1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2618_
timestamp 1751632746
transform 1 0 26768 0 -1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2619_
timestamp 1751632746
transform 1 0 25760 0 1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2620_
timestamp 1751632746
transform 1 0 25984 0 -1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2621_
timestamp 1751632746
transform 1 0 25088 0 -1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2622_
timestamp 1751632746
transform 1 0 21728 0 -1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2623_
timestamp 1751632746
transform -1 0 26432 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2624_
timestamp 1751632746
transform 1 0 13440 0 -1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2625_
timestamp 1751632746
transform -1 0 20496 0 1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2626_
timestamp 1751632746
transform 1 0 10192 0 -1 37632
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2627_
timestamp 1751632746
transform 1 0 10080 0 1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2628_
timestamp 1751632746
transform -1 0 20496 0 -1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2629_
timestamp 1751632746
transform 1 0 17920 0 1 45472
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2630_
timestamp 1751632746
transform 1 0 18368 0 -1 45472
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2631_
timestamp 1751632746
transform 1 0 17920 0 1 42336
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2632_
timestamp 1751632746
transform -1 0 16688 0 1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2633_
timestamp 1751632746
transform 1 0 11200 0 -1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2634_
timestamp 1751632746
transform 1 0 8288 0 1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2635_
timestamp 1751632746
transform 1 0 7840 0 1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2636_
timestamp 1751632746
transform -1 0 28784 0 1 29792
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2637_
timestamp 1751632746
transform 1 0 22736 0 1 29792
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2638_
timestamp 1751632746
transform -1 0 26208 0 1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2639_
timestamp 1751632746
transform -1 0 26992 0 1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2640_
timestamp 1751632746
transform 1 0 21728 0 -1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2641_
timestamp 1751632746
transform -1 0 24304 0 1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2642_
timestamp 1751632746
transform -1 0 26544 0 1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2643_
timestamp 1751632746
transform -1 0 28784 0 -1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2644_
timestamp 1751632746
transform 1 0 44688 0 1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2645_
timestamp 1751632746
transform -1 0 49392 0 1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2646_
timestamp 1751632746
transform 1 0 46368 0 1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2647_
timestamp 1751632746
transform 1 0 42896 0 -1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2648_
timestamp 1751632746
transform 1 0 43120 0 -1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2649_
timestamp 1751632746
transform 1 0 29344 0 -1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2650_
timestamp 1751632746
transform 1 0 32928 0 -1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2651_
timestamp 1751632746
transform 1 0 31024 0 1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2652_
timestamp 1751632746
transform -1 0 38080 0 -1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2653_
timestamp 1751632746
transform 1 0 33376 0 -1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2654_
timestamp 1751632746
transform 1 0 36848 0 1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2655_
timestamp 1751632746
transform -1 0 42560 0 1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2656_
timestamp 1751632746
transform -1 0 27552 0 1 3136
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2657_
timestamp 1751632746
transform 1 0 24864 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2658_
timestamp 1751632746
transform 1 0 28112 0 -1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2659_
timestamp 1751632746
transform 1 0 37744 0 1 37632
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2660_
timestamp 1751632746
transform 1 0 38080 0 1 39200
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2661_
timestamp 1751632746
transform 1 0 36400 0 -1 37632
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2662_
timestamp 1751632746
transform 1 0 37520 0 -1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2663_
timestamp 1751632746
transform 1 0 36848 0 1 45472
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2664_
timestamp 1751632746
transform -1 0 39424 0 -1 47040
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2665_
timestamp 1751632746
transform 1 0 36512 0 -1 43904
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2666_
timestamp 1751632746
transform 1 0 36624 0 -1 42336
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2667_
timestamp 1751632746
transform 1 0 29008 0 1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2668_
timestamp 1751632746
transform -1 0 32592 0 1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2669_
timestamp 1751632746
transform 1 0 25760 0 1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2670_
timestamp 1751632746
transform 1 0 24304 0 1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2671_
timestamp 1751632746
transform -1 0 36064 0 1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2672_
timestamp 1751632746
transform -1 0 35952 0 -1 39200
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2673_
timestamp 1751632746
transform 1 0 25872 0 -1 45472
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2674_
timestamp 1751632746
transform 1 0 25200 0 -1 43904
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2675_
timestamp 1751632746
transform 1 0 33600 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2676_
timestamp 1751632746
transform 1 0 40992 0 1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2677_
timestamp 1751632746
transform 1 0 38528 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2678_
timestamp 1751632746
transform 1 0 21168 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2679_
timestamp 1751632746
transform -1 0 33936 0 1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2680_
timestamp 1751632746
transform 1 0 23184 0 1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2681_
timestamp 1751632746
transform 1 0 25088 0 -1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2682_
timestamp 1751632746
transform 1 0 29008 0 1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2683_
timestamp 1751632746
transform -1 0 36176 0 -1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2684_
timestamp 1751632746
transform -1 0 38080 0 -1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2685_
timestamp 1751632746
transform 1 0 39424 0 1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2686_
timestamp 1751632746
transform -1 0 47824 0 1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2687_
timestamp 1751632746
transform 1 0 46368 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2688_
timestamp 1751632746
transform 1 0 45360 0 -1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2689_
timestamp 1751632746
transform -1 0 49392 0 1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2690_
timestamp 1751632746
transform 1 0 44688 0 1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2691_
timestamp 1751632746
transform -1 0 49392 0 1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2692_
timestamp 1751632746
transform -1 0 36624 0 1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2693_
timestamp 1751632746
transform 1 0 35280 0 -1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2694_
timestamp 1751632746
transform 1 0 37968 0 1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2695_
timestamp 1751632746
transform -1 0 42448 0 1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2696_
timestamp 1751632746
transform -1 0 49392 0 1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2697_
timestamp 1751632746
transform 1 0 46368 0 1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2698_
timestamp 1751632746
transform 1 0 42672 0 -1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2699_
timestamp 1751632746
transform -1 0 49392 0 1 37632
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2700_
timestamp 1751632746
transform 1 0 40768 0 -1 39200
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2701_
timestamp 1751632746
transform -1 0 45360 0 -1 47040
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2702_
timestamp 1751632746
transform -1 0 41328 0 1 43904
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2703_
timestamp 1751632746
transform 1 0 39648 0 1 47040
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2704_
timestamp 1751632746
transform 1 0 45360 0 -1 47040
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2705_
timestamp 1751632746
transform 1 0 46368 0 1 45472
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2706_
timestamp 1751632746
transform 1 0 46368 0 1 42336
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2707_
timestamp 1751632746
transform -1 0 49392 0 1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2708_
timestamp 1751632746
transform 1 0 41440 0 1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2709_
timestamp 1751632746
transform -1 0 32032 0 1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2710_
timestamp 1751632746
transform -1 0 28784 0 1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2711_
timestamp 1751632746
transform -1 0 27664 0 1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2712_
timestamp 1751632746
transform 1 0 20048 0 -1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2713_
timestamp 1751632746
transform 1 0 19712 0 -1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2714_
timestamp 1751632746
transform -1 0 19936 0 1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2715_
timestamp 1751632746
transform 1 0 13776 0 -1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2716_
timestamp 1751632746
transform 1 0 13440 0 1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2717_
timestamp 1751632746
transform 1 0 13664 0 1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2718_
timestamp 1751632746
transform 1 0 14000 0 -1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2719_
timestamp 1751632746
transform 1 0 14000 0 -1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2720_
timestamp 1751632746
transform 1 0 14336 0 1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2721_
timestamp 1751632746
transform 1 0 14000 0 -1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2722_
timestamp 1751632746
transform 1 0 20496 0 -1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2723_
timestamp 1751632746
transform 1 0 22848 0 1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2724_
timestamp 1751632746
transform 1 0 22736 0 1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2725_
timestamp 1751632746
transform 1 0 23408 0 1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2726_
timestamp 1751632746
transform -1 0 20944 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2727_
timestamp 1751632746
transform -1 0 20720 0 -1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2728_
timestamp 1751632746
transform 1 0 9632 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2729_
timestamp 1751632746
transform 1 0 10080 0 -1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2730_
timestamp 1751632746
transform -1 0 16128 0 -1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2731_
timestamp 1751632746
transform 1 0 14000 0 -1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2732_
timestamp 1751632746
transform 1 0 46368 0 1 29792
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2733_
timestamp 1751632746
transform 1 0 13328 0 1 37632
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2734_
timestamp 1751632746
transform -1 0 20720 0 -1 39200
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2735_
timestamp 1751632746
transform 1 0 8736 0 1 42336
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2736_
timestamp 1751632746
transform 1 0 9408 0 -1 45472
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2737_
timestamp 1751632746
transform 1 0 10192 0 -1 47040
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2738_
timestamp 1751632746
transform 1 0 14000 0 -1 47040
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2739_
timestamp 1751632746
transform 1 0 14896 0 1 45472
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2740_
timestamp 1751632746
transform 1 0 14000 0 -1 43904
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2741_
timestamp 1751632746
transform 1 0 6160 0 -1 43904
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2742_
timestamp 1751632746
transform 1 0 5488 0 1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2743_
timestamp 1751632746
transform -1 0 6272 0 -1 39200
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2744_
timestamp 1751632746
transform 1 0 5488 0 1 37632
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2745_
timestamp 1751632746
transform 1 0 21728 0 -1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2746_
timestamp 1751632746
transform 1 0 29680 0 1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2747_
timestamp 1751632746
transform 1 0 29008 0 1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2748_
timestamp 1751632746
transform 1 0 33040 0 1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2749_
timestamp 1751632746
transform 1 0 33040 0 1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2750_
timestamp 1751632746
transform 1 0 17808 0 1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2751_
timestamp 1751632746
transform -1 0 20944 0 1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2752_
timestamp 1751632746
transform 1 0 19040 0 -1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2753_
timestamp 1751632746
transform 1 0 16912 0 1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2754_
timestamp 1751632746
transform 1 0 17248 0 -1 29792
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2755_
timestamp 1751632746
transform 1 0 15792 0 1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2756_
timestamp 1751632746
transform 1 0 12992 0 -1 34496
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2757_
timestamp 1751632746
transform 1 0 9968 0 -1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2758_
timestamp 1751632746
transform 1 0 8288 0 1 29792
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2759_
timestamp 1751632746
transform -1 0 14112 0 -1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2760_
timestamp 1751632746
transform 1 0 6944 0 1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2761_
timestamp 1751632746
transform 1 0 7056 0 1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2762_
timestamp 1751632746
transform 1 0 17920 0 1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2763_
timestamp 1751632746
transform 1 0 25760 0 1 37632
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2764_
timestamp 1751632746
transform 1 0 21504 0 -1 37632
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2765_
timestamp 1751632746
transform 1 0 24416 0 1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2766_
timestamp 1751632746
transform -1 0 23520 0 -1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2767_
timestamp 1751632746
transform 1 0 21616 0 1 42336
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2768_
timestamp 1751632746
transform 1 0 21504 0 -1 45472
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2769_
timestamp 1751632746
transform 1 0 20160 0 -1 47040
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2770_
timestamp 1751632746
transform 1 0 23632 0 1 45472
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2771_
timestamp 1751632746
transform -1 0 30352 0 -1 47040
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2772_
timestamp 1751632746
transform 1 0 30016 0 1 45472
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2773_
timestamp 1751632746
transform -1 0 36400 0 -1 47040
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2774_
timestamp 1751632746
transform 1 0 32928 0 -1 45472
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2775_
timestamp 1751632746
transform 1 0 29008 0 1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2776_
timestamp 1751632746
transform 1 0 37072 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2777_
timestamp 1751632746
transform 1 0 37968 0 1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2778_
timestamp 1751632746
transform 1 0 38304 0 1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2779_
timestamp 1751632746
transform -1 0 43904 0 1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2780_
timestamp 1751632746
transform -1 0 47712 0 1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2781_
timestamp 1751632746
transform -1 0 49392 0 1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2782_
timestamp 1751632746
transform 1 0 41440 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2783_
timestamp 1751632746
transform -1 0 41664 0 1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2784_
timestamp 1751632746
transform 1 0 27552 0 -1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2785_
timestamp 1751632746
transform 1 0 28112 0 -1 29792
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2786_
timestamp 1751632746
transform -1 0 38080 0 -1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2787_
timestamp 1751632746
transform -1 0 38080 0 -1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2788_
timestamp 1751632746
transform 1 0 13328 0 1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2789_
timestamp 1751632746
transform 1 0 35728 0 -1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2790_
timestamp 1751632746
transform 1 0 36288 0 -1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2791_
timestamp 1751632746
transform 1 0 39200 0 1 29792
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2792_
timestamp 1751632746
transform 1 0 39872 0 1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2793_
timestamp 1751632746
transform 1 0 42784 0 -1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2794_
timestamp 1751632746
transform -1 0 47712 0 1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2795_
timestamp 1751632746
transform -1 0 48608 0 1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2796_
timestamp 1751632746
transform 1 0 42784 0 -1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2797_
timestamp 1751632746
transform -1 0 36624 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2798_
timestamp 1751632746
transform -1 0 37296 0 -1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2799_
timestamp 1751632746
transform 1 0 25088 0 1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2800_
timestamp 1751632746
transform 1 0 27776 0 -1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2801_
timestamp 1751632746
transform 1 0 41104 0 -1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2802_
timestamp 1751632746
transform 1 0 39200 0 1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2803_
timestamp 1751632746
transform 1 0 38192 0 1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _2804_
timestamp 1751632746
transform 1 0 41104 0 1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2824_
timestamp 1751534193
transform 1 0 43568 0 -1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2825_
timestamp 1751534193
transform -1 0 36624 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _2826_
timestamp 1751534193
transform 1 0 47264 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1272__S dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532392
transform 1 0 25760 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1274__S
timestamp 1751532392
transform 1 0 25872 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1276__S
timestamp 1751532392
transform 1 0 23520 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1278__S
timestamp 1751532392
transform 1 0 26432 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1331__A
timestamp 1751532392
transform -1 0 10528 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1341__A
timestamp 1751532392
transform 1 0 4928 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1393__A
timestamp 1751532392
transform 1 0 9856 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1397__A
timestamp 1751532392
transform 1 0 7952 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1421__A
timestamp 1751532392
transform -1 0 2688 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1432__C
timestamp 1751532392
transform 1 0 6496 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1457__A
timestamp 1751532392
transform 1 0 11760 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1460__A
timestamp 1751532392
transform 1 0 44912 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1461__A
timestamp 1751532392
transform -1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1466__A
timestamp 1751532392
transform -1 0 42784 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1467__C
timestamp 1751532392
transform -1 0 36176 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1467__D
timestamp 1751532392
transform 1 0 36400 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1470__A
timestamp 1751532392
transform -1 0 15232 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1471__A
timestamp 1751532392
transform 1 0 44800 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1473__A
timestamp 1751532392
transform 1 0 26880 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1475__B
timestamp 1751532392
transform 1 0 25312 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1477__A
timestamp 1751532392
transform 1 0 19824 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1479__A
timestamp 1751532392
transform 1 0 21840 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1480__A
timestamp 1751532392
transform -1 0 11536 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1482__A
timestamp 1751532392
transform -1 0 11536 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1483__A
timestamp 1751532392
transform -1 0 11984 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1485__A
timestamp 1751532392
transform -1 0 13328 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1488__A
timestamp 1751532392
transform 1 0 40320 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1490__A
timestamp 1751532392
transform 1 0 23408 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1490__B
timestamp 1751532392
transform 1 0 22400 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1494__A
timestamp 1751532392
transform -1 0 9856 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1495__A
timestamp 1751532392
transform 1 0 44128 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1497__A
timestamp 1751532392
transform 1 0 10528 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1497__B
timestamp 1751532392
transform -1 0 10528 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1498__A
timestamp 1751532392
transform 1 0 12768 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1500__A
timestamp 1751532392
transform 1 0 10864 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1502__A
timestamp 1751532392
transform 1 0 9856 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1507__A
timestamp 1751532392
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1510__A
timestamp 1751532392
transform -1 0 35392 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1514__A
timestamp 1751532392
transform -1 0 37632 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1515__A
timestamp 1751532392
transform 1 0 41888 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1517__A
timestamp 1751532392
transform 1 0 44912 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1523__A
timestamp 1751532392
transform 1 0 42784 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1527__A
timestamp 1751532392
transform 1 0 35616 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1531__A
timestamp 1751532392
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1537__C
timestamp 1751532392
transform 1 0 34272 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1541__A
timestamp 1751532392
transform 1 0 36960 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1544__A
timestamp 1751532392
transform 1 0 26656 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1550__A
timestamp 1751532392
transform -1 0 35056 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1551__A
timestamp 1751532392
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1553__A
timestamp 1751532392
transform 1 0 20272 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1554__A
timestamp 1751532392
transform 1 0 21392 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1562__A
timestamp 1751532392
transform 1 0 44128 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1566__A
timestamp 1751532392
transform 1 0 44240 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1617__A
timestamp 1751532392
transform -1 0 18480 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1649__A
timestamp 1751532392
transform 1 0 25312 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1654__A
timestamp 1751532392
transform -1 0 31248 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1655__A
timestamp 1751532392
transform -1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1657__A
timestamp 1751532392
transform 1 0 16128 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1659__A
timestamp 1751532392
transform 1 0 16016 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1661__A
timestamp 1751532392
transform 1 0 13552 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1667__A
timestamp 1751532392
transform -1 0 21280 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1669__A
timestamp 1751532392
transform 1 0 38192 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1670__A
timestamp 1751532392
transform -1 0 18816 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1672__A
timestamp 1751532392
transform -1 0 39872 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1673__A
timestamp 1751532392
transform -1 0 21056 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1676__A
timestamp 1751532392
transform 1 0 20944 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1681__A
timestamp 1751532392
transform -1 0 15680 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1682__A
timestamp 1751532392
transform 1 0 14560 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1682__B
timestamp 1751532392
transform -1 0 15232 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1683__A
timestamp 1751532392
transform 1 0 15680 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1685__A
timestamp 1751532392
transform 1 0 11648 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1687__A
timestamp 1751532392
transform 1 0 12768 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1691__A
timestamp 1751532392
transform 1 0 42560 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1694__A
timestamp 1751532392
transform 1 0 25984 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1696__A
timestamp 1751532392
transform 1 0 27664 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1698__A
timestamp 1751532392
transform 1 0 39872 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1699__A
timestamp 1751532392
transform 1 0 26544 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1701__A
timestamp 1751532392
transform 1 0 36288 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1702__A
timestamp 1751532392
transform -1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1704__A
timestamp 1751532392
transform 1 0 34496 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1705__A
timestamp 1751532392
transform 1 0 28448 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1709__A
timestamp 1751532392
transform 1 0 23968 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1711__A
timestamp 1751532392
transform 1 0 24080 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1713__A
timestamp 1751532392
transform -1 0 26656 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1715__A
timestamp 1751532392
transform 1 0 26768 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1734__A
timestamp 1751532392
transform 1 0 28000 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1761__A
timestamp 1751532392
transform 1 0 40432 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1762__A
timestamp 1751532392
transform 1 0 39312 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1763__A
timestamp 1751532392
transform -1 0 29456 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1767__A
timestamp 1751532392
transform 1 0 27216 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1768__A
timestamp 1751532392
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1770__A
timestamp 1751532392
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1775__A
timestamp 1751532392
transform 1 0 34272 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1777__A
timestamp 1751532392
transform 1 0 38864 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1779__A
timestamp 1751532392
transform 1 0 37072 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1781__A
timestamp 1751532392
transform 1 0 34384 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1783__A
timestamp 1751532392
transform 1 0 36400 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1788__A
timestamp 1751532392
transform -1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1790__A
timestamp 1751532392
transform 1 0 39424 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1792__A
timestamp 1751532392
transform 1 0 35168 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1794__A
timestamp 1751532392
transform 1 0 36400 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1798__A
timestamp 1751532392
transform 1 0 28224 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1800__A
timestamp 1751532392
transform 1 0 31584 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1802__A
timestamp 1751532392
transform 1 0 30576 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1804__A
timestamp 1751532392
transform 1 0 28112 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1806__A
timestamp 1751532392
transform 1 0 29232 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1810__A
timestamp 1751532392
transform 1 0 34384 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1812__A
timestamp 1751532392
transform 1 0 33264 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1814__A
timestamp 1751532392
transform 1 0 29456 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1816__A
timestamp 1751532392
transform -1 0 27552 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1818__A
timestamp 1751532392
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1821__A
timestamp 1751532392
transform -1 0 41552 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1823__B
timestamp 1751532392
transform -1 0 21168 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1825__A
timestamp 1751532392
transform 1 0 37072 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1830__A
timestamp 1751532392
transform 1 0 33824 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1832__A
timestamp 1751532392
transform -1 0 26992 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1834__A
timestamp 1751532392
transform -1 0 25872 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1836__A
timestamp 1751532392
transform -1 0 30688 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1838__A
timestamp 1751532392
transform 1 0 34832 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1840__A
timestamp 1751532392
transform -1 0 34608 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1926__A
timestamp 1751532392
transform 1 0 45248 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1929__B
timestamp 1751532392
transform -1 0 43568 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1930__A
timestamp 1751532392
transform 1 0 31136 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1933__A
timestamp 1751532392
transform 1 0 45360 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1933__B
timestamp 1751532392
transform -1 0 46032 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1935__A
timestamp 1751532392
transform 1 0 33824 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1937__C
timestamp 1751532392
transform -1 0 41776 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1938__A
timestamp 1751532392
transform 1 0 47264 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1939__A
timestamp 1751532392
transform -1 0 42224 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1941__B
timestamp 1751532392
transform 1 0 46704 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1945__A
timestamp 1751532392
transform 1 0 32704 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1946__B
timestamp 1751532392
transform 1 0 31808 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1947__A
timestamp 1751532392
transform -1 0 36288 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1952__C
timestamp 1751532392
transform 1 0 34832 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1980__A
timestamp 1751532392
transform 1 0 42448 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1998__A
timestamp 1751532392
transform 1 0 41440 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2002__A
timestamp 1751532392
transform 1 0 39872 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2014__S
timestamp 1751532392
transform 1 0 44240 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2032__A
timestamp 1751532392
transform 1 0 23968 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2037__A
timestamp 1751532392
transform -1 0 19488 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2053__A
timestamp 1751532392
transform -1 0 21280 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2068__A
timestamp 1751532392
transform -1 0 16464 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2082__C
timestamp 1751532392
transform -1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2097__A
timestamp 1751532392
transform 1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2111__A
timestamp 1751532392
transform -1 0 19936 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2114__B
timestamp 1751532392
transform -1 0 20384 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2118__B
timestamp 1751532392
transform -1 0 20384 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2186__B
timestamp 1751532392
transform -1 0 16128 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2187__A
timestamp 1751532392
transform -1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2189__B
timestamp 1751532392
transform -1 0 17696 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2193__C
timestamp 1751532392
transform -1 0 22512 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2193__D
timestamp 1751532392
transform -1 0 24416 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2194__C
timestamp 1751532392
transform -1 0 19264 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2235__A
timestamp 1751532392
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2236__A
timestamp 1751532392
transform -1 0 36512 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2238__A
timestamp 1751532392
transform 1 0 43456 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2241__A
timestamp 1751532392
transform 1 0 43904 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2244__A
timestamp 1751532392
transform 1 0 39088 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2304__A
timestamp 1751532392
transform 1 0 18256 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2306__B
timestamp 1751532392
transform 1 0 19824 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2310__C
timestamp 1751532392
transform 1 0 22064 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2310__D
timestamp 1751532392
transform 1 0 22288 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2311__C
timestamp 1751532392
transform 1 0 26432 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2349__D
timestamp 1751532392
transform 1 0 18144 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2403__C
timestamp 1751532392
transform -1 0 33936 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2404__A
timestamp 1751532392
transform 1 0 25312 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2404__B
timestamp 1751532392
transform -1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2406__B
timestamp 1751532392
transform 1 0 27664 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2410__C
timestamp 1751532392
transform 1 0 24640 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2410__D
timestamp 1751532392
transform 1 0 25648 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2411__C
timestamp 1751532392
transform 1 0 24528 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2417__A
timestamp 1751532392
transform 1 0 26320 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2437__A
timestamp 1751532392
transform 1 0 28560 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2444__A
timestamp 1751532392
transform 1 0 36848 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2446__A
timestamp 1751532392
transform 1 0 30128 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2447__B
timestamp 1751532392
transform 1 0 32704 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2450__B
timestamp 1751532392
transform 1 0 40992 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2460__A
timestamp 1751532392
transform -1 0 41776 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2464__A
timestamp 1751532392
transform 1 0 47264 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2468__A
timestamp 1751532392
transform 1 0 46032 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2472__A
timestamp 1751532392
transform 1 0 41664 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2474__A
timestamp 1751532392
transform -1 0 41216 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2474__B
timestamp 1751532392
transform 1 0 40992 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2475__A
timestamp 1751532392
transform -1 0 36736 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2475__B
timestamp 1751532392
transform 1 0 37520 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2476__A
timestamp 1751532392
transform -1 0 37296 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2479__A
timestamp 1751532392
transform -1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2483__A
timestamp 1751532392
transform -1 0 24416 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2490__C
timestamp 1751532392
transform -1 0 31024 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2495__C
timestamp 1751532392
transform 1 0 33824 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2500__C
timestamp 1751532392
transform 1 0 33264 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2504__B
timestamp 1751532392
transform 1 0 12208 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2509__A
timestamp 1751532392
transform 1 0 38304 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2519__A
timestamp 1751532392
transform 1 0 42448 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2521__A
timestamp 1751532392
transform 1 0 46368 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2523__A
timestamp 1751532392
transform 1 0 46144 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2528__A
timestamp 1751532392
transform 1 0 36288 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2529__A
timestamp 1751532392
transform 1 0 37744 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2534__A
timestamp 1751532392
transform -1 0 29456 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2535__A
timestamp 1751532392
transform 1 0 30464 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2539__A
timestamp 1751532392
transform -1 0 35056 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__2540__A
timestamp 1751532392
transform 1 0 40320 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_0_wb_clk_i_A
timestamp 1751532392
transform 1 0 25312 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_2_0__f_wb_clk_i_A
timestamp 1751532392
transform 1 0 17696 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_2_1__f_wb_clk_i_A
timestamp 1751532392
transform -1 0 17472 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_2_2__f_wb_clk_i_A
timestamp 1751532392
transform -1 0 36848 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_2_3__f_wb_clk_i_A
timestamp 1751532392
transform 1 0 36064 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_0_wb_clk_i_A
timestamp 1751532392
transform 1 0 13552 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_1_wb_clk_i_A
timestamp 1751532392
transform 1 0 6048 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_2_wb_clk_i_A
timestamp 1751532392
transform 1 0 10752 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_3_wb_clk_i_A
timestamp 1751532392
transform 1 0 12880 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_4_wb_clk_i_A
timestamp 1751532392
transform 1 0 18704 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_5_wb_clk_i_A
timestamp 1751532392
transform 1 0 16688 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_6_wb_clk_i_A
timestamp 1751532392
transform 1 0 8960 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_7_wb_clk_i_A
timestamp 1751532392
transform 1 0 9296 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_8_wb_clk_i_A
timestamp 1751532392
transform 1 0 8176 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_9_wb_clk_i_A
timestamp 1751532392
transform 1 0 12656 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_10_wb_clk_i_A
timestamp 1751532392
transform 1 0 18032 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_11_wb_clk_i_A
timestamp 1751532392
transform -1 0 22064 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_12_wb_clk_i_A
timestamp 1751532392
transform 1 0 20272 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_13_wb_clk_i_A
timestamp 1751532392
transform 1 0 21616 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_14_wb_clk_i_A
timestamp 1751532392
transform 1 0 32480 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_15_wb_clk_i_A
timestamp 1751532392
transform 1 0 37744 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_16_wb_clk_i_A
timestamp 1751532392
transform 1 0 28896 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_17_wb_clk_i_A
timestamp 1751532392
transform 1 0 38192 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_18_wb_clk_i_A
timestamp 1751532392
transform 1 0 40992 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_19_wb_clk_i_A
timestamp 1751532392
transform 1 0 40320 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_20_wb_clk_i_A
timestamp 1751532392
transform 1 0 41888 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_21_wb_clk_i_A
timestamp 1751532392
transform 1 0 40320 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_22_wb_clk_i_A
timestamp 1751532392
transform 1 0 44240 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_23_wb_clk_i_A
timestamp 1751532392
transform -1 0 42224 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_24_wb_clk_i_A
timestamp 1751532392
transform 1 0 39536 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_25_wb_clk_i_A
timestamp 1751532392
transform -1 0 32480 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_26_wb_clk_i_A
timestamp 1751532392
transform 1 0 36400 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_27_wb_clk_i_A
timestamp 1751532392
transform 1 0 44352 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_28_wb_clk_i_A
timestamp 1751532392
transform 1 0 45472 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_29_wb_clk_i_A
timestamp 1751532392
transform 1 0 44128 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_30_wb_clk_i_A
timestamp 1751532392
transform 1 0 44240 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_31_wb_clk_i_A
timestamp 1751532392
transform 1 0 48160 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_32_wb_clk_i_A
timestamp 1751532392
transform 1 0 34160 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_33_wb_clk_i_A
timestamp 1751532392
transform 1 0 39088 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_34_wb_clk_i_A
timestamp 1751532392
transform 1 0 33600 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_35_wb_clk_i_A
timestamp 1751532392
transform 1 0 32480 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_36_wb_clk_i_A
timestamp 1751532392
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_37_wb_clk_i_A
timestamp 1751532392
transform 1 0 23968 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_38_wb_clk_i_A
timestamp 1751532392
transform 1 0 19936 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_39_wb_clk_i_A
timestamp 1751532392
transform 1 0 21504 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_40_wb_clk_i_A
timestamp 1751532392
transform 1 0 26880 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_41_wb_clk_i_A
timestamp 1751532392
transform 1 0 15792 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_42_wb_clk_i_A
timestamp 1751532392
transform 1 0 7168 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_leaf_43_wb_clk_i_A
timestamp 1751532392
transform 1 0 9632 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload0_A
timestamp 1751532392
transform -1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload1_A
timestamp 1751532392
transform 1 0 35280 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input1_A
timestamp 1751532392
transform -1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input2_A
timestamp 1751532392
transform -1 0 44016 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input3_A
timestamp 1751532392
transform -1 0 38976 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input4_A
timestamp 1751532392
transform -1 0 49392 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input5_A
timestamp 1751532392
transform -1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input6_A
timestamp 1751532392
transform -1 0 49392 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input7_A
timestamp 1751532392
transform -1 0 43792 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input8_A
timestamp 1751532392
transform -1 0 30800 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input9_A
timestamp 1751532392
transform -1 0 39424 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input10_A
timestamp 1751532392
transform -1 0 19152 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0_wb_clk_i dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751661108
transform 1 0 25536 0 -1 28224
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_2_0__f_wb_clk_i
timestamp 1751661108
transform 1 0 15456 0 1 20384
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_2_1__f_wb_clk_i
timestamp 1751661108
transform -1 0 17808 0 1 31360
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_2_2__f_wb_clk_i
timestamp 1751661108
transform 1 0 35504 0 -1 20384
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_2_3__f_wb_clk_i
timestamp 1751661108
transform 1 0 36848 0 1 31360
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_0_wb_clk_i
timestamp 1751661108
transform 1 0 10752 0 -1 15680
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_1_wb_clk_i
timestamp 1751661108
transform -1 0 5264 0 1 18816
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_2_wb_clk_i
timestamp 1751661108
transform 1 0 6384 0 -1 23520
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_3_wb_clk_i
timestamp 1751661108
transform 1 0 13328 0 -1 20384
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_4_wb_clk_i
timestamp 1751661108
transform -1 0 21616 0 -1 25088
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_5_wb_clk_i
timestamp 1751661108
transform 1 0 13888 0 -1 32928
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_6_wb_clk_i
timestamp 1751661108
transform -1 0 7728 0 -1 29792
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_7_wb_clk_i
timestamp 1751661108
transform 1 0 6272 0 1 34496
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_8_wb_clk_i
timestamp 1751661108
transform 1 0 6160 0 -1 40768
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_9_wb_clk_i
timestamp 1751661108
transform -1 0 12320 0 1 43904
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_10_wb_clk_i
timestamp 1751661108
transform 1 0 14896 0 1 42336
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_11_wb_clk_i
timestamp 1751661108
transform 1 0 21280 0 1 43904
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_12_wb_clk_i
timestamp 1751661108
transform 1 0 21168 0 1 39200
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_13_wb_clk_i
timestamp 1751661108
transform 1 0 22064 0 -1 34496
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_14_wb_clk_i
timestamp 1751661108
transform -1 0 31584 0 -1 32928
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_15_wb_clk_i
timestamp 1751661108
transform -1 0 37296 0 -1 36064
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_16_wb_clk_i
timestamp 1751661108
transform -1 0 28672 0 -1 42336
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_17_wb_clk_i
timestamp 1751661108
transform -1 0 35616 0 1 47040
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_18_wb_clk_i
timestamp 1751661108
transform -1 0 40096 0 1 40768
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_19_wb_clk_i
timestamp 1751661108
transform -1 0 46256 0 1 47040
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_20_wb_clk_i
timestamp 1751661108
transform 1 0 45584 0 -1 42336
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_21_wb_clk_i
timestamp 1751661108
transform -1 0 44800 0 -1 37632
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_22_wb_clk_i
timestamp 1751661108
transform 1 0 45584 0 -1 32928
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_23_wb_clk_i
timestamp 1751661108
transform 1 0 41328 0 -1 29792
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_24_wb_clk_i
timestamp 1751661108
transform -1 0 39648 0 1 32928
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_25_wb_clk_i
timestamp 1751661108
transform -1 0 30912 0 -1 25088
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_26_wb_clk_i
timestamp 1751661108
transform -1 0 40096 0 -1 18816
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_27_wb_clk_i
timestamp 1751661108
transform 1 0 40768 0 -1 23520
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_28_wb_clk_i
timestamp 1751661108
transform 1 0 46592 0 1 21952
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_29_wb_clk_i
timestamp 1751661108
transform -1 0 46256 0 -1 15680
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_30_wb_clk_i
timestamp 1751661108
transform -1 0 47936 0 -1 10976
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_31_wb_clk_i
timestamp 1751661108
transform 1 0 45584 0 -1 7840
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_32_wb_clk_i
timestamp 1751661108
transform -1 0 43568 0 -1 7840
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_33_wb_clk_i
timestamp 1751661108
transform -1 0 38640 0 -1 10976
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_34_wb_clk_i
timestamp 1751661108
transform -1 0 32704 0 -1 4704
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_35_wb_clk_i
timestamp 1751661108
transform 1 0 28672 0 -1 12544
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_36_wb_clk_i
timestamp 1751661108
transform 1 0 29904 0 -1 17248
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_37_wb_clk_i
timestamp 1751661108
transform 1 0 25088 0 -1 20384
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_38_wb_clk_i
timestamp 1751661108
transform 1 0 20160 0 -1 15680
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_39_wb_clk_i
timestamp 1751661108
transform 1 0 22176 0 1 7840
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_40_wb_clk_i
timestamp 1751661108
transform -1 0 19152 0 1 7840
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_41_wb_clk_i
timestamp 1751661108
transform -1 0 16352 0 1 7840
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_42_wb_clk_i
timestamp 1751661108
transform -1 0 7392 0 -1 7840
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_leaf_43_wb_clk_i
timestamp 1751661108
transform 1 0 4592 0 -1 12544
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload0 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751896485
transform 1 0 15904 0 -1 29792
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkload1
timestamp 1751661108
transform 1 0 35504 0 -1 29792
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__inv_4  clkload2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751633659
transform 1 0 9968 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  clkload3
timestamp 1751532043
transform 1 0 2016 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_4  clkload4 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751558652
transform -1 0 8064 0 1 25088
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_4  clkload5
timestamp 1751558652
transform 1 0 13328 0 1 20384
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  clkload6
timestamp 1751532043
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkload7
timestamp 1751661108
transform 1 0 21168 0 1 14112
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  clkload8
timestamp 1751532043
transform 1 0 22288 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_4  clkload9
timestamp 1751633659
transform 1 0 13552 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_4  clkload10
timestamp 1751633659
transform 1 0 3696 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  clkload11
timestamp 1751532043
transform 1 0 2688 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_4  clkload12
timestamp 1751558652
transform 1 0 4256 0 1 28224
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  clkload13
timestamp 1751532043
transform 1 0 4816 0 1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_4  clkload14
timestamp 1751633659
transform 1 0 5376 0 -1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload15
timestamp 1751896485
transform 1 0 9520 0 1 45472
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_4  clkload16
timestamp 1751633659
transform 1 0 14896 0 1 43904
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_4  clkload17
timestamp 1751558652
transform 1 0 21280 0 1 45472
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__inv_4  clkload18
timestamp 1751633659
transform -1 0 21952 0 1 40768
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  clkload19
timestamp 1751532043
transform 1 0 23408 0 -1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload20
timestamp 1751896485
transform 1 0 26320 0 1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_4  clkload21
timestamp 1751633659
transform 1 0 36848 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload22
timestamp 1751896485
transform 1 0 47264 0 -1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload23
timestamp 1751896485
transform 1 0 43344 0 1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkload24
timestamp 1751661108
transform 1 0 45136 0 -1 9408
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__inv_4  clkload25
timestamp 1751633659
transform 1 0 48608 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload26
timestamp 1751896485
transform 1 0 39424 0 -1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload27
timestamp 1751896485
transform 1 0 36848 0 1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_4  clkload28
timestamp 1751558652
transform 1 0 29456 0 1 4704
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  clkload29
timestamp 1751532043
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkload30
timestamp 1751661108
transform 1 0 32032 0 1 17248
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload31
timestamp 1751896485
transform -1 0 35840 0 -1 37632
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload32
timestamp 1751896485
transform 1 0 25872 0 1 42336
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkload33
timestamp 1751661108
transform 1 0 33040 0 1 45472
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_4  clkload34
timestamp 1751558652
transform 1 0 35280 0 -1 40768
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkload35
timestamp 1751661108
transform 1 0 42784 0 -1 45472
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload36
timestamp 1751896485
transform 1 0 48272 0 1 43904
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload37
timestamp 1751896485
transform 1 0 42448 0 1 36064
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_4  clkload38
timestamp 1751633659
transform 1 0 48608 0 -1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_4  clkload39
timestamp 1751558652
transform 1 0 41328 0 -1 28224
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__inv_4  clkload40
timestamp 1751633659
transform 1 0 35504 0 -1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_0_6 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532312
transform 1 0 2016 0 1 3136
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_14 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532423
transform 1 0 2912 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_0_19
timestamp 1751532312
transform 1 0 3472 0 1 3136
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_27 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532246
transform 1 0 4368 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_31 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532440
transform 1 0 4816 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_33
timestamp 1751532423
transform 1 0 5040 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_40
timestamp 1751532246
transform 1 0 5824 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_44
timestamp 1751532440
transform 1 0 6272 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_46
timestamp 1751532423
transform 1 0 6496 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_0_51
timestamp 1751532312
transform 1 0 7056 0 1 3136
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_59
timestamp 1751532246
transform 1 0 7952 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_67
timestamp 1751532423
transform 1 0 8848 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_0_70
timestamp 1751532312
transform 1 0 9184 0 1 3136
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_78
timestamp 1751532423
transform 1 0 10080 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_0_83
timestamp 1751532312
transform 1 0 10640 0 1 3136
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_91
timestamp 1751532246
transform 1 0 11536 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_99
timestamp 1751532440
transform 1 0 12432 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_101
timestamp 1751532423
transform 1 0 12656 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_104
timestamp 1751532440
transform 1 0 12992 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_106
timestamp 1751532423
transform 1 0 13216 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_138
timestamp 1751532423
transform 1 0 16800 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_172
timestamp 1751532440
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_174
timestamp 1751532423
transform 1 0 20832 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_206
timestamp 1751532423
transform 1 0 24416 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_244
timestamp 1751532423
transform 1 0 28672 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_269
timestamp 1751532440
transform 1 0 31472 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_271
timestamp 1751532423
transform 1 0 31696 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_373
timestamp 1751532423
transform 1 0 43120 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_376
timestamp 1751532423
transform 1 0 43456 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_388
timestamp 1751532440
transform 1 0 44800 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_390
timestamp 1751532423
transform 1 0 45024 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_428
timestamp 1751532423
transform 1 0 49280 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532351
transform 1 0 1568 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_18
timestamp 1751532351
transform 1 0 3360 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_1_34
timestamp 1751532312
transform 1 0 5152 0 -1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_42
timestamp 1751532423
transform 1 0 6048 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_72
timestamp 1751532351
transform 1 0 9408 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_88
timestamp 1751532351
transform 1 0 11200 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_104
timestamp 1751532246
transform 1 0 12992 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_108
timestamp 1751532440
transform 1 0 13440 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_110
timestamp 1751532423
transform 1 0 13664 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_160
timestamp 1751532440
transform 1 0 19264 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_162
timestamp 1751532423
transform 1 0 19488 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_202
timestamp 1751532440
transform 1 0 23968 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_349
timestamp 1751532423
transform 1 0 40432 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_356
timestamp 1751532423
transform 1 0 41216 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_417
timestamp 1751532440
transform 1 0 48048 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_419
timestamp 1751532423
transform 1 0 48272 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_428
timestamp 1751532423
transform 1 0 49280 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_2_2
timestamp 1751532246
transform 1 0 1568 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_6
timestamp 1751532440
transform 1 0 2016 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_37
timestamp 1751532440
transform 1 0 5488 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_39
timestamp 1751532423
transform 1 0 5712 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_52
timestamp 1751532440
transform 1 0 7168 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_68
timestamp 1751532440
transform 1 0 8960 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_83
timestamp 1751532351
transform 1 0 10640 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_2_99
timestamp 1751532246
transform 1 0 12432 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_103
timestamp 1751532440
transform 1 0 12880 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_2_107
timestamp 1751532246
transform 1 0 13328 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_111
timestamp 1751532440
transform 1 0 13776 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_140
timestamp 1751532440
transform 1 0 17024 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_142
timestamp 1751532423
transform 1 0 17248 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_183
timestamp 1751532423
transform 1 0 21840 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_196
timestamp 1751532423
transform 1 0 23296 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_230
timestamp 1751532440
transform 1 0 27104 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_247
timestamp 1751532440
transform 1 0 29008 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_287
timestamp 1751532423
transform 1 0 33488 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_317
timestamp 1751532440
transform 1 0 36848 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_384
timestamp 1751532423
transform 1 0 44352 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_2
timestamp 1751532351
transform 1 0 1568 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_18
timestamp 1751532246
transform 1 0 3360 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_22
timestamp 1751532440
transform 1 0 3808 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_24
timestamp 1751532423
transform 1 0 4032 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_69
timestamp 1751532423
transform 1 0 9072 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_72
timestamp 1751532246
transform 1 0 9408 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_83
timestamp 1751532246
transform 1 0 10640 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_93
timestamp 1751532351
transform 1 0 11760 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_3_109
timestamp 1751532312
transform 1 0 13552 0 -1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_117
timestamp 1751532440
transform 1 0 14448 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_119
timestamp 1751532423
transform 1 0 14672 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_149
timestamp 1751532440
transform 1 0 18032 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_196
timestamp 1751532440
transform 1 0 23296 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_200
timestamp 1751532440
transform 1 0 23744 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_209
timestamp 1751532423
transform 1 0 24752 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_212
timestamp 1751532440
transform 1 0 25088 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_216
timestamp 1751532440
transform 1 0 25536 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_220
timestamp 1751532246
transform 1 0 25984 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_226
timestamp 1751532246
transform 1 0 26656 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_268
timestamp 1751532423
transform 1 0 31360 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_328
timestamp 1751532440
transform 1 0 38080 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_347
timestamp 1751532440
transform 1 0 40208 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_349
timestamp 1751532423
transform 1 0 40432 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_352
timestamp 1751532423
transform 1 0 40768 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_391
timestamp 1751532440
transform 1 0 45136 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_4_2
timestamp 1751532246
transform 1 0 1568 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_6
timestamp 1751532440
transform 1 0 2016 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_4_14
timestamp 1751532246
transform 1 0 2912 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_18
timestamp 1751532440
transform 1 0 3360 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_20
timestamp 1751532423
transform 1 0 3584 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_52
timestamp 1751532423
transform 1 0 7168 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_174
timestamp 1751532423
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_189
timestamp 1751532440
transform 1 0 22512 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_191
timestamp 1751532423
transform 1 0 22736 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_198
timestamp 1751532423
transform 1 0 23520 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_217
timestamp 1751532440
transform 1 0 25648 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_4_239
timestamp 1751532246
transform 1 0 28112 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_243
timestamp 1751532440
transform 1 0 28560 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_273
timestamp 1751532440
transform 1 0 31920 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_317
timestamp 1751532423
transform 1 0 36848 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_329
timestamp 1751532423
transform 1 0 38192 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_380
timestamp 1751532423
transform 1 0 43904 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_68
timestamp 1751532440
transform 1 0 8960 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_72
timestamp 1751532423
transform 1 0 9408 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_91
timestamp 1751532440
transform 1 0 11536 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_95
timestamp 1751532440
transform 1 0 11984 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_142
timestamp 1751532440
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_144
timestamp 1751532423
transform 1 0 17472 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_179
timestamp 1751532440
transform 1 0 21392 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_181
timestamp 1751532423
transform 1 0 21616 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_209
timestamp 1751532423
transform 1 0 24752 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_252
timestamp 1751532246
transform 1 0 29568 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_256
timestamp 1751532440
transform 1 0 30016 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_258
timestamp 1751532423
transform 1 0 30240 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_277
timestamp 1751532440
transform 1 0 32368 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_279
timestamp 1751532423
transform 1 0 32592 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_282
timestamp 1751532440
transform 1 0 32928 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_286
timestamp 1751532440
transform 1 0 33376 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_290
timestamp 1751532440
transform 1 0 33824 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_292
timestamp 1751532423
transform 1 0 34048 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_316
timestamp 1751532440
transform 1 0 36736 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_320
timestamp 1751532423
transform 1 0 37184 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_335
timestamp 1751532440
transform 1 0 38864 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_339
timestamp 1751532423
transform 1 0 39312 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_383
timestamp 1751532423
transform 1 0 44240 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_428
timestamp 1751532423
transform 1 0 49280 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_6_2
timestamp 1751532312
transform 1 0 1568 0 1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_10
timestamp 1751532246
transform 1 0 2464 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_14
timestamp 1751532423
transform 1 0 2912 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_48
timestamp 1751532246
transform 1 0 6720 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_92
timestamp 1751532440
transform 1 0 11648 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_94
timestamp 1751532423
transform 1 0 11872 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_107
timestamp 1751532440
transform 1 0 13328 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_159
timestamp 1751532440
transform 1 0 19152 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_174
timestamp 1751532423
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_177
timestamp 1751532440
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_179
timestamp 1751532423
transform 1 0 21392 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_218
timestamp 1751532440
transform 1 0 25760 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_226
timestamp 1751532440
transform 1 0 26656 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_241
timestamp 1751532246
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_247
timestamp 1751532440
transform 1 0 29008 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_296
timestamp 1751532440
transform 1 0 34496 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_298
timestamp 1751532423
transform 1 0 34720 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_314
timestamp 1751532423
transform 1 0 36512 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_317
timestamp 1751532423
transform 1 0 36848 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_381
timestamp 1751532440
transform 1 0 44016 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_387
timestamp 1751532440
transform 1 0 44688 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_389
timestamp 1751532423
transform 1 0 44912 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_401
timestamp 1751532423
transform 1 0 46256 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_29
timestamp 1751532423
transform 1 0 4592 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_44
timestamp 1751532440
transform 1 0 6272 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_48
timestamp 1751532423
transform 1 0 6720 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_55
timestamp 1751532423
transform 1 0 7504 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_68
timestamp 1751532440
transform 1 0 8960 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_78
timestamp 1751532246
transform 1 0 10080 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_82
timestamp 1751532423
transform 1 0 10528 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_110
timestamp 1751532440
transform 1 0 13664 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_112
timestamp 1751532423
transform 1 0 13888 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_152
timestamp 1751532440
transform 1 0 18368 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_168
timestamp 1751532440
transform 1 0 20160 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_170
timestamp 1751532423
transform 1 0 20384 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_204
timestamp 1751532246
transform 1 0 24192 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_218
timestamp 1751532440
transform 1 0 25760 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_254
timestamp 1751532246
transform 1 0 29792 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_264
timestamp 1751532440
transform 1 0 30912 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_266
timestamp 1751532423
transform 1 0 31136 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_274
timestamp 1751532246
transform 1 0 32032 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_278
timestamp 1751532440
transform 1 0 32480 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_282
timestamp 1751532440
transform 1 0 32928 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_338
timestamp 1751532423
transform 1 0 39200 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_349
timestamp 1751532423
transform 1 0 40432 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_390
timestamp 1751532423
transform 1 0 45024 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_428
timestamp 1751532423
transform 1 0 49280 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_2
timestamp 1751532246
transform 1 0 1568 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_6
timestamp 1751532423
transform 1 0 2016 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_13
timestamp 1751532246
transform 1 0 2800 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_17
timestamp 1751532423
transform 1 0 3248 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_29
timestamp 1751532246
transform 1 0 4592 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_33
timestamp 1751532440
transform 1 0 5040 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_48
timestamp 1751532246
transform 1 0 6720 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_66
timestamp 1751532351
transform 1 0 8736 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_82
timestamp 1751532423
transform 1 0 10528 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_100
timestamp 1751532246
transform 1 0 12544 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_104
timestamp 1751532423
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_107
timestamp 1751532440
transform 1 0 13328 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_154
timestamp 1751532423
transform 1 0 18592 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_191
timestamp 1751532423
transform 1 0 22736 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_8_219
timestamp 1751532312
transform 1 0 25872 0 1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_227
timestamp 1751532440
transform 1 0 26768 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_235
timestamp 1751532440
transform 1 0 27664 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_237
timestamp 1751532423
transform 1 0 27888 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_8_247
timestamp 1751532312
transform 1 0 29008 0 1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_255
timestamp 1751532440
transform 1 0 29904 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_257
timestamp 1751532423
transform 1 0 30128 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_264
timestamp 1751532246
transform 1 0 30912 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_268
timestamp 1751532423
transform 1 0 31360 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_295
timestamp 1751532440
transform 1 0 34384 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_314
timestamp 1751532423
transform 1 0 36512 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_317
timestamp 1751532440
transform 1 0 36848 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_368
timestamp 1751532440
transform 1 0 42560 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_372
timestamp 1751532423
transform 1 0 43008 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_380
timestamp 1751532440
transform 1 0 43904 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_384
timestamp 1751532423
transform 1 0 44352 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_387
timestamp 1751532440
transform 1 0 44688 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_391
timestamp 1751532423
transform 1 0 45136 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_56
timestamp 1751532440
transform 1 0 7616 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_83
timestamp 1751532440
transform 1 0 10640 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_85
timestamp 1751532423
transform 1 0 10864 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_142
timestamp 1751532440
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_174
timestamp 1751532440
transform 1 0 20832 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_208
timestamp 1751532440
transform 1 0 24640 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_227
timestamp 1751532246
transform 1 0 26768 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_231
timestamp 1751532440
transform 1 0 27216 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_233
timestamp 1751532423
transform 1 0 27440 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_240
timestamp 1751532440
transform 1 0 28224 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_242
timestamp 1751532423
transform 1 0 28448 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_277
timestamp 1751532440
transform 1 0 32368 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_279
timestamp 1751532423
transform 1 0 32592 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_289
timestamp 1751532246
transform 1 0 33712 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_293
timestamp 1751532423
transform 1 0 34160 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_307
timestamp 1751532423
transform 1 0 35728 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_359
timestamp 1751532440
transform 1 0 41552 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_361
timestamp 1751532423
transform 1 0 41776 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_416
timestamp 1751532440
transform 1 0 47936 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_428
timestamp 1751532423
transform 1 0 49280 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_2
timestamp 1751532246
transform 1 0 1568 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_6
timestamp 1751532423
transform 1 0 2016 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_13
timestamp 1751532423
transform 1 0 2800 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_32
timestamp 1751532440
transform 1 0 4928 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_34
timestamp 1751532423
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_91
timestamp 1751532440
transform 1 0 11536 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_104
timestamp 1751532423
transform 1 0 12992 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_10_121
timestamp 1751532312
transform 1 0 14896 0 1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_131
timestamp 1751532440
transform 1 0 16016 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_174
timestamp 1751532423
transform 1 0 20832 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_177
timestamp 1751532440
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_179
timestamp 1751532423
transform 1 0 21392 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_187
timestamp 1751532246
transform 1 0 22288 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_258
timestamp 1751532423
transform 1 0 30240 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_283
timestamp 1751532440
transform 1 0 33040 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_285
timestamp 1751532423
transform 1 0 33264 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_300
timestamp 1751532440
transform 1 0 34944 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_304
timestamp 1751532440
transform 1 0 35392 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_381
timestamp 1751532440
transform 1 0 44016 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_427
timestamp 1751532440
transform 1 0 49168 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_61
timestamp 1751532440
transform 1 0 8176 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_72
timestamp 1751532440
transform 1 0 9408 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_76
timestamp 1751532440
transform 1 0 9856 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_88
timestamp 1751532440
transform 1 0 11200 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_108
timestamp 1751532246
transform 1 0 13440 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_112
timestamp 1751532423
transform 1 0 13888 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_172
timestamp 1751532423
transform 1 0 20608 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_186
timestamp 1751532440
transform 1 0 22176 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_188
timestamp 1751532423
transform 1 0 22400 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_209
timestamp 1751532423
transform 1 0 24752 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_212
timestamp 1751532440
transform 1 0 25088 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_214
timestamp 1751532423
transform 1 0 25312 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_229
timestamp 1751532440
transform 1 0 26992 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_276
timestamp 1751532440
transform 1 0 32256 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_349
timestamp 1751532423
transform 1 0 40432 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_352
timestamp 1751532246
transform 1 0 40768 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_356
timestamp 1751532423
transform 1 0 41216 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_418
timestamp 1751532440
transform 1 0 48160 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_428
timestamp 1751532423
transform 1 0 49280 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_2
timestamp 1751532312
transform 1 0 1568 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_55
timestamp 1751532423
transform 1 0 7504 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_90
timestamp 1751532440
transform 1 0 11424 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_103
timestamp 1751532440
transform 1 0 12880 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_107
timestamp 1751532440
transform 1 0 13328 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_109
timestamp 1751532423
transform 1 0 13552 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_137
timestamp 1751532246
transform 1 0 16688 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_141
timestamp 1751532423
transform 1 0 17136 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_162
timestamp 1751532440
transform 1 0 19488 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_170
timestamp 1751532246
transform 1 0 20384 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_174
timestamp 1751532423
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_189
timestamp 1751532440
transform 1 0 22512 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_224
timestamp 1751532440
transform 1 0 26432 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_228
timestamp 1751532246
transform 1 0 26880 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_232
timestamp 1751532440
transform 1 0 27328 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_234
timestamp 1751532423
transform 1 0 27552 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_303
timestamp 1751532246
transform 1 0 35280 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_307
timestamp 1751532440
transform 1 0 35728 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_317
timestamp 1751532440
transform 1 0 36848 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_319
timestamp 1751532423
transform 1 0 37072 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_327
timestamp 1751532440
transform 1 0 37968 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_329
timestamp 1751532423
transform 1 0 38192 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_337
timestamp 1751532440
transform 1 0 39088 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_347
timestamp 1751532440
transform 1 0 40208 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_351
timestamp 1751532423
transform 1 0 40656 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_397
timestamp 1751532246
transform 1 0 45808 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_401
timestamp 1751532423
transform 1 0 46256 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_13_2
timestamp 1751532312
transform 1 0 1568 0 -1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_10
timestamp 1751532423
transform 1 0 2464 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_38
timestamp 1751532440
transform 1 0 5600 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_62
timestamp 1751532440
transform 1 0 8288 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_83
timestamp 1751532246
transform 1 0 10640 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_114
timestamp 1751532351
transform 1 0 14112 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_130
timestamp 1751532440
transform 1 0 15904 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_142
timestamp 1751532246
transform 1 0 17248 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_162
timestamp 1751532440
transform 1 0 19488 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_205
timestamp 1751532246
transform 1 0 24304 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_209
timestamp 1751532423
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_222
timestamp 1751532246
transform 1 0 26208 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_226
timestamp 1751532423
transform 1 0 26656 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_254
timestamp 1751532351
transform 1 0 29792 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_270
timestamp 1751532246
transform 1 0 31584 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_282
timestamp 1751532246
transform 1 0 32928 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_286
timestamp 1751532423
transform 1 0 33376 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_298
timestamp 1751532440
transform 1 0 34720 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_300
timestamp 1751532423
transform 1 0 34944 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_328
timestamp 1751532440
transform 1 0 38080 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_13_352
timestamp 1751532312
transform 1 0 40768 0 -1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_360
timestamp 1751532440
transform 1 0 41664 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_370
timestamp 1751532423
transform 1 0 42784 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_405
timestamp 1751532440
transform 1 0 46704 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_407
timestamp 1751532423
transform 1 0 46928 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_419
timestamp 1751532423
transform 1 0 48272 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_37
timestamp 1751532440
transform 1 0 5488 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_39
timestamp 1751532423
transform 1 0 5712 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_84
timestamp 1751532246
transform 1 0 10752 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_101
timestamp 1751532246
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_107
timestamp 1751532423
transform 1 0 13328 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_146
timestamp 1751532440
transform 1 0 17696 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_202
timestamp 1751532246
transform 1 0 23968 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_206
timestamp 1751532440
transform 1 0 24416 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_14_235
timestamp 1751532312
transform 1 0 27664 0 1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_243
timestamp 1751532440
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_247
timestamp 1751532423
transform 1 0 29008 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_266
timestamp 1751532440
transform 1 0 31136 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_268
timestamp 1751532423
transform 1 0 31360 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_282
timestamp 1751532246
transform 1 0 32928 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_286
timestamp 1751532440
transform 1 0 33376 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_295
timestamp 1751532246
transform 1 0 34384 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_299
timestamp 1751532440
transform 1 0 34832 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_312
timestamp 1751532440
transform 1 0 36288 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_314
timestamp 1751532423
transform 1 0 36512 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_401
timestamp 1751532423
transform 1 0 46256 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_2
timestamp 1751532246
transform 1 0 1568 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_6
timestamp 1751532440
transform 1 0 2016 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_15_14
timestamp 1751532312
transform 1 0 2912 0 -1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_22
timestamp 1751532246
transform 1 0 3808 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_26
timestamp 1751532423
transform 1 0 4256 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_38
timestamp 1751532440
transform 1 0 5600 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_47
timestamp 1751532440
transform 1 0 6608 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_49
timestamp 1751532423
transform 1 0 6832 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_57
timestamp 1751532440
transform 1 0 7728 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_15_61
timestamp 1751532312
transform 1 0 8176 0 -1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_69
timestamp 1751532423
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_72
timestamp 1751532423
transform 1 0 9408 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_109
timestamp 1751532440
transform 1 0 13552 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_138
timestamp 1751532440
transform 1 0 16800 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_152
timestamp 1751532440
transform 1 0 18368 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_164
timestamp 1751532440
transform 1 0 19712 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_193
timestamp 1751532423
transform 1 0 22960 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_209
timestamp 1751532423
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_218
timestamp 1751532246
transform 1 0 25760 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_15_226
timestamp 1751532312
transform 1 0 26656 0 -1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_234
timestamp 1751532440
transform 1 0 27552 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_263
timestamp 1751532423
transform 1 0 30800 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_275
timestamp 1751532246
transform 1 0 32144 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_279
timestamp 1751532423
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_289
timestamp 1751532440
transform 1 0 33712 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_319
timestamp 1751532440
transform 1 0 37072 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_321
timestamp 1751532423
transform 1 0 37296 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_324
timestamp 1751532246
transform 1 0 37632 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_328
timestamp 1751532423
transform 1 0 38080 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_347
timestamp 1751532440
transform 1 0 40208 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_349
timestamp 1751532423
transform 1 0 40432 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_352
timestamp 1751532246
transform 1 0 40768 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_356
timestamp 1751532440
transform 1 0 41216 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_358
timestamp 1751532423
transform 1 0 41440 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_375
timestamp 1751532423
transform 1 0 43344 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_408
timestamp 1751532440
transform 1 0 47040 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_419
timestamp 1751532423
transform 1 0 48272 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_428
timestamp 1751532423
transform 1 0 49280 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_2
timestamp 1751532246
transform 1 0 1568 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_6
timestamp 1751532440
transform 1 0 2016 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_37
timestamp 1751532423
transform 1 0 5488 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_55
timestamp 1751532246
transform 1 0 7504 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_59
timestamp 1751532440
transform 1 0 7952 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_61
timestamp 1751532423
transform 1 0 8176 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_89
timestamp 1751532423
transform 1 0 11312 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_96
timestamp 1751532312
transform 1 0 12096 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_104
timestamp 1751532423
transform 1 0 12992 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_107
timestamp 1751532440
transform 1 0 13328 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_125
timestamp 1751532312
transform 1 0 15344 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_133
timestamp 1751532440
transform 1 0 16240 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_170
timestamp 1751532423
transform 1 0 20384 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_177
timestamp 1751532423
transform 1 0 21168 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_188
timestamp 1751532440
transform 1 0 22400 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_190
timestamp 1751532423
transform 1 0 22624 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_211
timestamp 1751532440
transform 1 0 24976 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_213
timestamp 1751532423
transform 1 0 25200 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_297
timestamp 1751532440
transform 1 0 34608 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_299
timestamp 1751532423
transform 1 0 34832 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_311
timestamp 1751532440
transform 1 0 36176 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_350
timestamp 1751532440
transform 1 0 40544 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_352
timestamp 1751532423
transform 1 0 40768 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_380
timestamp 1751532440
transform 1 0 43904 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_384
timestamp 1751532423
transform 1 0 44352 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_420
timestamp 1751532246
transform 1 0 48384 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_424
timestamp 1751532440
transform 1 0 48832 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_426
timestamp 1751532423
transform 1 0 49056 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_40
timestamp 1751532440
transform 1 0 5824 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_58
timestamp 1751532440
transform 1 0 7840 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_60
timestamp 1751532423
transform 1 0 8064 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_68
timestamp 1751532440
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_139
timestamp 1751532423
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_142
timestamp 1751532440
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_144
timestamp 1751532423
transform 1 0 17472 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_165
timestamp 1751532440
transform 1 0 19824 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_17_212
timestamp 1751532312
transform 1 0 25088 0 -1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_240
timestamp 1751532423
transform 1 0 28224 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_253
timestamp 1751532440
transform 1 0 29680 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_282
timestamp 1751532440
transform 1 0 32928 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_313
timestamp 1751532440
transform 1 0 36400 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_317
timestamp 1751532440
transform 1 0 36848 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_321
timestamp 1751532440
transform 1 0 37296 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_329
timestamp 1751532423
transform 1 0 38192 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_352
timestamp 1751532440
transform 1 0 40768 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_356
timestamp 1751532246
transform 1 0 41216 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_376
timestamp 1751532246
transform 1 0 43456 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_380
timestamp 1751532423
transform 1 0 43904 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_388
timestamp 1751532440
transform 1 0 44800 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_17_411
timestamp 1751532312
transform 1 0 47376 0 -1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_419
timestamp 1751532423
transform 1 0 48272 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_422
timestamp 1751532423
transform 1 0 48608 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_37
timestamp 1751532440
transform 1 0 5488 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_59
timestamp 1751532423
transform 1 0 7952 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_74
timestamp 1751532440
transform 1 0 9632 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_18_78
timestamp 1751532312
transform 1 0 10080 0 1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_104
timestamp 1751532423
transform 1 0 12992 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_114
timestamp 1751532246
transform 1 0 14112 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_142
timestamp 1751532423
transform 1 0 17248 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_149
timestamp 1751532440
transform 1 0 18032 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_151
timestamp 1751532423
transform 1 0 18256 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_158
timestamp 1751532440
transform 1 0 19040 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_18_162
timestamp 1751532312
transform 1 0 19488 0 1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_170
timestamp 1751532246
transform 1 0 20384 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_174
timestamp 1751532423
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_187
timestamp 1751532440
transform 1 0 22288 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_205
timestamp 1751532423
transform 1 0 24304 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_236
timestamp 1751532440
transform 1 0 27776 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_240
timestamp 1751532246
transform 1 0 28224 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_244
timestamp 1751532423
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_312
timestamp 1751532440
transform 1 0 36288 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_314
timestamp 1751532423
transform 1 0 36512 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_374
timestamp 1751532423
transform 1 0 43232 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_382
timestamp 1751532440
transform 1 0 44128 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_384
timestamp 1751532423
transform 1 0 44352 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_387
timestamp 1751532440
transform 1 0 44688 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_389
timestamp 1751532423
transform 1 0 44912 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_397
timestamp 1751532440
transform 1 0 45808 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_401
timestamp 1751532423
transform 1 0 46256 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_2
timestamp 1751532246
transform 1 0 1568 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_16
timestamp 1751532423
transform 1 0 3136 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_63
timestamp 1751532246
transform 1 0 8400 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_67
timestamp 1751532440
transform 1 0 8848 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_69
timestamp 1751532423
transform 1 0 9072 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_19_72
timestamp 1751532351
transform 1 0 9408 0 -1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_88
timestamp 1751532440
transform 1 0 11200 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_104
timestamp 1751532440
transform 1 0 12992 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_149
timestamp 1751532440
transform 1 0 18032 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_162
timestamp 1751532440
transform 1 0 19488 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_166
timestamp 1751532440
transform 1 0 19936 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_170
timestamp 1751532440
transform 1 0 20384 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_172
timestamp 1751532423
transform 1 0 20608 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_177
timestamp 1751532423
transform 1 0 21168 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_198
timestamp 1751532246
transform 1 0 23520 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_212
timestamp 1751532246
transform 1 0 25088 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_216
timestamp 1751532440
transform 1 0 25536 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_224
timestamp 1751532246
transform 1 0 26432 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_228
timestamp 1751532440
transform 1 0 26880 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_230
timestamp 1751532423
transform 1 0 27104 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_266
timestamp 1751532440
transform 1 0 31136 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_268
timestamp 1751532423
transform 1 0 31360 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_293
timestamp 1751532423
transform 1 0 34160 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_346
timestamp 1751532440
transform 1 0 40096 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_373
timestamp 1751532440
transform 1 0 43120 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_405
timestamp 1751532423
transform 1 0 46704 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_418
timestamp 1751532440
transform 1 0 48160 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_2
timestamp 1751532440
transform 1 0 1568 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_44
timestamp 1751532440
transform 1 0 6272 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_46
timestamp 1751532423
transform 1 0 6496 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_101
timestamp 1751532440
transform 1 0 12656 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_142
timestamp 1751532246
transform 1 0 17248 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_244
timestamp 1751532423
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_258
timestamp 1751532423
transform 1 0 30240 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_317
timestamp 1751532440
transform 1 0 36848 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_353
timestamp 1751532423
transform 1 0 40880 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_387
timestamp 1751532440
transform 1 0 44688 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_391
timestamp 1751532440
transform 1 0 45136 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_395
timestamp 1751532440
transform 1 0 45584 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_399
timestamp 1751532440
transform 1 0 46032 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_401
timestamp 1751532423
transform 1 0 46256 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_69
timestamp 1751532423
transform 1 0 9072 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_72
timestamp 1751532351
transform 1 0 9408 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_132
timestamp 1751532423
transform 1 0 16128 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_166
timestamp 1751532440
transform 1 0 19936 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_170
timestamp 1751532246
transform 1 0 20384 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_174
timestamp 1751532423
transform 1 0 20832 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_177
timestamp 1751532440
transform 1 0 21168 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_188
timestamp 1751532423
transform 1 0 22400 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_195
timestamp 1751532440
transform 1 0 23184 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_199
timestamp 1751532440
transform 1 0 23632 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_201
timestamp 1751532423
transform 1 0 23856 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_275
timestamp 1751532440
transform 1 0 32144 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_279
timestamp 1751532423
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_282
timestamp 1751532440
transform 1 0 32928 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_304
timestamp 1751532423
transform 1 0 35392 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_337
timestamp 1751532440
transform 1 0 39088 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_359
timestamp 1751532423
transform 1 0 41552 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_366
timestamp 1751532440
transform 1 0 42336 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_390
timestamp 1751532440
transform 1 0 45024 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_394
timestamp 1751532440
transform 1 0 45472 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_396
timestamp 1751532423
transform 1 0 45696 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_2
timestamp 1751532440
transform 1 0 1568 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_37
timestamp 1751532440
transform 1 0 5488 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_22_59
timestamp 1751532312
transform 1 0 7952 0 1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_67
timestamp 1751532246
transform 1 0 8848 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_165
timestamp 1751532246
transform 1 0 19824 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_258
timestamp 1751532440
transform 1 0 30240 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_310
timestamp 1751532440
transform 1 0 36064 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_314
timestamp 1751532423
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_323
timestamp 1751532440
transform 1 0 37520 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_387
timestamp 1751532423
transform 1 0 44688 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_426
timestamp 1751532440
transform 1 0 49056 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_428
timestamp 1751532423
transform 1 0 49280 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_29
timestamp 1751532246
transform 1 0 4592 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_33
timestamp 1751532440
transform 1 0 5040 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_42
timestamp 1751532423
transform 1 0 6048 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_57
timestamp 1751532312
transform 1 0 7728 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_65
timestamp 1751532246
transform 1 0 8624 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_69
timestamp 1751532423
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_72
timestamp 1751532440
transform 1 0 9408 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_86
timestamp 1751532440
transform 1 0 10976 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_88
timestamp 1751532423
transform 1 0 11200 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_91
timestamp 1751532440
transform 1 0 11536 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_126
timestamp 1751532423
transform 1 0 15456 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_138
timestamp 1751532440
transform 1 0 16800 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_207
timestamp 1751532440
transform 1 0 24528 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_209
timestamp 1751532423
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_218
timestamp 1751532440
transform 1 0 25760 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_226
timestamp 1751532440
transform 1 0 26656 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_230
timestamp 1751532246
transform 1 0 27104 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_234
timestamp 1751532440
transform 1 0 27552 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_274
timestamp 1751532246
transform 1 0 32032 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_282
timestamp 1751532440
transform 1 0 32928 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_317
timestamp 1751532423
transform 1 0 36848 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_348
timestamp 1751532440
transform 1 0 40320 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_352
timestamp 1751532440
transform 1 0 40768 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_354
timestamp 1751532423
transform 1 0 40992 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_363
timestamp 1751532423
transform 1 0 42000 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_371
timestamp 1751532423
transform 1 0 42896 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_378
timestamp 1751532440
transform 1 0 43680 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_382
timestamp 1751532440
transform 1 0 44128 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_386
timestamp 1751532440
transform 1 0 44576 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_408
timestamp 1751532440
transform 1 0 47040 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_419
timestamp 1751532423
transform 1 0 48272 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_2
timestamp 1751532246
transform 1 0 1568 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_6
timestamp 1751532423
transform 1 0 2016 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_37
timestamp 1751532440
transform 1 0 5488 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_39
timestamp 1751532423
transform 1 0 5712 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_118
timestamp 1751532440
transform 1 0 14560 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_120
timestamp 1751532423
transform 1 0 14784 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_148
timestamp 1751532440
transform 1 0 17920 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_152
timestamp 1751532423
transform 1 0 18368 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_166
timestamp 1751532440
transform 1 0 19936 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_168
timestamp 1751532423
transform 1 0 20160 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_177
timestamp 1751532440
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_185
timestamp 1751532440
transform 1 0 22064 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_187
timestamp 1751532423
transform 1 0 22288 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_190
timestamp 1751532246
transform 1 0 22624 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_194
timestamp 1751532423
transform 1 0 23072 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_222
timestamp 1751532246
transform 1 0 26208 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_226
timestamp 1751532423
transform 1 0 26656 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_229
timestamp 1751532246
transform 1 0 26992 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_244
timestamp 1751532423
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_247
timestamp 1751532440
transform 1 0 29008 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_258
timestamp 1751532440
transform 1 0 30240 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_262
timestamp 1751532440
transform 1 0 30688 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_313
timestamp 1751532440
transform 1 0 36400 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_356
timestamp 1751532440
transform 1 0 41216 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_401
timestamp 1751532440
transform 1 0 46256 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_403
timestamp 1751532423
transform 1 0 46480 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_2
timestamp 1751532246
transform 1 0 1568 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_6
timestamp 1751532423
transform 1 0 2016 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_13
timestamp 1751532246
transform 1 0 2800 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_17
timestamp 1751532423
transform 1 0 3248 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_29
timestamp 1751532440
transform 1 0 4592 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_78
timestamp 1751532440
transform 1 0 10080 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_82
timestamp 1751532440
transform 1 0 10528 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_86
timestamp 1751532440
transform 1 0 10976 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_88
timestamp 1751532423
transform 1 0 11200 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_102
timestamp 1751532440
transform 1 0 12768 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_104
timestamp 1751532423
transform 1 0 12992 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_119
timestamp 1751532440
transform 1 0 14672 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_121
timestamp 1751532423
transform 1 0 14896 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_136
timestamp 1751532440
transform 1 0 16576 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_142
timestamp 1751532423
transform 1 0 17248 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_153
timestamp 1751532440
transform 1 0 18480 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_163
timestamp 1751532440
transform 1 0 19600 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_167
timestamp 1751532246
transform 1 0 20048 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_171
timestamp 1751532440
transform 1 0 20496 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_177
timestamp 1751532246
transform 1 0 21168 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_181
timestamp 1751532440
transform 1 0 21616 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_25_185
timestamp 1751532351
transform 1 0 22064 0 -1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_201
timestamp 1751532440
transform 1 0 23856 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_203
timestamp 1751532423
transform 1 0 24080 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_212
timestamp 1751532440
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_234
timestamp 1751532423
transform 1 0 27552 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_259
timestamp 1751532440
transform 1 0 30352 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_261
timestamp 1751532423
transform 1 0 30576 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_288
timestamp 1751532440
transform 1 0 33600 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_292
timestamp 1751532440
transform 1 0 34048 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_294
timestamp 1751532423
transform 1 0 34272 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_297
timestamp 1751532440
transform 1 0 34608 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_334
timestamp 1751532440
transform 1 0 38752 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_342
timestamp 1751532440
transform 1 0 39648 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_346
timestamp 1751532440
transform 1 0 40096 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_428
timestamp 1751532423
transform 1 0 49280 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_29
timestamp 1751532246
transform 1 0 4592 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_33
timestamp 1751532440
transform 1 0 5040 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_51
timestamp 1751532246
transform 1 0 7056 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_55
timestamp 1751532440
transform 1 0 7504 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_57
timestamp 1751532423
transform 1 0 7728 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_85
timestamp 1751532246
transform 1 0 10864 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_89
timestamp 1751532440
transform 1 0 11312 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_91
timestamp 1751532423
transform 1 0 11536 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_113
timestamp 1751532246
transform 1 0 14000 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_117
timestamp 1751532423
transform 1 0 14448 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_120
timestamp 1751532440
transform 1 0 14784 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_124
timestamp 1751532440
transform 1 0 15232 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_128
timestamp 1751532440
transform 1 0 15680 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_183
timestamp 1751532440
transform 1 0 21840 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_185
timestamp 1751532423
transform 1 0 22064 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_26_207
timestamp 1751532312
transform 1 0 24528 0 1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_215
timestamp 1751532440
transform 1 0 25424 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_237
timestamp 1751532423
transform 1 0 27888 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_286
timestamp 1751532423
transform 1 0 33376 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_294
timestamp 1751532440
transform 1 0 34272 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_310
timestamp 1751532440
transform 1 0 36064 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_314
timestamp 1751532423
transform 1 0 36512 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_374
timestamp 1751532440
transform 1 0 43232 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_378
timestamp 1751532440
transform 1 0 43680 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_380
timestamp 1751532423
transform 1 0 43904 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_397
timestamp 1751532440
transform 1 0 45808 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_399
timestamp 1751532423
transform 1 0 46032 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_424
timestamp 1751532246
transform 1 0 48832 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_428
timestamp 1751532423
transform 1 0 49280 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_27_2
timestamp 1751532312
transform 1 0 1568 0 -1 25088
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_10
timestamp 1751532440
transform 1 0 2464 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_26
timestamp 1751532423
transform 1 0 4256 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_61
timestamp 1751532440
transform 1 0 8176 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_63
timestamp 1751532423
transform 1 0 8400 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_27_72
timestamp 1751532246
transform 1 0 9408 0 -1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_76
timestamp 1751532423
transform 1 0 9856 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_128
timestamp 1751532440
transform 1 0 15680 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_181
timestamp 1751532423
transform 1 0 21616 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_209
timestamp 1751532423
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_278
timestamp 1751532440
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_288
timestamp 1751532440
transform 1 0 33600 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_296
timestamp 1751532440
transform 1 0 34496 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_298
timestamp 1751532423
transform 1 0 34720 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_335
timestamp 1751532440
transform 1 0 38864 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_352
timestamp 1751532440
transform 1 0 40768 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_354
timestamp 1751532423
transform 1 0 40992 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_392
timestamp 1751532440
transform 1 0 45248 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_403
timestamp 1751532440
transform 1 0 46480 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_405
timestamp 1751532423
transform 1 0 46704 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_28_29
timestamp 1751532246
transform 1 0 4592 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_33
timestamp 1751532440
transform 1 0 5040 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_48
timestamp 1751532440
transform 1 0 6720 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_50
timestamp 1751532423
transform 1 0 6944 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_60
timestamp 1751532440
transform 1 0 8064 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_100
timestamp 1751532440
transform 1 0 12544 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_104
timestamp 1751532423
transform 1 0 12992 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_107
timestamp 1751532440
transform 1 0 13328 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_109
timestamp 1751532423
transform 1 0 13552 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_137
timestamp 1751532440
transform 1 0 16688 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_172
timestamp 1751532440
transform 1 0 20608 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_174
timestamp 1751532423
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_177
timestamp 1751532440
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_179
timestamp 1751532423
transform 1 0 21392 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_28_184
timestamp 1751532246
transform 1 0 21952 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_188
timestamp 1751532423
transform 1 0 22400 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_222
timestamp 1751532423
transform 1 0 26208 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_243
timestamp 1751532440
transform 1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_274
timestamp 1751532440
transform 1 0 32032 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_278
timestamp 1751532440
transform 1 0 32480 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_282
timestamp 1751532440
transform 1 0 32928 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_284
timestamp 1751532423
transform 1 0 33152 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_314
timestamp 1751532423
transform 1 0 36512 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_317
timestamp 1751532440
transform 1 0 36848 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_319
timestamp 1751532423
transform 1 0 37072 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_326
timestamp 1751532423
transform 1 0 37856 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_365
timestamp 1751532440
transform 1 0 42224 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_381
timestamp 1751532440
transform 1 0 44016 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_391
timestamp 1751532423
transform 1 0 45136 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_29_2
timestamp 1751532312
transform 1 0 1568 0 -1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_10
timestamp 1751532423
transform 1 0 2464 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_29_18
timestamp 1751532312
transform 1 0 3360 0 -1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_26
timestamp 1751532246
transform 1 0 4256 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_30
timestamp 1751532440
transform 1 0 4704 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_47
timestamp 1751532423
transform 1 0 6608 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_55
timestamp 1751532246
transform 1 0 7504 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_59
timestamp 1751532423
transform 1 0 7952 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_67
timestamp 1751532440
transform 1 0 8848 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_69
timestamp 1751532423
transform 1 0 9072 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_82
timestamp 1751532423
transform 1 0 10528 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_90
timestamp 1751532440
transform 1 0 11424 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_92
timestamp 1751532423
transform 1 0 11648 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_103
timestamp 1751532440
transform 1 0 12880 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_126
timestamp 1751532440
transform 1 0 15456 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_130
timestamp 1751532246
transform 1 0 15904 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_134
timestamp 1751532440
transform 1 0 16352 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_138
timestamp 1751532440
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_154
timestamp 1751532246
transform 1 0 18592 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_29_195
timestamp 1751532312
transform 1 0 23184 0 -1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_203
timestamp 1751532423
transform 1 0 24080 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_206
timestamp 1751532440
transform 1 0 24416 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_233
timestamp 1751532423
transform 1 0 27440 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_261
timestamp 1751532440
transform 1 0 30576 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_279
timestamp 1751532423
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_282
timestamp 1751532423
transform 1 0 32928 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_300
timestamp 1751532423
transform 1 0 34944 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_328
timestamp 1751532440
transform 1 0 38080 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_349
timestamp 1751532423
transform 1 0 40432 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_352
timestamp 1751532440
transform 1 0 40768 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_354
timestamp 1751532423
transform 1 0 40992 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_361
timestamp 1751532440
transform 1 0 41776 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_365
timestamp 1751532440
transform 1 0 42224 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_369
timestamp 1751532246
transform 1 0 42672 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_373
timestamp 1751532423
transform 1 0 43120 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_380
timestamp 1751532440
transform 1 0 43904 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_384
timestamp 1751532246
transform 1 0 44352 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_402
timestamp 1751532246
transform 1 0 46368 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_406
timestamp 1751532440
transform 1 0 46816 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_408
timestamp 1751532423
transform 1 0 47040 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_419
timestamp 1751532423
transform 1 0 48272 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_428
timestamp 1751532423
transform 1 0 49280 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_33
timestamp 1751532440
transform 1 0 5040 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_48
timestamp 1751532440
transform 1 0 6720 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_50
timestamp 1751532423
transform 1 0 6944 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_96
timestamp 1751532440
transform 1 0 12096 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_118
timestamp 1751532423
transform 1 0 14560 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_136
timestamp 1751532440
transform 1 0 16576 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_138
timestamp 1751532423
transform 1 0 16800 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_149
timestamp 1751532440
transform 1 0 18032 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_164
timestamp 1751532440
transform 1 0 19712 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_173
timestamp 1751532440
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_181
timestamp 1751532423
transform 1 0 21616 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_196
timestamp 1751532246
transform 1 0 23296 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_200
timestamp 1751532440
transform 1 0 23744 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_235
timestamp 1751532440
transform 1 0 27664 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_244
timestamp 1751532423
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_259
timestamp 1751532440
transform 1 0 30352 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_282
timestamp 1751532440
transform 1 0 32928 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_284
timestamp 1751532423
transform 1 0 33152 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_311
timestamp 1751532440
transform 1 0 36176 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_317
timestamp 1751532440
transform 1 0 36848 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_321
timestamp 1751532440
transform 1 0 37296 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_325
timestamp 1751532423
transform 1 0 37744 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_333
timestamp 1751532440
transform 1 0 38640 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_348
timestamp 1751532423
transform 1 0 40320 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_382
timestamp 1751532440
transform 1 0 44128 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_384
timestamp 1751532423
transform 1 0 44352 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_421
timestamp 1751532440
transform 1 0 48496 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_2
timestamp 1751532423
transform 1 0 1568 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_55
timestamp 1751532423
transform 1 0 7504 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_82
timestamp 1751532246
transform 1 0 10528 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_86
timestamp 1751532423
transform 1 0 10976 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_114
timestamp 1751532246
transform 1 0 14112 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_118
timestamp 1751532423
transform 1 0 14560 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_136
timestamp 1751532440
transform 1 0 16576 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_153
timestamp 1751532423
transform 1 0 18480 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_31_200
timestamp 1751532312
transform 1 0 23744 0 -1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_208
timestamp 1751532440
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_212
timestamp 1751532440
transform 1 0 25088 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_260
timestamp 1751532246
transform 1 0 30464 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_31_302
timestamp 1751532312
transform 1 0 35168 0 -1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_312
timestamp 1751532440
transform 1 0 36288 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_352
timestamp 1751532440
transform 1 0 40768 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_356
timestamp 1751532423
transform 1 0 41216 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_366
timestamp 1751532440
transform 1 0 42336 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_397
timestamp 1751532351
transform 1 0 45808 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_413
timestamp 1751532246
transform 1 0 47600 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_417
timestamp 1751532423
transform 1 0 48048 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_422
timestamp 1751532423
transform 1 0 48608 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_32_2
timestamp 1751532312
transform 1 0 1568 0 1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_10
timestamp 1751532440
transform 1 0 2464 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_47
timestamp 1751532440
transform 1 0 6608 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_49
timestamp 1751532423
transform 1 0 6832 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_32_77
timestamp 1751532312
transform 1 0 9968 0 1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_85
timestamp 1751532440
transform 1 0 10864 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_87
timestamp 1751532423
transform 1 0 11088 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_102
timestamp 1751532440
transform 1 0 12768 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_104
timestamp 1751532423
transform 1 0 12992 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_32_113
timestamp 1751532246
transform 1 0 14000 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_117
timestamp 1751532440
transform 1 0 14448 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_136
timestamp 1751532423
transform 1 0 16576 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_155
timestamp 1751532440
transform 1 0 18704 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_157
timestamp 1751532423
transform 1 0 18928 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_32_164
timestamp 1751532312
transform 1 0 19712 0 1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_172
timestamp 1751532440
transform 1 0 20608 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_174
timestamp 1751532423
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_192
timestamp 1751532351
transform 1 0 22848 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_208
timestamp 1751532423
transform 1 0 24640 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_213
timestamp 1751532440
transform 1 0 25200 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_215
timestamp 1751532423
transform 1 0 25424 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_240
timestamp 1751532440
transform 1 0 28224 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_244
timestamp 1751532423
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_254
timestamp 1751532440
transform 1 0 29792 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_256
timestamp 1751532423
transform 1 0 30016 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_288
timestamp 1751532440
transform 1 0 33600 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_290
timestamp 1751532423
transform 1 0 33824 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_306
timestamp 1751532440
transform 1 0 35616 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_308
timestamp 1751532423
transform 1 0 35840 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_311
timestamp 1751532440
transform 1 0 36176 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_331
timestamp 1751532440
transform 1 0 38416 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_384
timestamp 1751532423
transform 1 0 44352 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_32_414
timestamp 1751532312
transform 1 0 47712 0 1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_32_422
timestamp 1751532246
transform 1 0 48608 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_426
timestamp 1751532423
transform 1 0 49056 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_2
timestamp 1751532440
transform 1 0 1568 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_4
timestamp 1751532423
transform 1 0 1792 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_57
timestamp 1751532440
transform 1 0 7728 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_66
timestamp 1751532440
transform 1 0 8736 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_104
timestamp 1751532351
transform 1 0 12992 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_124
timestamp 1751532440
transform 1 0 15232 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_169
timestamp 1751532246
transform 1 0 20272 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_173
timestamp 1751532423
transform 1 0 20720 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_199
timestamp 1751532440
transform 1 0 23632 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_201
timestamp 1751532423
transform 1 0 23856 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_212
timestamp 1751532440
transform 1 0 25088 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_231
timestamp 1751532423
transform 1 0 27216 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_273
timestamp 1751532246
transform 1 0 31920 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_277
timestamp 1751532440
transform 1 0 32368 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_279
timestamp 1751532423
transform 1 0 32592 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_282
timestamp 1751532246
transform 1 0 32928 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_301
timestamp 1751532440
transform 1 0 35056 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_341
timestamp 1751532440
transform 1 0 39536 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_343
timestamp 1751532423
transform 1 0 39760 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_352
timestamp 1751532440
transform 1 0 40768 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_356
timestamp 1751532423
transform 1 0 41216 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_382
timestamp 1751532423
transform 1 0 44128 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_400
timestamp 1751532440
transform 1 0 46144 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_404
timestamp 1751532440
transform 1 0 46592 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_422
timestamp 1751532246
transform 1 0 48608 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_426
timestamp 1751532440
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_428
timestamp 1751532423
transform 1 0 49280 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_2
timestamp 1751532246
transform 1 0 1568 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_6
timestamp 1751532440
transform 1 0 2016 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_14
timestamp 1751532246
transform 1 0 2912 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_18
timestamp 1751532440
transform 1 0 3360 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_20
timestamp 1751532423
transform 1 0 3584 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_61
timestamp 1751532423
transform 1 0 8176 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_89
timestamp 1751532423
transform 1 0 11312 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_101
timestamp 1751532246
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_107
timestamp 1751532246
transform 1 0 13328 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_111
timestamp 1751532423
transform 1 0 13776 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_137
timestamp 1751532423
transform 1 0 16688 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_163
timestamp 1751532440
transform 1 0 19600 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_167
timestamp 1751532423
transform 1 0 20048 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_188
timestamp 1751532440
transform 1 0 22400 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_190
timestamp 1751532423
transform 1 0 22624 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_247
timestamp 1751532351
transform 1 0 29008 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_263
timestamp 1751532246
transform 1 0 30800 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_267
timestamp 1751532440
transform 1 0 31248 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_269
timestamp 1751532423
transform 1 0 31472 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_312
timestamp 1751532440
transform 1 0 36288 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_314
timestamp 1751532423
transform 1 0 36512 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_317
timestamp 1751532440
transform 1 0 36848 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_319
timestamp 1751532423
transform 1 0 37072 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_337
timestamp 1751532423
transform 1 0 39088 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_371
timestamp 1751532440
transform 1 0 42896 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_384
timestamp 1751532423
transform 1 0 44352 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_398
timestamp 1751532440
transform 1 0 45920 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_29
timestamp 1751532440
transform 1 0 4592 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_41
timestamp 1751532423
transform 1 0 5936 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_35_56
timestamp 1751532312
transform 1 0 7616 0 -1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_64
timestamp 1751532246
transform 1 0 8512 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_68
timestamp 1751532440
transform 1 0 8960 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_35_72
timestamp 1751532312
transform 1 0 9408 0 -1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_82
timestamp 1751532246
transform 1 0 10528 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_156
timestamp 1751532423
transform 1 0 18816 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_179
timestamp 1751532440
transform 1 0 21392 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_223
timestamp 1751532440
transform 1 0 26320 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_233
timestamp 1751532440
transform 1 0 27440 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_237
timestamp 1751532246
transform 1 0 27888 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_241
timestamp 1751532423
transform 1 0 28336 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_35_249
timestamp 1751532312
transform 1 0 29232 0 -1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_263
timestamp 1751532440
transform 1 0 30800 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_267
timestamp 1751532423
transform 1 0 31248 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_279
timestamp 1751532423
transform 1 0 32592 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_282
timestamp 1751532440
transform 1 0 32928 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_286
timestamp 1751532423
transform 1 0 33376 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_298
timestamp 1751532440
transform 1 0 34720 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_345
timestamp 1751532423
transform 1 0 39984 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_369
timestamp 1751532423
transform 1 0 42672 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_403
timestamp 1751532440
transform 1 0 46480 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_418
timestamp 1751532440
transform 1 0 48160 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_428
timestamp 1751532423
transform 1 0 49280 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_36_2
timestamp 1751532312
transform 1 0 1568 0 1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_36_10
timestamp 1751532246
transform 1 0 2464 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_14
timestamp 1751532423
transform 1 0 2912 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_36_22
timestamp 1751532246
transform 1 0 3808 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_26
timestamp 1751532440
transform 1 0 4256 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_44
timestamp 1751532423
transform 1 0 6272 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_72
timestamp 1751532423
transform 1 0 9408 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_80
timestamp 1751532440
transform 1 0 10304 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_174
timestamp 1751532423
transform 1 0 20832 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_202
timestamp 1751532440
transform 1 0 23968 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_242
timestamp 1751532440
transform 1 0 28448 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_244
timestamp 1751532423
transform 1 0 28672 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_281
timestamp 1751532440
transform 1 0 32816 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_314
timestamp 1751532423
transform 1 0 36512 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_342
timestamp 1751532440
transform 1 0 39648 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_383
timestamp 1751532440
transform 1 0 44240 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_387
timestamp 1751532440
transform 1 0 44688 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_389
timestamp 1751532423
transform 1 0 44912 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_394
timestamp 1751532423
transform 1 0 45472 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_428
timestamp 1751532423
transform 1 0 49280 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_37_2
timestamp 1751532246
transform 1 0 1568 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_6
timestamp 1751532423
transform 1 0 2016 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_37_34
timestamp 1751532351
transform 1 0 5152 0 -1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_37_57
timestamp 1751532246
transform 1 0 7728 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_61
timestamp 1751532440
transform 1 0 8176 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_63
timestamp 1751532423
transform 1 0 8400 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_72
timestamp 1751532440
transform 1 0 9408 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_76
timestamp 1751532423
transform 1 0 9856 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_111
timestamp 1751532423
transform 1 0 13776 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_137
timestamp 1751532440
transform 1 0 16688 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_139
timestamp 1751532423
transform 1 0 16912 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_180
timestamp 1751532440
transform 1 0 21504 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_209
timestamp 1751532423
transform 1 0 24752 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_276
timestamp 1751532440
transform 1 0 32256 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_304
timestamp 1751532423
transform 1 0 35392 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_358
timestamp 1751532440
transform 1 0 41440 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_360
timestamp 1751532423
transform 1 0 41664 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_378
timestamp 1751532440
transform 1 0 43680 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_380
timestamp 1751532423
transform 1 0 43904 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_38_2
timestamp 1751532351
transform 1 0 1568 0 1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_38_18
timestamp 1751532351
transform 1 0 3360 0 1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_34
timestamp 1751532423
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_38_37
timestamp 1751532312
transform 1 0 5488 0 1 32928
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_38_45
timestamp 1751532246
transform 1 0 6384 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_49
timestamp 1751532423
transform 1 0 6832 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_88
timestamp 1751532423
transform 1 0 11200 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_96
timestamp 1751532440
transform 1 0 12096 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_128
timestamp 1751532423
transform 1 0 15680 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_156
timestamp 1751532440
transform 1 0 18816 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_173
timestamp 1751532440
transform 1 0 20720 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_177
timestamp 1751532440
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_179
timestamp 1751532423
transform 1 0 21392 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_197
timestamp 1751532423
transform 1 0 23408 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_225
timestamp 1751532440
transform 1 0 26544 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_38_229
timestamp 1751532351
transform 1 0 26992 0 1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_38_247
timestamp 1751532246
transform 1 0 29008 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_251
timestamp 1751532440
transform 1 0 29456 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_280
timestamp 1751532440
transform 1 0 32704 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_282
timestamp 1751532423
transform 1 0 32928 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_310
timestamp 1751532440
transform 1 0 36064 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_314
timestamp 1751532423
transform 1 0 36512 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_348
timestamp 1751532423
transform 1 0 40320 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_365
timestamp 1751532440
transform 1 0 42224 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_382
timestamp 1751532440
transform 1 0 44128 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_384
timestamp 1751532423
transform 1 0 44352 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_39_2
timestamp 1751532351
transform 1 0 1568 0 -1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_39_18
timestamp 1751532351
transform 1 0 3360 0 -1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_34
timestamp 1751532440
transform 1 0 5152 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_36
timestamp 1751532423
transform 1 0 5376 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_100
timestamp 1751532440
transform 1 0 12544 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_131
timestamp 1751532440
transform 1 0 16016 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_170
timestamp 1751532423
transform 1 0 20384 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_218
timestamp 1751532440
transform 1 0 25760 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_222
timestamp 1751532440
transform 1 0 26208 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_226
timestamp 1751532440
transform 1 0 26656 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_39_234
timestamp 1751532312
transform 1 0 27552 0 -1 34496
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_242
timestamp 1751532440
transform 1 0 28448 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_261
timestamp 1751532423
transform 1 0 30576 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_268
timestamp 1751532440
transform 1 0 31360 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_39_272
timestamp 1751532312
transform 1 0 31808 0 -1 34496
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_282
timestamp 1751532440
transform 1 0 32928 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_284
timestamp 1751532423
transform 1 0 33152 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_295
timestamp 1751532440
transform 1 0 34384 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_348
timestamp 1751532440
transform 1 0 40320 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_352
timestamp 1751532423
transform 1 0 40768 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_375
timestamp 1751532440
transform 1 0 43344 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_397
timestamp 1751532440
transform 1 0 45808 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_419
timestamp 1751532423
transform 1 0 48272 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_422
timestamp 1751532423
transform 1 0 48608 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_40_2
timestamp 1751532351
transform 1 0 1568 0 1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_40_18
timestamp 1751532312
transform 1 0 3360 0 1 34496
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_40_26
timestamp 1751532246
transform 1 0 4256 0 1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_30
timestamp 1751532423
transform 1 0 4704 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_37
timestamp 1751532423
transform 1 0 5488 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_69
timestamp 1751532440
transform 1 0 9072 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_73
timestamp 1751532440
transform 1 0 9520 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_75
timestamp 1751532423
transform 1 0 9744 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_40_107
timestamp 1751532312
transform 1 0 13328 0 1 34496
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_130
timestamp 1751532440
transform 1 0 15904 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_134
timestamp 1751532440
transform 1 0 16352 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_136
timestamp 1751532423
transform 1 0 16576 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_139
timestamp 1751532440
transform 1 0 16912 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_141
timestamp 1751532423
transform 1 0 17136 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_177
timestamp 1751532423
transform 1 0 21168 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_216
timestamp 1751532440
transform 1 0 25536 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_274
timestamp 1751532440
transform 1 0 32032 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_297
timestamp 1751532440
transform 1 0 34608 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_354
timestamp 1751532440
transform 1 0 40992 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_356
timestamp 1751532423
transform 1 0 41216 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_372
timestamp 1751532440
transform 1 0 43008 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_380
timestamp 1751532440
transform 1 0 43904 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_382
timestamp 1751532423
transform 1 0 44128 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_397
timestamp 1751532423
transform 1 0 45808 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_41_2
timestamp 1751532351
transform 1 0 1568 0 -1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_41_18
timestamp 1751532351
transform 1 0 3360 0 -1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_61
timestamp 1751532440
transform 1 0 8176 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_63
timestamp 1751532423
transform 1 0 8400 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_83
timestamp 1751532440
transform 1 0 10640 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_41_87
timestamp 1751532246
transform 1 0 11088 0 -1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_91
timestamp 1751532440
transform 1 0 11536 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_41_104
timestamp 1751532246
transform 1 0 12992 0 -1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_135
timestamp 1751532440
transform 1 0 16464 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_137
timestamp 1751532423
transform 1 0 16688 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_149
timestamp 1751532423
transform 1 0 18032 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_162
timestamp 1751532440
transform 1 0 19488 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_164
timestamp 1751532423
transform 1 0 19712 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_41_182
timestamp 1751532246
transform 1 0 21728 0 -1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_186
timestamp 1751532423
transform 1 0 22176 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_189
timestamp 1751532440
transform 1 0 22512 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_201
timestamp 1751532440
transform 1 0 23856 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_205
timestamp 1751532440
transform 1 0 24304 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_209
timestamp 1751532423
transform 1 0 24752 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_212
timestamp 1751532440
transform 1 0 25088 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_222
timestamp 1751532440
transform 1 0 26208 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_237
timestamp 1751532440
transform 1 0 27888 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_241
timestamp 1751532423
transform 1 0 28336 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_259
timestamp 1751532440
transform 1 0 30352 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_263
timestamp 1751532440
transform 1 0 30800 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_265
timestamp 1751532423
transform 1 0 31024 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_289
timestamp 1751532423
transform 1 0 33712 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_339
timestamp 1751532440
transform 1 0 39312 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_417
timestamp 1751532440
transform 1 0 48048 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_419
timestamp 1751532423
transform 1 0 48272 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_42_2
timestamp 1751532351
transform 1 0 1568 0 1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_42_18
timestamp 1751532351
transform 1 0 3360 0 1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_34
timestamp 1751532423
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_42_37
timestamp 1751532246
transform 1 0 5488 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_41
timestamp 1751532423
transform 1 0 5936 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_42_48
timestamp 1751532246
transform 1 0 6720 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_52
timestamp 1751532423
transform 1 0 7168 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_42_80
timestamp 1751532312
transform 1 0 10304 0 1 36064
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_107
timestamp 1751532440
transform 1 0 13328 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_42_111
timestamp 1751532246
transform 1 0 13776 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_115
timestamp 1751532440
transform 1 0 14224 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_117
timestamp 1751532423
transform 1 0 14448 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_42_124
timestamp 1751532246
transform 1 0 15232 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_128
timestamp 1751532440
transform 1 0 15680 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_130
timestamp 1751532423
transform 1 0 15904 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_171
timestamp 1751532440
transform 1 0 20496 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_42_177
timestamp 1751532246
transform 1 0 21168 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_183
timestamp 1751532440
transform 1 0 21840 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_187
timestamp 1751532423
transform 1 0 22288 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_243
timestamp 1751532440
transform 1 0 28560 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_247
timestamp 1751532440
transform 1 0 29008 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_251
timestamp 1751532423
transform 1 0 29456 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_285
timestamp 1751532440
transform 1 0 33264 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_287
timestamp 1751532423
transform 1 0 33488 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_323
timestamp 1751532440
transform 1 0 37520 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_327
timestamp 1751532440
transform 1 0 37968 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_331
timestamp 1751532440
transform 1 0 38416 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_333
timestamp 1751532423
transform 1 0 38640 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_384
timestamp 1751532423
transform 1 0 44352 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_394
timestamp 1751532423
transform 1 0 45472 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_2
timestamp 1751532351
transform 1 0 1568 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_18
timestamp 1751532351
transform 1 0 3360 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_43_34
timestamp 1751532246
transform 1 0 5152 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_38
timestamp 1751532440
transform 1 0 5600 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_47
timestamp 1751532351
transform 1 0 6608 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_67
timestamp 1751532440
transform 1 0 8848 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_69
timestamp 1751532423
transform 1 0 9072 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_76
timestamp 1751532440
transform 1 0 9856 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_78
timestamp 1751532423
transform 1 0 10080 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_43_112
timestamp 1751532312
transform 1 0 13888 0 -1 37632
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_43_120
timestamp 1751532246
transform 1 0 14784 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_124
timestamp 1751532440
transform 1 0 15232 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_126
timestamp 1751532423
transform 1 0 15456 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_133
timestamp 1751532440
transform 1 0 16240 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_135
timestamp 1751532423
transform 1 0 16464 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_156
timestamp 1751532440
transform 1 0 18816 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_173
timestamp 1751532423
transform 1 0 20720 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_207
timestamp 1751532440
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_209
timestamp 1751532423
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_43_212
timestamp 1751532246
transform 1 0 25088 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_216
timestamp 1751532423
transform 1 0 25536 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_233
timestamp 1751532440
transform 1 0 27440 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_237
timestamp 1751532440
transform 1 0 27888 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_239
timestamp 1751532423
transform 1 0 28112 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_255
timestamp 1751532440
transform 1 0 29904 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_43_267
timestamp 1751532246
transform 1 0 31248 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_271
timestamp 1751532423
transform 1 0 31696 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_282
timestamp 1751532440
transform 1 0 32928 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_308
timestamp 1751532440
transform 1 0 35840 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_312
timestamp 1751532423
transform 1 0 36288 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_340
timestamp 1751532440
transform 1 0 39424 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_43_344
timestamp 1751532246
transform 1 0 39872 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_388
timestamp 1751532423
transform 1 0 44800 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_393
timestamp 1751532440
transform 1 0 45360 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_395
timestamp 1751532423
transform 1 0 45584 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_422
timestamp 1751532423
transform 1 0 48608 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_2
timestamp 1751532351
transform 1 0 1568 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_18
timestamp 1751532351
transform 1 0 3360 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_34
timestamp 1751532423
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_44_85
timestamp 1751532246
transform 1 0 10864 0 1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_89
timestamp 1751532423
transform 1 0 11312 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_96
timestamp 1751532440
transform 1 0 12096 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_149
timestamp 1751532423
transform 1 0 18032 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_163
timestamp 1751532440
transform 1 0 19600 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_191
timestamp 1751532440
transform 1 0 22736 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_193
timestamp 1751532423
transform 1 0 22960 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_215
timestamp 1751532440
transform 1 0 25424 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_217
timestamp 1751532423
transform 1 0 25648 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_247
timestamp 1751532423
transform 1 0 29008 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_44_274
timestamp 1751532246
transform 1 0 32032 0 1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_278
timestamp 1751532440
transform 1 0 32480 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_288
timestamp 1751532440
transform 1 0 33600 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_292
timestamp 1751532440
transform 1 0 34048 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_294
timestamp 1751532423
transform 1 0 34272 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_323
timestamp 1751532440
transform 1 0 37520 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_352
timestamp 1751532440
transform 1 0 40768 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_354
timestamp 1751532423
transform 1 0 40992 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_362
timestamp 1751532423
transform 1 0 41888 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_384
timestamp 1751532423
transform 1 0 44352 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_394
timestamp 1751532440
transform 1 0 45472 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_45_2
timestamp 1751532312
transform 1 0 1568 0 -1 39200
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_45_10
timestamp 1751532246
transform 1 0 2464 0 -1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_14
timestamp 1751532440
transform 1 0 2912 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_16
timestamp 1751532423
transform 1 0 3136 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_58
timestamp 1751532440
transform 1 0 7840 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_60
timestamp 1751532423
transform 1 0 8064 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_97
timestamp 1751532423
transform 1 0 12208 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_45_109
timestamp 1751532312
transform 1 0 13552 0 -1 39200
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_131
timestamp 1751532440
transform 1 0 16016 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_142
timestamp 1751532440
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_180
timestamp 1751532440
transform 1 0 21504 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_182
timestamp 1751532423
transform 1 0 21728 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_197
timestamp 1751532440
transform 1 0 23408 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_206
timestamp 1751532440
transform 1 0 24416 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_237
timestamp 1751532440
transform 1 0 27888 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_239
timestamp 1751532423
transform 1 0 28112 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_268
timestamp 1751532423
transform 1 0 31360 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_326
timestamp 1751532423
transform 1 0 37856 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_333
timestamp 1751532440
transform 1 0 38640 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_45_337
timestamp 1751532312
transform 1 0 39088 0 -1 39200
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_45_345
timestamp 1751532246
transform 1 0 39984 0 -1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_349
timestamp 1751532423
transform 1 0 40432 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_379
timestamp 1751532423
transform 1 0 43792 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_418
timestamp 1751532440
transform 1 0 48160 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_428
timestamp 1751532423
transform 1 0 49280 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_46_2
timestamp 1751532351
transform 1 0 1568 0 1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_46_18
timestamp 1751532351
transform 1 0 3360 0 1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_34
timestamp 1751532423
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_80
timestamp 1751532440
transform 1 0 10304 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_82
timestamp 1751532423
transform 1 0 10528 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_93
timestamp 1751532423
transform 1 0 11760 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_46_107
timestamp 1751532246
transform 1 0 13328 0 1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_111
timestamp 1751532423
transform 1 0 13776 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_123
timestamp 1751532440
transform 1 0 15120 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_46_145
timestamp 1751532246
transform 1 0 17584 0 1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_149
timestamp 1751532423
transform 1 0 18032 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_173
timestamp 1751532440
transform 1 0 20720 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_202
timestamp 1751532440
transform 1 0 23968 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_46_219
timestamp 1751532246
transform 1 0 25872 0 1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_46_225
timestamp 1751532312
transform 1 0 26544 0 1 39200
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_233
timestamp 1751532423
transform 1 0 27440 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_244
timestamp 1751532423
transform 1 0 28672 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_247
timestamp 1751532440
transform 1 0 29008 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_283
timestamp 1751532440
transform 1 0 33040 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_287
timestamp 1751532440
transform 1 0 33488 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_291
timestamp 1751532440
transform 1 0 33936 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_293
timestamp 1751532423
transform 1 0 34160 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_303
timestamp 1751532423
transform 1 0 35280 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_310
timestamp 1751532440
transform 1 0 36064 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_312
timestamp 1751532423
transform 1 0 36288 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_46_355
timestamp 1751532246
transform 1 0 41104 0 1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_361
timestamp 1751532440
transform 1 0 41776 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_365
timestamp 1751532440
transform 1 0 42224 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_380
timestamp 1751532440
transform 1 0 43904 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_382
timestamp 1751532423
transform 1 0 44128 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_391
timestamp 1751532423
transform 1 0 45136 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_426
timestamp 1751532440
transform 1 0 49056 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_428
timestamp 1751532423
transform 1 0 49280 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_47_2
timestamp 1751532351
transform 1 0 1568 0 -1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_47_18
timestamp 1751532351
transform 1 0 3360 0 -1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_34
timestamp 1751532440
transform 1 0 5152 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_68
timestamp 1751532440
transform 1 0 8960 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_47_97
timestamp 1751532246
transform 1 0 12208 0 -1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_101
timestamp 1751532423
transform 1 0 12656 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_123
timestamp 1751532440
transform 1 0 15120 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_125
timestamp 1751532423
transform 1 0 15344 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_142
timestamp 1751532440
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_198
timestamp 1751532423
transform 1 0 23520 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_223
timestamp 1751532423
transform 1 0 26320 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_249
timestamp 1751532423
transform 1 0 29232 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_261
timestamp 1751532440
transform 1 0 30576 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_277
timestamp 1751532440
transform 1 0 32368 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_279
timestamp 1751532423
transform 1 0 32592 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_293
timestamp 1751532440
transform 1 0 34160 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_47_352
timestamp 1751532246
transform 1 0 40768 0 -1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_356
timestamp 1751532423
transform 1 0 41216 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_405
timestamp 1751532423
transform 1 0 46704 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_2
timestamp 1751532351
transform 1 0 1568 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_18
timestamp 1751532351
transform 1 0 3360 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_48_34
timestamp 1751532423
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_71
timestamp 1751532440
transform 1 0 9296 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_48_73
timestamp 1751532423
transform 1 0 9520 0 1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_89
timestamp 1751532440
transform 1 0 11312 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_128
timestamp 1751532440
transform 1 0 15680 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_147
timestamp 1751532440
transform 1 0 17808 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_48_151
timestamp 1751532312
transform 1 0 18256 0 1 40768
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_159
timestamp 1751532440
transform 1 0 19152 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_167
timestamp 1751532440
transform 1 0 20048 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_171
timestamp 1751532440
transform 1 0 20496 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_184
timestamp 1751532440
transform 1 0 21952 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_48_186
timestamp 1751532423
transform 1 0 22176 0 1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_48_244
timestamp 1751532423
transform 1 0 28672 0 1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_261
timestamp 1751532440
transform 1 0 30576 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_48_277
timestamp 1751532246
transform 1 0 32368 0 1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_281
timestamp 1751532440
transform 1 0 32816 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_310
timestamp 1751532440
transform 1 0 36064 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_48_312
timestamp 1751532423
transform 1 0 36288 0 1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_317
timestamp 1751532440
transform 1 0 36848 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_352
timestamp 1751532440
transform 1 0 40768 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_356
timestamp 1751532440
transform 1 0 41216 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_360
timestamp 1751532440
transform 1 0 41664 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_48_375
timestamp 1751532246
transform 1 0 43344 0 1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_48_401
timestamp 1751532423
transform 1 0 46256 0 1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_49_2
timestamp 1751532351
transform 1 0 1568 0 -1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_49_18
timestamp 1751532351
transform 1 0 3360 0 -1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_34
timestamp 1751532423
transform 1 0 5152 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_62
timestamp 1751532423
transform 1 0 8288 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_72
timestamp 1751532440
transform 1 0 9408 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_74
timestamp 1751532423
transform 1 0 9632 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_81
timestamp 1751532423
transform 1 0 10416 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_107
timestamp 1751532423
transform 1 0 13328 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_49_119
timestamp 1751532246
transform 1 0 14672 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_123
timestamp 1751532440
transform 1 0 15120 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_125
timestamp 1751532423
transform 1 0 15344 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_137
timestamp 1751532440
transform 1 0 16688 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_139
timestamp 1751532423
transform 1 0 16912 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_174
timestamp 1751532440
transform 1 0 20832 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_178
timestamp 1751532423
transform 1 0 21280 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_49_192
timestamp 1751532312
transform 1 0 22848 0 -1 42336
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_49_204
timestamp 1751532246
transform 1 0 24192 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_208
timestamp 1751532440
transform 1 0 24640 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_212
timestamp 1751532423
transform 1 0 25088 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_217
timestamp 1751532440
transform 1 0 25648 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_244
timestamp 1751532440
transform 1 0 28672 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_248
timestamp 1751532440
transform 1 0 29120 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_268
timestamp 1751532423
transform 1 0 31360 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_49_276
timestamp 1751532246
transform 1 0 32256 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_49_282
timestamp 1751532246
transform 1 0 32928 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_286
timestamp 1751532440
transform 1 0 33376 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_288
timestamp 1751532423
transform 1 0 33600 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_295
timestamp 1751532423
transform 1 0 34384 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_300
timestamp 1751532440
transform 1 0 34944 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_348
timestamp 1751532440
transform 1 0 40320 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_428
timestamp 1751532423
transform 1 0 49280 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_50_2
timestamp 1751532351
transform 1 0 1568 0 1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_50_18
timestamp 1751532351
transform 1 0 3360 0 1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_50_34
timestamp 1751532423
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_50_37
timestamp 1751532312
transform 1 0 5488 0 1 42336
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_50_45
timestamp 1751532246
transform 1 0 6384 0 1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_50_49
timestamp 1751532423
transform 1 0 6832 0 1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_50_64
timestamp 1751532440
transform 1 0 8512 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_50_93
timestamp 1751532423
transform 1 0 11760 0 1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_50_146
timestamp 1751532440
transform 1 0 17696 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_50_208
timestamp 1751532423
transform 1 0 24640 0 1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_50_229
timestamp 1751532440
transform 1 0 26992 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_50_242
timestamp 1751532440
transform 1 0 28448 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_50_244
timestamp 1751532423
transform 1 0 28672 0 1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_50_261
timestamp 1751532440
transform 1 0 30576 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_50_284
timestamp 1751532246
transform 1 0 33152 0 1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_50_288
timestamp 1751532440
transform 1 0 33600 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_50_340
timestamp 1751532440
transform 1 0 39424 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_50_373
timestamp 1751532423
transform 1 0 43120 0 1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_50_384
timestamp 1751532423
transform 1 0 44352 0 1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_50_387
timestamp 1751532423
transform 1 0 44688 0 1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_50_399
timestamp 1751532440
transform 1 0 46032 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_50_401
timestamp 1751532423
transform 1 0 46256 0 1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_51_2
timestamp 1751532351
transform 1 0 1568 0 -1 43904
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_51_18
timestamp 1751532351
transform 1 0 3360 0 -1 43904
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_51_34
timestamp 1751532312
transform 1 0 5152 0 -1 43904
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_51_42
timestamp 1751532423
transform 1 0 6048 0 -1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_51_78
timestamp 1751532440
transform 1 0 10080 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_51_105
timestamp 1751532423
transform 1 0 13104 0 -1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_51_173
timestamp 1751532440
transform 1 0 20720 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_51_177
timestamp 1751532423
transform 1 0 21168 0 -1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_51_212
timestamp 1751532423
transform 1 0 25088 0 -1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_51_251
timestamp 1751532440
transform 1 0 29456 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_51_277
timestamp 1751532440
transform 1 0 32368 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_51_279
timestamp 1751532423
transform 1 0 32592 0 -1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_51_292
timestamp 1751532440
transform 1 0 34048 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_51_312
timestamp 1751532440
transform 1 0 36288 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_51_341
timestamp 1751532440
transform 1 0 39536 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_51_343
timestamp 1751532423
transform 1 0 39760 0 -1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_51_368
timestamp 1751532440
transform 1 0 42560 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_51_370
timestamp 1751532423
transform 1 0 42784 0 -1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_51_403
timestamp 1751532440
transform 1 0 46480 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_51_418
timestamp 1751532440
transform 1 0 48160 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_51_428
timestamp 1751532423
transform 1 0 49280 0 -1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_52_2
timestamp 1751532351
transform 1 0 1568 0 1 43904
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_52_18
timestamp 1751532351
transform 1 0 3360 0 1 43904
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_52_34
timestamp 1751532423
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_52_37
timestamp 1751532351
transform 1 0 5488 0 1 43904
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_52_60
timestamp 1751532246
transform 1 0 8064 0 1 43904
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_52_64
timestamp 1751532440
transform 1 0 8512 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_52_66
timestamp 1751532423
transform 1 0 8736 0 1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_52_115
timestamp 1751532246
transform 1 0 14224 0 1 43904
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_52_119
timestamp 1751532440
transform 1 0 14672 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_52_152
timestamp 1751532440
transform 1 0 18368 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_52_173
timestamp 1751532440
transform 1 0 20720 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_52_177
timestamp 1751532423
transform 1 0 21168 0 1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_52_214
timestamp 1751532351
transform 1 0 25312 0 1 43904
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_52_230
timestamp 1751532440
transform 1 0 27104 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_52_254
timestamp 1751532440
transform 1 0 29792 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_52_285
timestamp 1751532423
transform 1 0 33264 0 1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_52_314
timestamp 1751532423
transform 1 0 36512 0 1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_52_364
timestamp 1751532440
transform 1 0 42112 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_52_408
timestamp 1751532423
transform 1 0 47040 0 1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_52_416
timestamp 1751532440
transform 1 0 47936 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_52_418
timestamp 1751532423
transform 1 0 48160 0 1 43904
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_53_2
timestamp 1751532351
transform 1 0 1568 0 -1 45472
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_53_18
timestamp 1751532351
transform 1 0 3360 0 -1 45472
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_53_34
timestamp 1751532351
transform 1 0 5152 0 -1 45472
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_53_50
timestamp 1751532351
transform 1 0 6944 0 -1 45472
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_53_66
timestamp 1751532246
transform 1 0 8736 0 -1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_53_99
timestamp 1751532440
transform 1 0 12432 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_53_103
timestamp 1751532440
transform 1 0 12880 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_53_130
timestamp 1751532246
transform 1 0 15904 0 -1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_53_134
timestamp 1751532440
transform 1 0 16352 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_53_149
timestamp 1751532440
transform 1 0 18032 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_53_151
timestamp 1751532423
transform 1 0 18256 0 -1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_53_179
timestamp 1751532423
transform 1 0 21392 0 -1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_53_207
timestamp 1751532440
transform 1 0 24528 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_53_209
timestamp 1751532423
transform 1 0 24752 0 -1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_53_246
timestamp 1751532246
transform 1 0 28896 0 -1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_53_250
timestamp 1751532423
transform 1 0 29344 0 -1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_53_253
timestamp 1751532246
transform 1 0 29680 0 -1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_53_257
timestamp 1751532440
transform 1 0 30128 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_53_259
timestamp 1751532423
transform 1 0 30352 0 -1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_53_278
timestamp 1751532440
transform 1 0 32480 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_53_309
timestamp 1751532423
transform 1 0 35952 0 -1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_53_338
timestamp 1751532440
transform 1 0 39200 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_53_342
timestamp 1751532440
transform 1 0 39648 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_53_346
timestamp 1751532440
transform 1 0 40096 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_53_406
timestamp 1751532440
transform 1 0 46816 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_53_408
timestamp 1751532423
transform 1 0 47040 0 -1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_54_2
timestamp 1751532351
transform 1 0 1568 0 1 45472
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_54_18
timestamp 1751532351
transform 1 0 3360 0 1 45472
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_54_34
timestamp 1751532423
transform 1 0 5152 0 1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_54_37
timestamp 1751532351
transform 1 0 5488 0 1 45472
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_54_53
timestamp 1751532351
transform 1 0 7280 0 1 45472
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_54_69
timestamp 1751532246
transform 1 0 9072 0 1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_54_83
timestamp 1751532440
transform 1 0 10640 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_54_103
timestamp 1751532440
transform 1 0 12880 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_54_177
timestamp 1751532423
transform 1 0 21168 0 1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_54_187
timestamp 1751532440
transform 1 0 22288 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_54_196
timestamp 1751532440
transform 1 0 23296 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_54_198
timestamp 1751532423
transform 1 0 23520 0 1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_54_226
timestamp 1751532246
transform 1 0 26656 0 1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_54_240
timestamp 1751532440
transform 1 0 28224 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_54_242
timestamp 1751532423
transform 1 0 28448 0 1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_54_254
timestamp 1751532440
transform 1 0 29792 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_54_308
timestamp 1751532246
transform 1 0 35840 0 1 45472
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_54_312
timestamp 1751532423
transform 1 0 36288 0 1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_54_344
timestamp 1751532440
transform 1 0 39872 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_54_346
timestamp 1751532423
transform 1 0 40096 0 1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_54_382
timestamp 1751532440
transform 1 0 44128 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_54_384
timestamp 1751532423
transform 1 0 44352 0 1 45472
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_55_2
timestamp 1751532351
transform 1 0 1568 0 -1 47040
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_55_18
timestamp 1751532351
transform 1 0 3360 0 -1 47040
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_55_34
timestamp 1751532351
transform 1 0 5152 0 -1 47040
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_55_50
timestamp 1751532351
transform 1 0 6944 0 -1 47040
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_55_66
timestamp 1751532246
transform 1 0 8736 0 -1 47040
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_55_72
timestamp 1751532246
transform 1 0 9408 0 -1 47040
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_55_76
timestamp 1751532440
transform 1 0 9856 0 -1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_55_78
timestamp 1751532423
transform 1 0 10080 0 -1 47040
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_55_146
timestamp 1751532312
transform 1 0 17696 0 -1 47040
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_55_154
timestamp 1751532246
transform 1 0 18592 0 -1 47040
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_55_158
timestamp 1751532440
transform 1 0 19040 0 -1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_55_160
timestamp 1751532423
transform 1 0 19264 0 -1 47040
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_55_167
timestamp 1751532423
transform 1 0 20048 0 -1 47040
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_55_209
timestamp 1751532423
transform 1 0 24752 0 -1 47040
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_55_226
timestamp 1751532246
transform 1 0 26656 0 -1 47040
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_55_230
timestamp 1751532440
transform 1 0 27104 0 -1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_55_273
timestamp 1751532423
transform 1 0 31920 0 -1 47040
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_55_340
timestamp 1751532440
transform 1 0 39424 0 -1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_55_342
timestamp 1751532423
transform 1 0 39648 0 -1 47040
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_55_352
timestamp 1751532440
transform 1 0 40768 0 -1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_55_364
timestamp 1751532440
transform 1 0 42112 0 -1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_55_428
timestamp 1751532423
transform 1 0 49280 0 -1 47040
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_56_2
timestamp 1751532351
transform 1 0 1568 0 1 47040
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_56_18
timestamp 1751532351
transform 1 0 3360 0 1 47040
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_56_36
timestamp 1751532351
transform 1 0 5376 0 1 47040
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_56_52
timestamp 1751532351
transform 1 0 7168 0 1 47040
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_56_70
timestamp 1751532351
transform 1 0 9184 0 1 47040
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_56_86
timestamp 1751532440
transform 1 0 10976 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_56_94
timestamp 1751532312
transform 1 0 11872 0 1 47040
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_56_104
timestamp 1751532423
transform 1 0 12992 0 1 47040
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_56_126
timestamp 1751532312
transform 1 0 15456 0 1 47040
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_56_134
timestamp 1751532440
transform 1 0 16352 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_56_138
timestamp 1751532351
transform 1 0 16800 0 1 47040
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_56_154
timestamp 1751532440
transform 1 0 18592 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_56_156
timestamp 1751532423
transform 1 0 18816 0 1 47040
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_56_165
timestamp 1751532246
transform 1 0 19824 0 1 47040
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_56_169
timestamp 1751532423
transform 1 0 20272 0 1 47040
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_56_172
timestamp 1751532440
transform 1 0 20608 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_56_176
timestamp 1751532423
transform 1 0 21056 0 1 47040
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_56_181
timestamp 1751532440
transform 1 0 21616 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_56_185
timestamp 1751532440
transform 1 0 22064 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_56_198
timestamp 1751532246
transform 1 0 23520 0 1 47040
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_56_202
timestamp 1751532440
transform 1 0 23968 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_56_213
timestamp 1751532312
transform 1 0 25200 0 1 47040
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_56_228
timestamp 1751532312
transform 1 0 26880 0 1 47040
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_56_236
timestamp 1751532440
transform 1 0 27776 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_56_254
timestamp 1751532440
transform 1 0 29792 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_56_256
timestamp 1751532423
transform 1 0 30016 0 1 47040
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_56_259
timestamp 1751532440
transform 1 0 30352 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_56_269
timestamp 1751532440
transform 1 0 31472 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_56_271
timestamp 1751532423
transform 1 0 31696 0 1 47040
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_56_315
timestamp 1751532440
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_56_319
timestamp 1751532440
transform 1 0 37072 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_56_327
timestamp 1751532440
transform 1 0 37968 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_56_331
timestamp 1751532440
transform 1 0 38416 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_56_333
timestamp 1751532423
transform 1 0 38640 0 1 47040
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_56_336
timestamp 1751532440
transform 1 0 38976 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_56_369
timestamp 1751532423
transform 1 0 42672 0 1 47040
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input1
timestamp 1751534193
transform -1 0 49392 0 -1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input2
timestamp 1751534193
transform -1 0 47376 0 -1 43904
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_4  input3 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751546029
transform -1 0 49392 0 1 47040
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input4
timestamp 1751534193
transform -1 0 49392 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input5
timestamp 1751534193
transform -1 0 49392 0 1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input6
timestamp 1751534193
transform -1 0 49392 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input7
timestamp 1751534193
transform -1 0 49392 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input8
timestamp 1751534193
transform 1 0 32032 0 -1 47040
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input9
timestamp 1751534193
transform 1 0 47264 0 1 47040
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input10
timestamp 1751534193
transform 1 0 19152 0 1 47040
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output11
timestamp 1751661108
transform 1 0 19152 0 -1 6272
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output12
timestamp 1751661108
transform 1 0 20944 0 1 3136
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output13
timestamp 1751661108
transform -1 0 34832 0 1 3136
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output14
timestamp 1751661108
transform 1 0 35840 0 1 3136
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output15
timestamp 1751661108
transform -1 0 38080 0 -1 6272
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output16
timestamp 1751661108
transform -1 0 42448 0 1 3136
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output17
timestamp 1751661108
transform 1 0 41552 0 1 4704
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output18
timestamp 1751661108
transform 1 0 13776 0 1 3136
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output19
timestamp 1751661108
transform 1 0 17360 0 1 4704
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_0_Left_57 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532504
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_0_Right_0
timestamp 1751532504
transform -1 0 49616 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_1_Left_58
timestamp 1751532504
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_1_Right_1
timestamp 1751532504
transform -1 0 49616 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_2_Left_59
timestamp 1751532504
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_2_Right_2
timestamp 1751532504
transform -1 0 49616 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_3_Left_60
timestamp 1751532504
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_3_Right_3
timestamp 1751532504
transform -1 0 49616 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_4_Left_61
timestamp 1751532504
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_4_Right_4
timestamp 1751532504
transform -1 0 49616 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_5_Left_62
timestamp 1751532504
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_5_Right_5
timestamp 1751532504
transform -1 0 49616 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_6_Left_63
timestamp 1751532504
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_6_Right_6
timestamp 1751532504
transform -1 0 49616 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_7_Left_64
timestamp 1751532504
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_7_Right_7
timestamp 1751532504
transform -1 0 49616 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_8_Left_65
timestamp 1751532504
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_8_Right_8
timestamp 1751532504
transform -1 0 49616 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_9_Left_66
timestamp 1751532504
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_9_Right_9
timestamp 1751532504
transform -1 0 49616 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_10_Left_67
timestamp 1751532504
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_10_Right_10
timestamp 1751532504
transform -1 0 49616 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_11_Left_68
timestamp 1751532504
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_11_Right_11
timestamp 1751532504
transform -1 0 49616 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_12_Left_69
timestamp 1751532504
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_12_Right_12
timestamp 1751532504
transform -1 0 49616 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_13_Left_70
timestamp 1751532504
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_13_Right_13
timestamp 1751532504
transform -1 0 49616 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_14_Left_71
timestamp 1751532504
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_14_Right_14
timestamp 1751532504
transform -1 0 49616 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_15_Left_72
timestamp 1751532504
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_15_Right_15
timestamp 1751532504
transform -1 0 49616 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_16_Left_73
timestamp 1751532504
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_16_Right_16
timestamp 1751532504
transform -1 0 49616 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_17_Left_74
timestamp 1751532504
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_17_Right_17
timestamp 1751532504
transform -1 0 49616 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_18_Left_75
timestamp 1751532504
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_18_Right_18
timestamp 1751532504
transform -1 0 49616 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_19_Left_76
timestamp 1751532504
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_19_Right_19
timestamp 1751532504
transform -1 0 49616 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_20_Left_77
timestamp 1751532504
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_20_Right_20
timestamp 1751532504
transform -1 0 49616 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_21_Left_78
timestamp 1751532504
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_21_Right_21
timestamp 1751532504
transform -1 0 49616 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_22_Left_79
timestamp 1751532504
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_22_Right_22
timestamp 1751532504
transform -1 0 49616 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_23_Left_80
timestamp 1751532504
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_23_Right_23
timestamp 1751532504
transform -1 0 49616 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_24_Left_81
timestamp 1751532504
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_24_Right_24
timestamp 1751532504
transform -1 0 49616 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_25_Left_82
timestamp 1751532504
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_25_Right_25
timestamp 1751532504
transform -1 0 49616 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_26_Left_83
timestamp 1751532504
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_26_Right_26
timestamp 1751532504
transform -1 0 49616 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_27_Left_84
timestamp 1751532504
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_27_Right_27
timestamp 1751532504
transform -1 0 49616 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_28_Left_85
timestamp 1751532504
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_28_Right_28
timestamp 1751532504
transform -1 0 49616 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_29_Left_86
timestamp 1751532504
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_29_Right_29
timestamp 1751532504
transform -1 0 49616 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_30_Left_87
timestamp 1751532504
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_30_Right_30
timestamp 1751532504
transform -1 0 49616 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_31_Left_88
timestamp 1751532504
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_31_Right_31
timestamp 1751532504
transform -1 0 49616 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_32_Left_89
timestamp 1751532504
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_32_Right_32
timestamp 1751532504
transform -1 0 49616 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_33_Left_90
timestamp 1751532504
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_33_Right_33
timestamp 1751532504
transform -1 0 49616 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_34_Left_91
timestamp 1751532504
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_34_Right_34
timestamp 1751532504
transform -1 0 49616 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_35_Left_92
timestamp 1751532504
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_35_Right_35
timestamp 1751532504
transform -1 0 49616 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_36_Left_93
timestamp 1751532504
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_36_Right_36
timestamp 1751532504
transform -1 0 49616 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_37_Left_94
timestamp 1751532504
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_37_Right_37
timestamp 1751532504
transform -1 0 49616 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_38_Left_95
timestamp 1751532504
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_38_Right_38
timestamp 1751532504
transform -1 0 49616 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_39_Left_96
timestamp 1751532504
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_39_Right_39
timestamp 1751532504
transform -1 0 49616 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_40_Left_97
timestamp 1751532504
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_40_Right_40
timestamp 1751532504
transform -1 0 49616 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_41_Left_98
timestamp 1751532504
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_41_Right_41
timestamp 1751532504
transform -1 0 49616 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_42_Left_99
timestamp 1751532504
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_42_Right_42
timestamp 1751532504
transform -1 0 49616 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_43_Left_100
timestamp 1751532504
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_43_Right_43
timestamp 1751532504
transform -1 0 49616 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_44_Left_101
timestamp 1751532504
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_44_Right_44
timestamp 1751532504
transform -1 0 49616 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_45_Left_102
timestamp 1751532504
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_45_Right_45
timestamp 1751532504
transform -1 0 49616 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_46_Left_103
timestamp 1751532504
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_46_Right_46
timestamp 1751532504
transform -1 0 49616 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_47_Left_104
timestamp 1751532504
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_47_Right_47
timestamp 1751532504
transform -1 0 49616 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_48_Left_105
timestamp 1751532504
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_48_Right_48
timestamp 1751532504
transform -1 0 49616 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_49_Left_106
timestamp 1751532504
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_49_Right_49
timestamp 1751532504
transform -1 0 49616 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_50_Left_107
timestamp 1751532504
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_50_Right_50
timestamp 1751532504
transform -1 0 49616 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_51_Left_108
timestamp 1751532504
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_51_Right_51
timestamp 1751532504
transform -1 0 49616 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_52_Left_109
timestamp 1751532504
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_52_Right_52
timestamp 1751532504
transform -1 0 49616 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_53_Left_110
timestamp 1751532504
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_53_Right_53
timestamp 1751532504
transform -1 0 49616 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_54_Left_111
timestamp 1751532504
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_54_Right_54
timestamp 1751532504
transform -1 0 49616 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_55_Left_112
timestamp 1751532504
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_55_Right_55
timestamp 1751532504
transform -1 0 49616 0 -1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_56_Left_113
timestamp 1751532504
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_56_Right_56
timestamp 1751532504
transform -1 0 49616 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_114
timestamp 1751532504
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_115
timestamp 1751532504
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_116
timestamp 1751532504
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_117
timestamp 1751532504
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_118
timestamp 1751532504
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_119
timestamp 1751532504
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_120
timestamp 1751532504
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_121
timestamp 1751532504
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_122
timestamp 1751532504
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_123
timestamp 1751532504
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_124
timestamp 1751532504
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_125
timestamp 1751532504
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_126
timestamp 1751532504
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_127
timestamp 1751532504
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_128
timestamp 1751532504
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_129
timestamp 1751532504
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_130
timestamp 1751532504
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_131
timestamp 1751532504
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_132
timestamp 1751532504
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_133
timestamp 1751532504
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_134
timestamp 1751532504
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_135
timestamp 1751532504
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_136
timestamp 1751532504
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_137
timestamp 1751532504
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_138
timestamp 1751532504
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_139
timestamp 1751532504
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_140
timestamp 1751532504
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_141
timestamp 1751532504
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_142
timestamp 1751532504
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_143
timestamp 1751532504
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_144
timestamp 1751532504
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_145
timestamp 1751532504
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_146
timestamp 1751532504
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_147
timestamp 1751532504
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_148
timestamp 1751532504
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_149
timestamp 1751532504
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_150
timestamp 1751532504
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_151
timestamp 1751532504
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_152
timestamp 1751532504
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_153
timestamp 1751532504
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_154
timestamp 1751532504
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_155
timestamp 1751532504
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_156
timestamp 1751532504
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_157
timestamp 1751532504
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_158
timestamp 1751532504
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_159
timestamp 1751532504
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_160
timestamp 1751532504
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_161
timestamp 1751532504
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_162
timestamp 1751532504
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_163
timestamp 1751532504
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_164
timestamp 1751532504
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_165
timestamp 1751532504
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_166
timestamp 1751532504
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_167
timestamp 1751532504
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_168
timestamp 1751532504
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_169
timestamp 1751532504
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_170
timestamp 1751532504
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_171
timestamp 1751532504
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_172
timestamp 1751532504
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_173
timestamp 1751532504
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_174
timestamp 1751532504
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_175
timestamp 1751532504
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_176
timestamp 1751532504
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_177
timestamp 1751532504
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_178
timestamp 1751532504
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_179
timestamp 1751532504
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_180
timestamp 1751532504
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_181
timestamp 1751532504
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_182
timestamp 1751532504
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_183
timestamp 1751532504
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_184
timestamp 1751532504
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_185
timestamp 1751532504
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_186
timestamp 1751532504
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_187
timestamp 1751532504
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_188
timestamp 1751532504
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_189
timestamp 1751532504
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_190
timestamp 1751532504
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_191
timestamp 1751532504
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_192
timestamp 1751532504
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_193
timestamp 1751532504
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_194
timestamp 1751532504
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_195
timestamp 1751532504
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_196
timestamp 1751532504
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_197
timestamp 1751532504
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_198
timestamp 1751532504
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_199
timestamp 1751532504
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_200
timestamp 1751532504
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_201
timestamp 1751532504
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_202
timestamp 1751532504
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_203
timestamp 1751532504
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_204
timestamp 1751532504
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_205
timestamp 1751532504
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_206
timestamp 1751532504
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_207
timestamp 1751532504
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_208
timestamp 1751532504
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_209
timestamp 1751532504
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_210
timestamp 1751532504
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_211
timestamp 1751532504
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_212
timestamp 1751532504
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_213
timestamp 1751532504
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_214
timestamp 1751532504
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_215
timestamp 1751532504
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_216
timestamp 1751532504
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_217
timestamp 1751532504
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_218
timestamp 1751532504
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_219
timestamp 1751532504
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_220
timestamp 1751532504
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_221
timestamp 1751532504
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_222
timestamp 1751532504
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_223
timestamp 1751532504
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_224
timestamp 1751532504
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_225
timestamp 1751532504
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_226
timestamp 1751532504
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_227
timestamp 1751532504
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_228
timestamp 1751532504
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_229
timestamp 1751532504
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_230
timestamp 1751532504
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_231
timestamp 1751532504
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_232
timestamp 1751532504
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_233
timestamp 1751532504
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_234
timestamp 1751532504
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_235
timestamp 1751532504
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_236
timestamp 1751532504
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_237
timestamp 1751532504
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_238
timestamp 1751532504
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_239
timestamp 1751532504
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_240
timestamp 1751532504
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_241
timestamp 1751532504
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_242
timestamp 1751532504
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_243
timestamp 1751532504
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_244
timestamp 1751532504
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_245
timestamp 1751532504
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_246
timestamp 1751532504
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_247
timestamp 1751532504
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_248
timestamp 1751532504
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_249
timestamp 1751532504
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_250
timestamp 1751532504
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_251
timestamp 1751532504
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_252
timestamp 1751532504
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_253
timestamp 1751532504
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_254
timestamp 1751532504
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_255
timestamp 1751532504
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_256
timestamp 1751532504
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_257
timestamp 1751532504
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_258
timestamp 1751532504
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_259
timestamp 1751532504
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_260
timestamp 1751532504
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_261
timestamp 1751532504
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_262
timestamp 1751532504
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_263
timestamp 1751532504
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_264
timestamp 1751532504
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_265
timestamp 1751532504
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_266
timestamp 1751532504
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_267
timestamp 1751532504
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_268
timestamp 1751532504
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_269
timestamp 1751532504
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_270
timestamp 1751532504
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_271
timestamp 1751532504
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_272
timestamp 1751532504
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_273
timestamp 1751532504
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_274
timestamp 1751532504
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_275
timestamp 1751532504
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_276
timestamp 1751532504
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_277
timestamp 1751532504
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_278
timestamp 1751532504
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_279
timestamp 1751532504
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_280
timestamp 1751532504
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_281
timestamp 1751532504
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_282
timestamp 1751532504
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_283
timestamp 1751532504
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_284
timestamp 1751532504
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_285
timestamp 1751532504
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_286
timestamp 1751532504
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_287
timestamp 1751532504
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_288
timestamp 1751532504
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_289
timestamp 1751532504
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_290
timestamp 1751532504
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_291
timestamp 1751532504
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_292
timestamp 1751532504
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_293
timestamp 1751532504
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_294
timestamp 1751532504
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_295
timestamp 1751532504
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_296
timestamp 1751532504
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_297
timestamp 1751532504
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_298
timestamp 1751532504
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_299
timestamp 1751532504
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_300
timestamp 1751532504
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_301
timestamp 1751532504
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_302
timestamp 1751532504
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_303
timestamp 1751532504
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_304
timestamp 1751532504
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_305
timestamp 1751532504
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_306
timestamp 1751532504
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_307
timestamp 1751532504
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_308
timestamp 1751532504
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_309
timestamp 1751532504
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_310
timestamp 1751532504
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_311
timestamp 1751532504
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_312
timestamp 1751532504
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_313
timestamp 1751532504
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_314
timestamp 1751532504
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_315
timestamp 1751532504
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_316
timestamp 1751532504
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_317
timestamp 1751532504
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_318
timestamp 1751532504
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_319
timestamp 1751532504
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_320
timestamp 1751532504
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_321
timestamp 1751532504
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_322
timestamp 1751532504
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_323
timestamp 1751532504
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_324
timestamp 1751532504
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_325
timestamp 1751532504
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_326
timestamp 1751532504
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_327
timestamp 1751532504
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_328
timestamp 1751532504
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_329
timestamp 1751532504
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_330
timestamp 1751532504
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_331
timestamp 1751532504
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_332
timestamp 1751532504
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_333
timestamp 1751532504
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_334
timestamp 1751532504
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_335
timestamp 1751532504
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_336
timestamp 1751532504
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_337
timestamp 1751532504
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_338
timestamp 1751532504
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_339
timestamp 1751532504
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_340
timestamp 1751532504
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_341
timestamp 1751532504
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_342
timestamp 1751532504
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_343
timestamp 1751532504
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_344
timestamp 1751532504
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_345
timestamp 1751532504
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_346
timestamp 1751532504
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_347
timestamp 1751532504
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_348
timestamp 1751532504
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_349
timestamp 1751532504
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_350
timestamp 1751532504
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_351
timestamp 1751532504
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_352
timestamp 1751532504
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_353
timestamp 1751532504
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_354
timestamp 1751532504
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_355
timestamp 1751532504
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_356
timestamp 1751532504
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_357
timestamp 1751532504
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_358
timestamp 1751532504
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_359
timestamp 1751532504
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_360
timestamp 1751532504
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_361
timestamp 1751532504
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_362
timestamp 1751532504
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_363
timestamp 1751532504
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_364
timestamp 1751532504
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_365
timestamp 1751532504
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_366
timestamp 1751532504
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_367
timestamp 1751532504
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_368
timestamp 1751532504
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_369
timestamp 1751532504
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_370
timestamp 1751532504
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_371
timestamp 1751532504
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_372
timestamp 1751532504
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_373
timestamp 1751532504
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_374
timestamp 1751532504
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_375
timestamp 1751532504
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_376
timestamp 1751532504
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_377
timestamp 1751532504
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_43_378
timestamp 1751532504
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_43_379
timestamp 1751532504
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_43_380
timestamp 1751532504
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_43_381
timestamp 1751532504
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_43_382
timestamp 1751532504
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_43_383
timestamp 1751532504
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_44_384
timestamp 1751532504
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_44_385
timestamp 1751532504
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_44_386
timestamp 1751532504
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_44_387
timestamp 1751532504
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_44_388
timestamp 1751532504
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_44_389
timestamp 1751532504
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_45_390
timestamp 1751532504
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_45_391
timestamp 1751532504
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_45_392
timestamp 1751532504
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_45_393
timestamp 1751532504
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_45_394
timestamp 1751532504
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_45_395
timestamp 1751532504
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_46_396
timestamp 1751532504
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_46_397
timestamp 1751532504
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_46_398
timestamp 1751532504
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_46_399
timestamp 1751532504
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_46_400
timestamp 1751532504
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_46_401
timestamp 1751532504
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_47_402
timestamp 1751532504
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_47_403
timestamp 1751532504
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_47_404
timestamp 1751532504
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_47_405
timestamp 1751532504
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_47_406
timestamp 1751532504
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_47_407
timestamp 1751532504
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_48_408
timestamp 1751532504
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_48_409
timestamp 1751532504
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_48_410
timestamp 1751532504
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_48_411
timestamp 1751532504
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_48_412
timestamp 1751532504
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_48_413
timestamp 1751532504
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_414
timestamp 1751532504
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_415
timestamp 1751532504
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_416
timestamp 1751532504
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_417
timestamp 1751532504
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_418
timestamp 1751532504
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_419
timestamp 1751532504
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_50_420
timestamp 1751532504
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_50_421
timestamp 1751532504
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_50_422
timestamp 1751532504
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_50_423
timestamp 1751532504
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_50_424
timestamp 1751532504
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_50_425
timestamp 1751532504
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_51_426
timestamp 1751532504
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_51_427
timestamp 1751532504
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_51_428
timestamp 1751532504
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_51_429
timestamp 1751532504
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_51_430
timestamp 1751532504
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_51_431
timestamp 1751532504
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_52_432
timestamp 1751532504
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_52_433
timestamp 1751532504
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_52_434
timestamp 1751532504
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_52_435
timestamp 1751532504
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_52_436
timestamp 1751532504
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_52_437
timestamp 1751532504
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_53_438
timestamp 1751532504
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_53_439
timestamp 1751532504
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_53_440
timestamp 1751532504
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_53_441
timestamp 1751532504
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_53_442
timestamp 1751532504
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_53_443
timestamp 1751532504
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_54_444
timestamp 1751532504
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_54_445
timestamp 1751532504
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_54_446
timestamp 1751532504
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_54_447
timestamp 1751532504
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_54_448
timestamp 1751532504
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_54_449
timestamp 1751532504
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_55_450
timestamp 1751532504
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_55_451
timestamp 1751532504
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_55_452
timestamp 1751532504
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_55_453
timestamp 1751532504
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_55_454
timestamp 1751532504
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_55_455
timestamp 1751532504
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_56_456
timestamp 1751532504
transform 1 0 5152 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_56_457
timestamp 1751532504
transform 1 0 8960 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_56_458
timestamp 1751532504
transform 1 0 12768 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_56_459
timestamp 1751532504
transform 1 0 16576 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_56_460
timestamp 1751532504
transform 1 0 20384 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_56_461
timestamp 1751532504
transform 1 0 24192 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_56_462
timestamp 1751532504
transform 1 0 28000 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_56_463
timestamp 1751532504
transform 1 0 31808 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_56_464
timestamp 1751532504
transform 1 0 35616 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_56_465
timestamp 1751532504
transform 1 0 39424 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_56_466
timestamp 1751532504
transform 1 0 43232 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_56_467
timestamp 1751532504
transform 1 0 47040 0 1 47040
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_ay8913_20 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532612
transform 1 0 1568 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_ay8913_21
timestamp 1751532612
transform 1 0 3024 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_ay8913_22
timestamp 1751532612
transform 1 0 5376 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_ay8913_23
timestamp 1751532612
transform 1 0 6608 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_ay8913_24
timestamp 1751532612
transform 1 0 8400 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_ay8913_25
timestamp 1751532612
transform 1 0 10192 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_ay8913_26
timestamp 1751532612
transform 1 0 11984 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_ay8913_27
timestamp 1751532612
transform -1 0 13776 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_ay8913_28
timestamp 1751532612
transform -1 0 20384 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_ay8913_29
timestamp 1751532612
transform -1 0 24192 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_ay8913_30
timestamp 1751532612
transform 1 0 26432 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_ay8913_31
timestamp 1751532612
transform 1 0 28224 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_ay8913_32
timestamp 1751532612
transform -1 0 28000 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_ay8913_33
timestamp 1751532612
transform 1 0 45920 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_ay8913_34
timestamp 1751532612
transform 1 0 48944 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_ay8913_35
timestamp 1751532612
transform -1 0 44464 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_ay8913_36
timestamp 1751532612
transform 1 0 47936 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_ay8913_37
timestamp 1751532612
transform -1 0 49392 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__tiel_4  wrapped_ay8913_38
timestamp 1751532612
transform 1 0 40768 0 -1 4704
box -86 -86 534 870
<< labels >>
flabel metal3 s 50200 36064 51000 36176 0 FreeSans 448 0 0 0 custom_settings[0]
port 0 nsew signal input
flabel metal3 s 50200 40320 51000 40432 0 FreeSans 448 0 0 0 custom_settings[1]
port 1 nsew signal input
flabel metal3 s 50200 44576 51000 44688 0 FreeSans 448 0 0 0 custom_settings[2]
port 2 nsew signal input
flabel metal3 s 50200 48832 51000 48944 0 FreeSans 448 0 0 0 custom_settings[3]
port 3 nsew signal input
flabel metal3 s 50200 2016 51000 2128 0 FreeSans 448 0 0 0 io_in_1[0]
port 4 nsew signal input
flabel metal3 s 50200 6272 51000 6384 0 FreeSans 448 0 0 0 io_in_1[1]
port 5 nsew signal input
flabel metal3 s 50200 10528 51000 10640 0 FreeSans 448 0 0 0 io_in_1[2]
port 6 nsew signal input
flabel metal3 s 50200 14784 51000 14896 0 FreeSans 448 0 0 0 io_in_1[3]
port 7 nsew signal input
flabel metal3 s 50200 19040 51000 19152 0 FreeSans 448 0 0 0 io_in_1[4]
port 8 nsew signal input
flabel metal3 s 50200 23296 51000 23408 0 FreeSans 448 0 0 0 io_in_1[5]
port 9 nsew signal input
flabel metal3 s 50200 27552 51000 27664 0 FreeSans 448 0 0 0 io_in_1[6]
port 10 nsew signal input
flabel metal3 s 50200 31808 51000 31920 0 FreeSans 448 0 0 0 io_in_1[7]
port 11 nsew signal input
flabel metal2 s 31808 50200 31920 51000 0 FreeSans 448 90 0 0 io_in_2[0]
port 12 nsew signal input
flabel metal2 s 44576 50200 44688 51000 0 FreeSans 448 90 0 0 io_in_2[1]
port 13 nsew signal input
flabel metal2 s 1120 0 1232 800 0 FreeSans 448 90 0 0 io_out[0]
port 14 nsew signal output
flabel metal2 s 19040 0 19152 800 0 FreeSans 448 90 0 0 io_out[10]
port 15 nsew signal output
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 io_out[11]
port 16 nsew signal output
flabel metal2 s 22624 0 22736 800 0 FreeSans 448 90 0 0 io_out[12]
port 17 nsew signal output
flabel metal2 s 24416 0 24528 800 0 FreeSans 448 90 0 0 io_out[13]
port 18 nsew signal output
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 io_out[14]
port 19 nsew signal output
flabel metal2 s 28000 0 28112 800 0 FreeSans 448 90 0 0 io_out[15]
port 20 nsew signal output
flabel metal2 s 29792 0 29904 800 0 FreeSans 448 90 0 0 io_out[16]
port 21 nsew signal output
flabel metal2 s 31584 0 31696 800 0 FreeSans 448 90 0 0 io_out[17]
port 22 nsew signal output
flabel metal2 s 33376 0 33488 800 0 FreeSans 448 90 0 0 io_out[18]
port 23 nsew signal output
flabel metal2 s 35168 0 35280 800 0 FreeSans 448 90 0 0 io_out[19]
port 24 nsew signal output
flabel metal2 s 2912 0 3024 800 0 FreeSans 448 90 0 0 io_out[1]
port 25 nsew signal output
flabel metal2 s 36960 0 37072 800 0 FreeSans 448 90 0 0 io_out[20]
port 26 nsew signal output
flabel metal2 s 38752 0 38864 800 0 FreeSans 448 90 0 0 io_out[21]
port 27 nsew signal output
flabel metal2 s 40544 0 40656 800 0 FreeSans 448 90 0 0 io_out[22]
port 28 nsew signal output
flabel metal2 s 42336 0 42448 800 0 FreeSans 448 90 0 0 io_out[23]
port 29 nsew signal output
flabel metal2 s 44128 0 44240 800 0 FreeSans 448 90 0 0 io_out[24]
port 30 nsew signal output
flabel metal2 s 45920 0 46032 800 0 FreeSans 448 90 0 0 io_out[25]
port 31 nsew signal output
flabel metal2 s 47712 0 47824 800 0 FreeSans 448 90 0 0 io_out[26]
port 32 nsew signal output
flabel metal2 s 49504 0 49616 800 0 FreeSans 448 90 0 0 io_out[27]
port 33 nsew signal output
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 io_out[2]
port 34 nsew signal output
flabel metal2 s 6496 0 6608 800 0 FreeSans 448 90 0 0 io_out[3]
port 35 nsew signal output
flabel metal2 s 8288 0 8400 800 0 FreeSans 448 90 0 0 io_out[4]
port 36 nsew signal output
flabel metal2 s 10080 0 10192 800 0 FreeSans 448 90 0 0 io_out[5]
port 37 nsew signal output
flabel metal2 s 11872 0 11984 800 0 FreeSans 448 90 0 0 io_out[6]
port 38 nsew signal output
flabel metal2 s 13664 0 13776 800 0 FreeSans 448 90 0 0 io_out[7]
port 39 nsew signal output
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 io_out[8]
port 40 nsew signal output
flabel metal2 s 17248 0 17360 800 0 FreeSans 448 90 0 0 io_out[9]
port 41 nsew signal output
flabel metal2 s 19040 50200 19152 51000 0 FreeSans 448 90 0 0 rst_n
port 42 nsew signal input
flabel metal4 s 4448 3076 4768 47884 0 FreeSans 1280 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 35168 3076 35488 47884 0 FreeSans 1280 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 19808 3076 20128 47884 0 FreeSans 1280 90 0 0 vss
port 44 nsew ground bidirectional
flabel metal2 s 6272 50200 6384 51000 0 FreeSans 448 90 0 0 wb_clk_i
port 45 nsew signal input
rlabel metal1 25480 47824 25480 47824 0 vdd
rlabel metal1 25480 47040 25480 47040 0 vss
rlabel metal2 2744 28896 2744 28896 0 _0000_
rlabel metal2 2464 30408 2464 30408 0 _0001_
rlabel metal2 7560 32256 7560 32256 0 _0002_
rlabel metal2 3640 31892 3640 31892 0 _0003_
rlabel metal2 4872 28280 4872 28280 0 _0004_
rlabel metal2 2352 27160 2352 27160 0 _0005_
rlabel metal2 7336 24808 7336 24808 0 _0006_
rlabel metal2 2408 23632 2408 23632 0 _0007_
rlabel metal2 3752 25872 3752 25872 0 _0008_
rlabel metal2 2072 21224 2072 21224 0 _0009_
rlabel metal2 2072 19656 2072 19656 0 _0010_
rlabel metal2 6664 22736 6664 22736 0 _0011_
rlabel metal2 8120 18704 8120 18704 0 _0012_
rlabel metal2 2408 17976 2408 17976 0 _0013_
rlabel metal2 2464 16296 2464 16296 0 _0014_
rlabel metal2 2408 14840 2408 14840 0 _0015_
rlabel metal2 10472 16408 10472 16408 0 _0016_
rlabel metal3 8008 14616 8008 14616 0 _0017_
rlabel metal2 3416 13384 3416 13384 0 _0018_
rlabel metal2 9240 13272 9240 13272 0 _0019_
rlabel metal2 11928 14000 11928 14000 0 _0020_
rlabel metal2 12880 8344 12880 8344 0 _0021_
rlabel metal2 9352 11088 9352 11088 0 _0022_
rlabel metal2 2408 11816 2408 11816 0 _0023_
rlabel metal2 2408 10248 2408 10248 0 _0024_
rlabel metal3 3696 8344 3696 8344 0 _0025_
rlabel metal2 2464 6888 2464 6888 0 _0026_
rlabel metal2 3080 5432 3080 5432 0 _0027_
rlabel metal2 8344 4760 8344 4760 0 _0028_
rlabel metal2 8232 7896 8232 7896 0 _0029_
rlabel metal2 11480 6272 11480 6272 0 _0030_
rlabel metal2 11592 9324 11592 9324 0 _0031_
rlabel metal2 15736 22680 15736 22680 0 _0032_
rlabel metal2 9912 22064 9912 22064 0 _0033_
rlabel metal2 13272 21896 13272 21896 0 _0034_
rlabel metal2 10136 21112 10136 21112 0 _0035_
rlabel metal3 22344 21560 22344 21560 0 _0036_
rlabel metal2 7784 33656 7784 33656 0 _0037_
rlabel metal2 8120 36176 8120 36176 0 _0038_
rlabel metal3 6104 34104 6104 34104 0 _0039_
rlabel metal2 5992 35784 5992 35784 0 _0040_
rlabel metal3 38472 4312 38472 4312 0 _0041_
rlabel metal2 39144 6384 39144 6384 0 _0042_
rlabel metal2 37128 8456 37128 8456 0 _0043_
rlabel metal2 40152 11704 40152 11704 0 _0044_
rlabel metal2 36792 12432 36792 12432 0 _0045_
rlabel metal2 35336 9296 35336 9296 0 _0046_
rlabel metal2 35112 6216 35112 6216 0 _0047_
rlabel metal2 31192 3752 31192 3752 0 _0048_
rlabel metal2 31528 5656 31528 5656 0 _0049_
rlabel metal2 41608 9296 41608 9296 0 _0050_
rlabel metal2 41160 8792 41160 8792 0 _0051_
rlabel metal3 42280 3752 42280 3752 0 _0052_
rlabel metal2 42168 4928 42168 4928 0 _0053_
rlabel metal3 47432 3752 47432 3752 0 _0054_
rlabel metal2 49000 3976 49000 3976 0 _0055_
rlabel metal2 49000 14056 49000 14056 0 _0056_
rlabel metal2 49000 5600 49000 5600 0 _0057_
rlabel metal2 47768 5320 47768 5320 0 _0058_
rlabel metal2 47432 10136 47432 10136 0 _0059_
rlabel metal2 30296 8792 30296 8792 0 _0060_
rlabel metal3 28616 5880 28616 5880 0 _0061_
rlabel metal2 27664 4312 27664 4312 0 _0062_
rlabel metal2 14728 3864 14728 3864 0 _0063_
rlabel metal2 14840 5432 14840 5432 0 _0064_
rlabel metal2 14840 8008 14840 8008 0 _0065_
rlabel metal2 18424 7728 18424 7728 0 _0066_
rlabel metal2 20440 4592 20440 4592 0 _0067_
rlabel metal2 32648 14784 32648 14784 0 _0068_
rlabel metal2 28616 15316 28616 15316 0 _0069_
rlabel metal2 27888 13160 27888 13160 0 _0070_
rlabel metal2 26600 11088 26600 11088 0 _0071_
rlabel metal2 26824 9296 26824 9296 0 _0072_
rlabel metal2 25928 7728 25928 7728 0 _0073_
rlabel metal2 23128 6944 23128 6944 0 _0074_
rlabel metal2 24528 4536 24528 4536 0 _0075_
rlabel metal2 14280 36176 14280 36176 0 _0076_
rlabel metal2 19432 35896 19432 35896 0 _0077_
rlabel metal2 11368 36680 11368 36680 0 _0078_
rlabel metal3 11592 34328 11592 34328 0 _0079_
rlabel metal2 19656 40656 19656 40656 0 _0080_
rlabel metal2 18760 46200 18760 46200 0 _0081_
rlabel metal2 19152 44520 19152 44520 0 _0082_
rlabel metal2 18760 43064 18760 43064 0 _0083_
rlabel metal2 15848 25648 15848 25648 0 _0084_
rlabel metal2 12040 24808 12040 24808 0 _0085_
rlabel metal2 9128 25816 9128 25816 0 _0086_
rlabel metal2 8736 24024 8736 24024 0 _0087_
rlabel metal2 27944 30408 27944 30408 0 _0088_
rlabel metal3 24024 29624 24024 29624 0 _0089_
rlabel metal2 25480 26208 25480 26208 0 _0090_
rlabel metal2 26152 27888 26152 27888 0 _0091_
rlabel metal2 22568 32816 22568 32816 0 _0092_
rlabel metal2 23408 35000 23408 35000 0 _0093_
rlabel metal2 25704 33656 25704 33656 0 _0094_
rlabel metal2 26600 32144 26600 32144 0 _0095_
rlabel metal3 45472 3304 45472 3304 0 _0096_
rlabel metal2 49000 12656 49000 12656 0 _0097_
rlabel metal3 47656 15848 47656 15848 0 _0098_
rlabel metal2 43792 13608 43792 13608 0 _0099_
rlabel metal2 41944 12460 41944 12460 0 _0100_
rlabel metal2 30352 10024 30352 10024 0 _0101_
rlabel metal2 32648 11816 32648 11816 0 _0102_
rlabel metal2 31864 13272 31864 13272 0 _0103_
rlabel metal2 37240 14000 37240 14000 0 _0104_
rlabel metal2 34216 17080 34216 17080 0 _0105_
rlabel metal3 38976 16072 38976 16072 0 _0106_
rlabel metal3 40992 13944 40992 13944 0 _0107_
rlabel metal2 26768 3640 26768 3640 0 _0108_
rlabel metal2 25984 18648 25984 18648 0 _0109_
rlabel metal3 28336 18312 28336 18312 0 _0110_
rlabel metal2 38360 38360 38360 38360 0 _0111_
rlabel metal2 38920 39816 38920 39816 0 _0112_
rlabel metal2 37240 37520 37240 37520 0 _0113_
rlabel metal2 39144 41944 39144 41944 0 _0114_
rlabel metal2 37576 45976 37576 45976 0 _0115_
rlabel metal2 38864 45304 38864 45304 0 _0116_
rlabel metal2 37408 43512 37408 43512 0 _0117_
rlabel metal3 36848 41944 36848 41944 0 _0118_
rlabel metal3 30072 34328 30072 34328 0 _0119_
rlabel metal3 31136 36568 31136 36568 0 _0120_
rlabel metal2 26600 34608 26600 34608 0 _0121_
rlabel metal3 25480 35896 25480 35896 0 _0122_
rlabel metal3 34664 41272 34664 41272 0 _0123_
rlabel metal3 34216 38696 34216 38696 0 _0124_
rlabel metal2 26712 45360 26712 45360 0 _0125_
rlabel metal3 25760 42952 25760 42952 0 _0126_
rlabel metal2 34440 4816 34440 4816 0 _0127_
rlabel metal2 41496 10248 41496 10248 0 _0128_
rlabel metal2 43624 6692 43624 6692 0 _0129_
rlabel metal2 20944 18508 20944 18508 0 _0130_
rlabel metal2 33096 22680 33096 22680 0 _0131_
rlabel metal2 24024 22680 24024 22680 0 _0132_
rlabel metal2 25928 24864 25928 24864 0 _0133_
rlabel metal3 29232 23128 29232 23128 0 _0134_
rlabel metal2 34328 21112 34328 21112 0 _0135_
rlabel metal2 37240 22792 37240 22792 0 _0136_
rlabel metal2 38808 25872 38808 25872 0 _0137_
rlabel metal3 46536 20216 46536 20216 0 _0138_
rlabel metal2 47152 18648 47152 18648 0 _0139_
rlabel metal3 47600 23016 47600 23016 0 _0140_
rlabel metal2 48552 25816 48552 25816 0 _0141_
rlabel metal2 46032 25592 46032 25592 0 _0142_
rlabel metal2 49000 31976 49000 31976 0 _0143_
rlabel metal3 36064 38584 36064 38584 0 _0144_
rlabel metal2 36008 34552 36008 34552 0 _0145_
rlabel metal2 38808 35616 38808 35616 0 _0146_
rlabel metal3 42000 35896 42000 35896 0 _0147_
rlabel metal3 48272 34328 48272 34328 0 _0148_
rlabel metal2 47208 35280 47208 35280 0 _0149_
rlabel metal2 43736 36120 43736 36120 0 _0150_
rlabel metal2 49112 43288 49112 43288 0 _0151_
rlabel metal2 41664 38696 41664 38696 0 _0152_
rlabel metal3 45472 47544 45472 47544 0 _0153_
rlabel metal3 40992 44408 40992 44408 0 _0154_
rlabel metal2 40264 47124 40264 47124 0 _0155_
rlabel metal3 47600 46536 47600 46536 0 _0156_
rlabel metal2 44072 45024 44072 45024 0 _0157_
rlabel metal2 47208 42952 47208 42952 0 _0158_
rlabel metal2 48776 40712 48776 40712 0 _0159_
rlabel metal2 43288 21840 43288 21840 0 _0160_
rlabel metal3 26824 16912 26824 16912 0 _0161_
rlabel metal2 25704 16856 25704 16856 0 _0162_
rlabel metal3 26152 15064 26152 15064 0 _0163_
rlabel metal2 20888 17136 20888 17136 0 _0164_
rlabel metal2 20552 13776 20552 13776 0 _0165_
rlabel metal2 19096 16296 19096 16296 0 _0166_
rlabel metal3 16352 15176 16352 15176 0 _0167_
rlabel metal2 14280 13776 14280 13776 0 _0168_
rlabel metal2 14504 12600 14504 12600 0 _0169_
rlabel metal3 17304 12040 17304 12040 0 _0170_
rlabel metal3 16296 10472 16296 10472 0 _0171_
rlabel metal2 19432 9184 19432 9184 0 _0172_
rlabel metal2 14840 9352 14840 9352 0 _0173_
rlabel metal2 21336 9352 21336 9352 0 _0174_
rlabel metal3 23184 9912 23184 9912 0 _0175_
rlabel metal2 23464 11480 23464 11480 0 _0176_
rlabel metal2 24472 12600 24472 12600 0 _0177_
rlabel metal2 20104 19544 20104 19544 0 _0178_
rlabel metal2 19768 21560 19768 21560 0 _0179_
rlabel metal2 10472 19600 10472 19600 0 _0180_
rlabel metal3 11312 16296 11312 16296 0 _0181_
rlabel metal2 15288 16688 15288 16688 0 _0182_
rlabel metal2 14840 18032 14840 18032 0 _0183_
rlabel metal2 47040 29904 47040 29904 0 _0184_
rlabel metal2 13608 37744 13608 37744 0 _0185_
rlabel metal2 19320 38472 19320 38472 0 _0186_
rlabel metal3 9800 42168 9800 42168 0 _0187_
rlabel metal3 9688 44520 9688 44520 0 _0188_
rlabel metal2 11032 46928 11032 46928 0 _0189_
rlabel metal2 14840 47096 14840 47096 0 _0190_
rlabel metal2 15736 45416 15736 45416 0 _0191_
rlabel metal2 14840 43960 14840 43960 0 _0192_
rlabel metal2 7448 44184 7448 44184 0 _0193_
rlabel metal3 5992 41272 5992 41272 0 _0194_
rlabel metal2 5544 39704 5544 39704 0 _0195_
rlabel metal2 6440 37576 6440 37576 0 _0196_
rlabel metal2 22568 24976 22568 24976 0 _0197_
rlabel metal2 30520 33656 30520 33656 0 _0198_
rlabel metal2 29848 32088 29848 32088 0 _0199_
rlabel metal2 33880 32144 33880 32144 0 _0200_
rlabel metal2 33936 33432 33936 33432 0 _0201_
rlabel metal3 17640 31192 17640 31192 0 _0202_
rlabel metal2 19880 34300 19880 34300 0 _0203_
rlabel metal3 20104 25704 20104 25704 0 _0204_
rlabel metal2 17752 25816 17752 25816 0 _0205_
rlabel metal2 18424 28896 18424 28896 0 _0206_
rlabel metal2 16632 33712 16632 33712 0 _0207_
rlabel metal2 13832 33880 13832 33880 0 _0208_
rlabel metal2 11144 33432 11144 33432 0 _0209_
rlabel metal2 9576 29568 9576 29568 0 _0210_
rlabel metal2 13272 28224 13272 28224 0 _0211_
rlabel metal2 7784 29008 7784 29008 0 _0212_
rlabel metal2 7896 26964 7896 26964 0 _0213_
rlabel metal2 19320 23464 19320 23464 0 _0214_
rlabel metal2 26600 38416 26600 38416 0 _0215_
rlabel metal2 22680 38696 22680 38696 0 _0216_
rlabel metal2 25368 39816 25368 39816 0 _0217_
rlabel metal2 22680 40600 22680 40600 0 _0218_
rlabel metal2 21672 42056 21672 42056 0 _0219_
rlabel metal2 22624 45976 22624 45976 0 _0220_
rlabel metal3 21784 47544 21784 47544 0 _0221_
rlabel metal2 24808 46788 24808 46788 0 _0222_
rlabel metal2 29512 46256 29512 46256 0 _0223_
rlabel metal4 31192 46480 31192 46480 0 _0224_
rlabel metal2 36008 47096 36008 47096 0 _0225_
rlabel metal3 33264 47544 33264 47544 0 _0226_
rlabel metal2 29960 26824 29960 26824 0 _0227_
rlabel metal2 37912 19600 37912 19600 0 _0228_
rlabel metal2 38808 21112 38808 21112 0 _0229_
rlabel metal2 39760 17080 39760 17080 0 _0230_
rlabel metal2 42392 15400 42392 15400 0 _0231_
rlabel metal2 46872 16464 46872 16464 0 _0232_
rlabel metal2 48552 17976 48552 17976 0 _0233_
rlabel metal2 42840 17920 42840 17920 0 _0234_
rlabel metal2 40264 28224 40264 28224 0 _0235_
rlabel metal2 28392 26544 28392 26544 0 _0236_
rlabel metal2 29400 28112 29400 28112 0 _0237_
rlabel metal2 37240 24808 37240 24808 0 _0238_
rlabel metal3 36568 26824 36568 26824 0 _0239_
rlabel metal3 13944 6776 13944 6776 0 _0240_
rlabel metal2 36568 32032 36568 32032 0 _0241_
rlabel metal2 37352 34608 37352 34608 0 _0242_
rlabel metal2 40096 29624 40096 29624 0 _0243_
rlabel metal2 40712 32088 40712 32088 0 _0244_
rlabel metal2 43624 27104 43624 27104 0 _0245_
rlabel metal2 46872 28840 46872 28840 0 _0246_
rlabel metal3 46984 31192 46984 31192 0 _0247_
rlabel metal2 43624 31248 43624 31248 0 _0248_
rlabel metal3 36232 19320 36232 19320 0 _0249_
rlabel metal3 36456 18536 36456 18536 0 _0250_
rlabel metal2 25928 21112 25928 21112 0 _0251_
rlabel metal2 28392 21224 28392 21224 0 _0252_
rlabel metal2 41888 24696 41888 24696 0 _0253_
rlabel metal2 40040 26208 40040 26208 0 _0254_
rlabel metal2 39032 22680 39032 22680 0 _0255_
rlabel metal3 41384 27160 41384 27160 0 _0256_
rlabel metal2 34496 12852 34496 12852 0 _0257_
rlabel metal2 34888 12264 34888 12264 0 _0258_
rlabel metal2 33040 11368 33040 11368 0 _0259_
rlabel metal2 34216 14392 34216 14392 0 _0260_
rlabel metal3 36176 15064 36176 15064 0 _0261_
rlabel metal3 33208 13720 33208 13720 0 _0262_
rlabel metal2 35672 14540 35672 14540 0 _0263_
rlabel metal2 35840 14504 35840 14504 0 _0264_
rlabel metal2 36008 14420 36008 14420 0 _0265_
rlabel metal2 35616 15176 35616 15176 0 _0266_
rlabel metal2 39368 16800 39368 16800 0 _0267_
rlabel metal2 35672 16772 35672 16772 0 _0268_
rlabel metal2 39592 19040 39592 19040 0 _0269_
rlabel metal2 38808 15876 38808 15876 0 _0270_
rlabel metal2 39760 15288 39760 15288 0 _0271_
rlabel metal2 39144 15484 39144 15484 0 _0272_
rlabel metal2 39088 14420 39088 14420 0 _0273_
rlabel metal3 39340 14504 39340 14504 0 _0274_
rlabel metal2 39256 14308 39256 14308 0 _0275_
rlabel metal2 38864 16632 38864 16632 0 _0276_
rlabel metal2 27048 5824 27048 5824 0 _0277_
rlabel metal2 35252 28840 35252 28840 0 _0278_
rlabel metal3 29176 28616 29176 28616 0 _0279_
rlabel metal2 28840 20076 28840 20076 0 _0280_
rlabel metal2 28616 19670 28616 19670 0 _0281_
rlabel metal2 26376 18480 26376 18480 0 _0282_
rlabel metal2 28056 18592 28056 18592 0 _0283_
rlabel metal2 35168 30968 35168 30968 0 _0284_
rlabel metal2 38696 41664 38696 41664 0 _0285_
rlabel metal2 35728 39368 35728 39368 0 _0286_
rlabel metal2 40152 40936 40152 40936 0 _0287_
rlabel via2 36792 40390 36792 40390 0 _0288_
rlabel metal3 37828 38808 37828 38808 0 _0289_
rlabel metal2 39704 41216 39704 41216 0 _0290_
rlabel metal3 36652 38024 36652 38024 0 _0291_
rlabel metal2 38808 41664 38808 41664 0 _0292_
rlabel metal3 42308 26152 42308 26152 0 _0293_
rlabel metal2 38248 45164 38248 45164 0 _0294_
rlabel metal2 40488 41888 40488 41888 0 _0295_
rlabel metal2 37520 45472 37520 45472 0 _0296_
rlabel metal3 37828 45080 37828 45080 0 _0297_
rlabel metal2 37856 43064 37856 43064 0 _0298_
rlabel metal2 35616 42112 35616 42112 0 _0299_
rlabel metal2 28840 35672 28840 35672 0 _0300_
rlabel metal2 28840 35448 28840 35448 0 _0301_
rlabel metal2 29008 38808 29008 38808 0 _0302_
rlabel metal2 29624 36372 29624 36372 0 _0303_
rlabel metal2 29820 34104 29820 34104 0 _0304_
rlabel metal2 30156 35784 30156 35784 0 _0305_
rlabel metal2 26824 34944 26824 34944 0 _0306_
rlabel metal2 26152 35840 26152 35840 0 _0307_
rlabel metal2 29176 43470 29176 43470 0 _0308_
rlabel metal2 28952 43358 28952 43358 0 _0309_
rlabel metal2 33908 40488 33908 40488 0 _0310_
rlabel metal2 32480 38668 32480 38668 0 _0311_
rlabel metal2 28420 43624 28420 43624 0 _0312_
rlabel metal3 26628 42728 26628 42728 0 _0313_
rlabel metal2 43064 11200 43064 11200 0 _0314_
rlabel via1 42159 10584 42159 10584 0 _0315_
rlabel metal2 41776 9800 41776 9800 0 _0316_
rlabel metal3 21336 18424 21336 18424 0 _0317_
rlabel metal2 38528 21784 38528 21784 0 _0318_
rlabel metal2 33208 23912 33208 23912 0 _0319_
rlabel via1 26432 23159 26432 23159 0 _0320_
rlabel metal3 33376 24024 33376 24024 0 _0321_
rlabel metal3 27020 23576 27020 23576 0 _0322_
rlabel metal3 32340 23128 32340 23128 0 _0323_
rlabel metal3 25284 23128 25284 23128 0 _0324_
rlabel metal2 26880 24248 26880 24248 0 _0325_
rlabel metal2 29204 23128 29204 23128 0 _0326_
rlabel metal2 33992 21504 33992 21504 0 _0327_
rlabel metal2 36540 22344 36540 22344 0 _0328_
rlabel metal4 38696 25760 38696 25760 0 _0329_
rlabel metal2 47656 24920 47656 24920 0 _0330_
rlabel metal2 44912 25760 44912 25760 0 _0331_
rlabel metal3 45556 26264 45556 26264 0 _0332_
rlabel metal2 45864 25760 45864 25760 0 _0333_
rlabel metal2 45528 21638 45528 21638 0 _0334_
rlabel metal2 49168 21056 49168 21056 0 _0335_
rlabel metal2 46424 21467 46424 21467 0 _0336_
rlabel metal3 44884 23912 44884 23912 0 _0337_
rlabel metal3 47040 21560 47040 21560 0 _0338_
rlabel metal2 46424 20272 46424 20272 0 _0339_
rlabel metal2 46648 20104 46648 20104 0 _0340_
rlabel metal2 48608 20776 48608 20776 0 _0341_
rlabel metal2 47432 18984 47432 18984 0 _0342_
rlabel metal2 47656 22064 47656 22064 0 _0343_
rlabel metal3 48132 23912 48132 23912 0 _0344_
rlabel metal2 47768 23436 47768 23436 0 _0345_
rlabel metal2 48552 24696 48552 24696 0 _0346_
rlabel metal3 48160 24696 48160 24696 0 _0347_
rlabel metal2 49196 24808 49196 24808 0 _0348_
rlabel metal2 49168 19712 49168 19712 0 _0349_
rlabel metal2 45640 25284 45640 25284 0 _0350_
rlabel metal2 44240 40684 44240 40684 0 _0351_
rlabel metal2 46480 40880 46480 40880 0 _0352_
rlabel metal2 45192 41440 45192 41440 0 _0353_
rlabel metal3 45024 41272 45024 41272 0 _0354_
rlabel metal2 44772 45640 44772 45640 0 _0355_
rlabel metal2 45192 43596 45192 43596 0 _0356_
rlabel metal2 45752 43120 45752 43120 0 _0357_
rlabel metal2 46872 44464 46872 44464 0 _0358_
rlabel metal3 44408 44072 44408 44072 0 _0359_
rlabel metal2 42392 41020 42392 41020 0 _0360_
rlabel metal2 42000 40656 42000 40656 0 _0361_
rlabel metal2 45416 42764 45416 42764 0 _0362_
rlabel metal2 43736 42280 43736 42280 0 _0363_
rlabel metal2 42056 42392 42056 42392 0 _0364_
rlabel metal2 42616 42840 42616 42840 0 _0365_
rlabel metal2 43512 42056 43512 42056 0 _0366_
rlabel metal2 40992 43442 40992 43442 0 _0367_
rlabel metal3 40600 45080 40600 45080 0 _0368_
rlabel metal2 40488 42812 40488 42812 0 _0369_
rlabel metal2 43400 43008 43400 43008 0 _0370_
rlabel metal3 43932 42952 43932 42952 0 _0371_
rlabel metal2 45752 46424 45752 46424 0 _0372_
rlabel metal2 46088 45038 46088 45038 0 _0373_
rlabel metal3 45808 43848 45808 43848 0 _0374_
rlabel metal3 45080 43512 45080 43512 0 _0375_
rlabel metal2 45808 40460 45808 40460 0 _0376_
rlabel metal2 46984 39704 46984 39704 0 _0377_
rlabel metal2 45416 38724 45416 38724 0 _0378_
rlabel metal2 45248 31948 45248 31948 0 _0379_
rlabel metal2 45752 32620 45752 32620 0 _0380_
rlabel metal2 45640 33236 45640 33236 0 _0381_
rlabel metal2 42280 33712 42280 33712 0 _0382_
rlabel metal2 42280 32340 42280 32340 0 _0383_
rlabel metal2 40320 31472 40320 31472 0 _0384_
rlabel metal2 42000 33600 42000 33600 0 _0385_
rlabel metal2 38920 34468 38920 34468 0 _0386_
rlabel via2 40936 33300 40936 33300 0 _0387_
rlabel metal3 42168 32536 42168 32536 0 _0388_
rlabel via1 42784 33302 42784 33302 0 _0389_
rlabel metal2 42952 33236 42952 33236 0 _0390_
rlabel metal2 43026 32667 43026 32667 0 _0391_
rlabel metal3 44408 32424 44408 32424 0 _0392_
rlabel metal2 45304 32984 45304 32984 0 _0393_
rlabel metal2 47936 31304 47936 31304 0 _0394_
rlabel metal2 45192 32844 45192 32844 0 _0395_
rlabel metal2 44884 33208 44884 33208 0 _0396_
rlabel metal2 45602 38742 45602 38742 0 _0397_
rlabel metal2 45976 38920 45976 38920 0 _0398_
rlabel metal2 45640 41412 45640 41412 0 _0399_
rlabel metal2 44296 41888 44296 41888 0 _0400_
rlabel metal3 45752 39592 45752 39592 0 _0401_
rlabel metal2 42840 40236 42840 40236 0 _0402_
rlabel metal2 44912 40104 44912 40104 0 _0403_
rlabel metal2 43848 40376 43848 40376 0 _0404_
rlabel metal2 45640 39704 45640 39704 0 _0405_
rlabel metal3 46760 39704 46760 39704 0 _0406_
rlabel metal2 42392 21038 42392 21038 0 _0407_
rlabel metal3 41720 19880 41720 19880 0 _0408_
rlabel metal2 41412 18984 41412 18984 0 _0409_
rlabel metal2 24724 38696 24724 38696 0 _0410_
rlabel metal2 32984 34944 32984 34944 0 _0411_
rlabel metal2 44016 19992 44016 19992 0 _0412_
rlabel metal2 44072 18956 44072 18956 0 _0413_
rlabel metal2 43736 19908 43736 19908 0 _0414_
rlabel metal2 24164 39704 24164 39704 0 _0415_
rlabel metal3 35280 35672 35280 35672 0 _0416_
rlabel metal2 47262 39396 47262 39396 0 _0417_
rlabel via1 47264 38825 47264 38825 0 _0418_
rlabel metal2 42112 39200 42112 39200 0 _0419_
rlabel metal2 48720 38696 48720 38696 0 _0420_
rlabel metal2 49000 39088 49000 39088 0 _0421_
rlabel via1 47706 38822 47706 38822 0 _0422_
rlabel metal2 47936 38528 47936 38528 0 _0423_
rlabel metal2 45304 45584 45304 45584 0 _0424_
rlabel metal2 19300 20888 19300 20888 0 _0425_
rlabel metal2 34552 37352 34552 37352 0 _0426_
rlabel metal3 35448 38808 35448 38808 0 _0427_
rlabel metal3 40936 38024 40936 38024 0 _0428_
rlabel metal2 23800 36232 23800 36232 0 _0429_
rlabel metal2 20328 37968 20328 37968 0 _0430_
rlabel metal3 34692 33880 34692 33880 0 _0431_
rlabel metal2 41720 34944 41720 34944 0 _0432_
rlabel metal2 35672 35140 35672 35140 0 _0433_
rlabel metal3 49224 41720 49224 41720 0 _0434_
rlabel metal2 42056 34804 42056 34804 0 _0435_
rlabel metal2 41272 35573 41272 35573 0 _0436_
rlabel metal2 41104 34496 41104 34496 0 _0437_
rlabel metal2 39368 36344 39368 36344 0 _0438_
rlabel metal2 40264 36428 40264 36428 0 _0439_
rlabel metal2 43288 34944 43288 34944 0 _0440_
rlabel metal2 43624 35168 43624 35168 0 _0441_
rlabel metal2 41720 36540 41720 36540 0 _0442_
rlabel metal3 47824 35672 47824 35672 0 _0443_
rlabel metal3 46452 36344 46452 36344 0 _0444_
rlabel metal2 48776 35728 48776 35728 0 _0445_
rlabel metal2 47096 36092 47096 36092 0 _0446_
rlabel metal2 47320 34720 47320 34720 0 _0447_
rlabel metal2 44884 35112 44884 35112 0 _0448_
rlabel metal3 45584 36456 45584 36456 0 _0449_
rlabel via2 43848 36448 43848 36448 0 _0450_
rlabel metal2 45276 37912 45276 37912 0 _0451_
rlabel metal3 44016 38136 44016 38136 0 _0452_
rlabel metal2 44632 39172 44632 39172 0 _0453_
rlabel via2 41608 38016 41608 38016 0 _0454_
rlabel metal2 46592 46088 46592 46088 0 _0455_
rlabel metal2 41832 45920 41832 45920 0 _0456_
rlabel metal2 42840 44352 42840 44352 0 _0457_
rlabel metal2 43848 46200 43848 46200 0 _0458_
rlabel metal2 42560 44576 42560 44576 0 _0459_
rlabel metal2 41692 44240 41692 44240 0 _0460_
rlabel metal2 40824 46144 40824 46144 0 _0461_
rlabel metal2 45976 44520 45976 44520 0 _0462_
rlabel metal2 40264 46487 40264 46487 0 _0463_
rlabel metal2 45668 44520 45668 44520 0 _0464_
rlabel metal2 46424 44464 46424 44464 0 _0465_
rlabel metal2 46088 46172 46088 46172 0 _0466_
rlabel metal2 47768 44763 47768 44763 0 _0467_
rlabel metal3 47712 45080 47712 45080 0 _0468_
rlabel metal3 45976 44296 45976 44296 0 _0469_
rlabel metal2 48104 40600 48104 40600 0 _0470_
rlabel metal2 48776 39816 48776 39816 0 _0471_
rlabel metal2 44072 23016 44072 23016 0 _0472_
rlabel metal2 44856 23856 44856 23856 0 _0473_
rlabel metal3 44072 24696 44072 24696 0 _0474_
rlabel metal2 45134 24192 45134 24192 0 _0475_
rlabel via1 45732 22328 45732 22328 0 _0476_
rlabel metal2 45976 22904 45976 22904 0 _0477_
rlabel metal2 43624 22232 43624 22232 0 _0478_
rlabel metal2 26600 16184 26600 16184 0 _0479_
rlabel metal2 23128 17808 23128 17808 0 _0480_
rlabel metal2 23240 16744 23240 16744 0 _0481_
rlabel metal2 23128 10430 23128 10430 0 _0482_
rlabel metal2 21448 17388 21448 17388 0 _0483_
rlabel metal2 24640 17360 24640 17360 0 _0484_
rlabel metal2 23128 16968 23128 16968 0 _0485_
rlabel metal2 24136 16996 24136 16996 0 _0486_
rlabel metal3 27468 16856 27468 16856 0 _0487_
rlabel metal3 24920 17640 24920 17640 0 _0488_
rlabel metal2 25872 17696 25872 17696 0 _0489_
rlabel metal2 23016 15792 23016 15792 0 _0490_
rlabel metal2 23352 16156 23352 16156 0 _0491_
rlabel metal3 24696 21000 24696 21000 0 _0492_
rlabel metal3 25200 23912 25200 23912 0 _0493_
rlabel metal2 24528 16072 24528 16072 0 _0494_
rlabel metal2 25144 15624 25144 15624 0 _0495_
rlabel metal2 20720 16352 20720 16352 0 _0496_
rlabel metal2 19130 17155 19130 17155 0 _0497_
rlabel metal2 22176 17332 22176 17332 0 _0498_
rlabel metal2 19544 15736 19544 15736 0 _0499_
rlabel metal3 24304 15624 24304 15624 0 _0500_
rlabel metal2 20664 13832 20664 13832 0 _0501_
rlabel metal2 19712 14560 19712 14560 0 _0502_
rlabel metal2 18200 16744 18200 16744 0 _0503_
rlabel metal2 17752 15848 17752 15848 0 _0504_
rlabel metal2 18872 15792 18872 15792 0 _0505_
rlabel metal2 16800 13580 16800 13580 0 _0506_
rlabel metal2 18256 15596 18256 15596 0 _0507_
rlabel metal2 17864 13216 17864 13216 0 _0508_
rlabel metal3 19741 11368 19741 11368 0 _0509_
rlabel metal2 18256 13244 18256 13244 0 _0510_
rlabel metal2 17640 11256 17640 11256 0 _0511_
rlabel metal3 19320 12936 19320 12936 0 _0512_
rlabel metal2 18256 12236 18256 12236 0 _0513_
rlabel metal2 19320 10920 19320 10920 0 _0514_
rlabel metal2 19768 11648 19768 11648 0 _0515_
rlabel metal2 19600 12096 19600 12096 0 _0516_
rlabel metal2 18760 9856 18760 9856 0 _0517_
rlabel metal2 17584 10668 17584 10668 0 _0518_
rlabel metal2 19208 9800 19208 9800 0 _0519_
rlabel metal2 19030 10721 19030 10721 0 _0520_
rlabel metal2 19600 9268 19600 9268 0 _0521_
rlabel metal3 20720 9800 20720 9800 0 _0522_
rlabel metal2 21560 10640 21560 10640 0 _0523_
rlabel metal2 19712 10108 19712 10108 0 _0524_
rlabel metal2 21448 10528 21448 10528 0 _0525_
rlabel metal2 20832 9856 20832 9856 0 _0526_
rlabel metal2 24472 10808 24472 10808 0 _0527_
rlabel metal2 22512 10528 22512 10528 0 _0528_
rlabel metal2 25256 13552 25256 13552 0 _0529_
rlabel metal2 23800 11088 23800 11088 0 _0530_
rlabel metal2 17864 10500 17864 10500 0 _0531_
rlabel metal2 18144 11704 18144 11704 0 _0532_
rlabel metal3 23688 11368 23688 11368 0 _0533_
rlabel metal2 21700 11592 21700 11592 0 _0534_
rlabel metal2 21952 12320 21952 12320 0 _0535_
rlabel metal2 17416 14420 17416 14420 0 _0536_
rlabel metal2 23240 14084 23240 14084 0 _0537_
rlabel metal2 23800 14616 23800 14616 0 _0538_
rlabel metal2 24024 12908 24024 12908 0 _0539_
rlabel metal3 25536 16072 25536 16072 0 _0540_
rlabel metal2 24640 12068 24640 12068 0 _0541_
rlabel metal3 18592 19992 18592 19992 0 _0542_
rlabel metal2 17528 23044 17528 23044 0 _0543_
rlabel metal2 17472 21112 17472 21112 0 _0544_
rlabel metal2 12320 20076 12320 20076 0 _0545_
rlabel metal2 12600 20132 12600 20132 0 _0546_
rlabel metal2 14222 19488 14222 19488 0 _0547_
rlabel metal2 16464 19292 16464 19292 0 _0548_
rlabel metal2 15624 19068 15624 19068 0 _0549_
rlabel metal2 13776 18760 13776 18760 0 _0550_
rlabel metal2 16744 19432 16744 19432 0 _0551_
rlabel metal2 17528 18480 17528 18480 0 _0552_
rlabel metal3 15708 19208 15708 19208 0 _0553_
rlabel metal2 17024 19488 17024 19488 0 _0554_
rlabel metal2 17808 18816 17808 18816 0 _0555_
rlabel metal2 18760 19712 18760 19712 0 _0556_
rlabel metal2 18648 19852 18648 19852 0 _0557_
rlabel metal2 19264 18760 19264 18760 0 _0558_
rlabel metal2 19544 21112 19544 21112 0 _0559_
rlabel metal2 19180 22344 19180 22344 0 _0560_
rlabel metal2 16184 17528 16184 17528 0 _0561_
rlabel metal2 16184 18648 16184 18648 0 _0562_
rlabel metal2 11648 18536 11648 18536 0 _0563_
rlabel metal3 12684 17640 12684 17640 0 _0564_
rlabel metal2 12264 17682 12264 17682 0 _0565_
rlabel metal2 15176 16632 15176 16632 0 _0566_
rlabel metal2 12040 16772 12040 16772 0 _0567_
rlabel metal2 16408 16934 16408 16934 0 _0568_
rlabel metal2 15960 17506 15960 17506 0 _0569_
rlabel metal2 9576 41160 9576 41160 0 _0570_
rlabel metal3 10416 41160 10416 41160 0 _0571_
rlabel metal2 10696 40432 10696 40432 0 _0572_
rlabel metal3 10472 40264 10472 40264 0 _0573_
rlabel metal2 21224 46144 21224 46144 0 _0574_
rlabel metal3 17164 44632 17164 44632 0 _0575_
rlabel metal2 17304 37884 17304 37884 0 _0576_
rlabel metal2 16772 37464 16772 37464 0 _0577_
rlabel metal2 15512 39312 15512 39312 0 _0578_
rlabel metal2 15624 39760 15624 39760 0 _0579_
rlabel metal2 12824 40376 12824 40376 0 _0580_
rlabel metal2 13272 40572 13272 40572 0 _0581_
rlabel metal2 14840 39900 14840 39900 0 _0582_
rlabel metal2 16632 39648 16632 39648 0 _0583_
rlabel metal2 12600 42252 12600 42252 0 _0584_
rlabel metal2 12992 42728 12992 42728 0 _0585_
rlabel metal2 14168 42588 14168 42588 0 _0586_
rlabel metal2 14590 40916 14590 40916 0 _0587_
rlabel metal2 16744 39648 16744 39648 0 _0588_
rlabel metal2 15904 38892 15904 38892 0 _0589_
rlabel metal2 16968 40488 16968 40488 0 _0590_
rlabel via2 18088 44282 18088 44282 0 _0591_
rlabel metal2 17360 43932 17360 43932 0 _0592_
rlabel metal2 18816 41636 18816 41636 0 _0593_
rlabel metal3 17836 46424 17836 46424 0 _0594_
rlabel metal2 18424 43204 18424 43204 0 _0595_
rlabel metal2 17528 42252 17528 42252 0 _0596_
rlabel metal2 19096 41384 19096 41384 0 _0597_
rlabel metal2 16688 44072 16688 44072 0 _0598_
rlabel metal2 15960 41678 15960 41678 0 _0599_
rlabel metal3 17556 41944 17556 41944 0 _0600_
rlabel metal2 19376 39816 19376 39816 0 _0601_
rlabel metal2 11480 40516 11480 40516 0 _0602_
rlabel metal2 9016 38976 9016 38976 0 _0603_
rlabel metal3 9968 38024 9968 38024 0 _0604_
rlabel metal2 9240 38388 9240 38388 0 _0605_
rlabel metal3 10276 38248 10276 38248 0 _0606_
rlabel metal3 12320 38808 12320 38808 0 _0607_
rlabel metal2 11086 39340 11086 39340 0 _0608_
rlabel metal2 12040 39630 12040 39630 0 _0609_
rlabel metal2 10472 38976 10472 38976 0 _0610_
rlabel metal2 12488 38864 12488 38864 0 _0611_
rlabel metal2 15848 40712 15848 40712 0 _0612_
rlabel metal2 16520 40096 16520 40096 0 _0613_
rlabel metal2 10248 41020 10248 41020 0 _0614_
rlabel metal2 15848 37912 15848 37912 0 _0615_
rlabel metal2 14672 38892 14672 38892 0 _0616_
rlabel metal2 15736 39144 15736 39144 0 _0617_
rlabel metal3 12880 40264 12880 40264 0 _0618_
rlabel metal2 14056 40376 14056 40376 0 _0619_
rlabel metal2 13160 39536 13160 39536 0 _0620_
rlabel metal2 12432 39508 12432 39508 0 _0621_
rlabel metal2 16184 41432 16184 41432 0 _0622_
rlabel metal2 16072 40936 16072 40936 0 _0623_
rlabel metal2 12992 28056 12992 28056 0 _0624_
rlabel metal2 17640 24276 17640 24276 0 _0625_
rlabel metal2 12096 38024 12096 38024 0 _0626_
rlabel metal3 12040 38024 12040 38024 0 _0627_
rlabel metal2 12600 37688 12600 37688 0 _0628_
rlabel metal2 13272 37576 13272 37576 0 _0629_
rlabel metal2 16184 44184 16184 44184 0 _0630_
rlabel metal2 10808 43030 10808 43030 0 _0631_
rlabel metal2 20216 37576 20216 37576 0 _0632_
rlabel metal2 18648 37722 18648 37722 0 _0633_
rlabel metal2 11256 40544 11256 40544 0 _0634_
rlabel metal2 10920 43456 10920 43456 0 _0635_
rlabel metal2 11816 42616 11816 42616 0 _0636_
rlabel metal2 10360 42056 10360 42056 0 _0637_
rlabel metal2 13496 45864 13496 45864 0 _0638_
rlabel metal2 12488 43960 12488 43960 0 _0639_
rlabel metal2 9464 44240 9464 44240 0 _0640_
rlabel metal3 13076 46424 13076 46424 0 _0641_
rlabel metal3 11760 45864 11760 45864 0 _0642_
rlabel metal2 11816 47152 11816 47152 0 _0643_
rlabel metal2 14952 47592 14952 47592 0 _0644_
rlabel metal2 13888 44968 13888 44968 0 _0645_
rlabel metal2 15624 45158 15624 45158 0 _0646_
rlabel via1 14382 42728 14382 42728 0 _0647_
rlabel metal2 15960 44106 15960 44106 0 _0648_
rlabel metal2 7467 42896 7467 42896 0 _0649_
rlabel metal2 7224 43120 7224 43120 0 _0650_
rlabel metal3 7364 41944 7364 41944 0 _0651_
rlabel metal2 6888 39628 6888 39628 0 _0652_
rlabel metal2 6664 39872 6664 39872 0 _0653_
rlabel metal2 5880 41104 5880 41104 0 _0654_
rlabel metal3 6160 38920 6160 38920 0 _0655_
rlabel metal2 6272 37324 6272 37324 0 _0656_
rlabel metal3 23352 23912 23352 23912 0 _0657_
rlabel metal2 23940 24136 23940 24136 0 _0658_
rlabel metal2 32172 30408 32172 30408 0 _0659_
rlabel metal2 33880 32676 33880 32676 0 _0660_
rlabel via2 33656 32550 33656 32550 0 _0661_
rlabel metal2 33152 32704 33152 32704 0 _0662_
rlabel metal2 38808 31136 38808 31136 0 _0663_
rlabel metal2 31612 31080 31612 31080 0 _0664_
rlabel via2 40936 30985 40936 30985 0 _0665_
rlabel metal2 34496 31304 34496 31304 0 _0666_
rlabel metal3 39088 26488 39088 26488 0 _0667_
rlabel metal2 35140 32648 35140 32648 0 _0668_
rlabel metal3 11368 27048 11368 27048 0 _0669_
rlabel metal2 10696 27104 10696 27104 0 _0670_
rlabel metal3 14952 27384 14952 27384 0 _0671_
rlabel metal3 12964 27048 12964 27048 0 _0672_
rlabel metal2 14784 27832 14784 27832 0 _0673_
rlabel metal2 11424 30184 11424 30184 0 _0674_
rlabel metal2 14112 30044 14112 30044 0 _0675_
rlabel via2 13384 30985 13384 30985 0 _0676_
rlabel metal2 12740 31024 12740 31024 0 _0677_
rlabel metal2 15064 30506 15064 30506 0 _0678_
rlabel metal2 13944 31668 13944 31668 0 _0679_
rlabel metal2 14056 31444 14056 31444 0 _0680_
rlabel metal2 14728 33208 14728 33208 0 _0681_
rlabel metal3 14672 32648 14672 32648 0 _0682_
rlabel metal2 19992 33236 19992 33236 0 _0683_
rlabel metal2 20636 32312 20636 32312 0 _0684_
rlabel metal2 22512 31668 22512 31668 0 _0685_
rlabel metal2 23016 30912 23016 30912 0 _0686_
rlabel metal2 22568 30744 22568 30744 0 _0687_
rlabel metal2 20440 31052 20440 31052 0 _0688_
rlabel metal3 21812 30968 21812 30968 0 _0689_
rlabel via2 22456 27850 22456 27850 0 _0690_
rlabel metal2 23016 27552 23016 27552 0 _0691_
rlabel metal2 21336 29176 21336 29176 0 _0692_
rlabel via1 21728 30152 21728 30152 0 _0693_
rlabel metal2 21700 25704 21700 25704 0 _0694_
rlabel metal2 21224 27552 21224 27552 0 _0695_
rlabel metal2 21896 28826 21896 28826 0 _0696_
rlabel metal2 22176 28448 22176 28448 0 _0697_
rlabel via1 21952 30152 21952 30152 0 _0698_
rlabel metal2 22092 30408 22092 30408 0 _0699_
rlabel via2 19768 33306 19768 33306 0 _0700_
rlabel metal2 20468 33208 20468 33208 0 _0701_
rlabel metal2 14504 31794 14504 31794 0 _0702_
rlabel via1 14784 30166 14784 30166 0 _0703_
rlabel metal2 14952 28112 14952 28112 0 _0704_
rlabel metal3 12796 26936 12796 26936 0 _0705_
rlabel metal2 15098 27907 15098 27907 0 _0706_
rlabel metal2 15736 27328 15736 27328 0 _0707_
rlabel metal2 16296 28664 16296 28664 0 _0708_
rlabel metal2 16184 27664 16184 27664 0 _0709_
rlabel metal2 18648 30072 18648 30072 0 _0710_
rlabel metal3 16576 27832 16576 27832 0 _0711_
rlabel metal2 15176 27216 15176 27216 0 _0712_
rlabel metal2 14896 27440 14896 27440 0 _0713_
rlabel metal3 13832 31080 13832 31080 0 _0714_
rlabel metal2 21952 29400 21952 29400 0 _0715_
rlabel metal2 22568 29484 22568 29484 0 _0716_
rlabel metal2 17416 31136 17416 31136 0 _0717_
rlabel metal2 15680 29680 15680 29680 0 _0718_
rlabel metal2 16014 30464 16014 30464 0 _0719_
rlabel metal2 21112 29478 21112 29478 0 _0720_
rlabel metal3 22064 29288 22064 29288 0 _0721_
rlabel metal2 15288 28896 15288 28896 0 _0722_
rlabel metal3 14672 28616 14672 28616 0 _0723_
rlabel metal2 15932 27048 15932 27048 0 _0724_
rlabel metal2 17304 24416 17304 24416 0 _0725_
rlabel metal2 17304 26572 17304 26572 0 _0726_
rlabel metal2 12824 29624 12824 29624 0 _0727_
rlabel metal2 19096 30268 19096 30268 0 _0728_
rlabel metal2 19376 30296 19376 30296 0 _0729_
rlabel metal2 12488 33264 12488 33264 0 _0730_
rlabel metal2 21000 34552 21000 34552 0 _0731_
rlabel metal3 20580 35672 20580 35672 0 _0732_
rlabel metal2 20104 34238 20104 34238 0 _0733_
rlabel metal2 10024 29064 10024 29064 0 _0734_
rlabel metal2 18984 27202 18984 27202 0 _0735_
rlabel metal2 19740 27048 19740 27048 0 _0736_
rlabel metal2 19600 26152 19600 26152 0 _0737_
rlabel metal2 17864 27972 17864 27972 0 _0738_
rlabel metal3 18424 27832 18424 27832 0 _0739_
rlabel metal2 17808 27496 17808 27496 0 _0740_
rlabel metal3 17369 34104 17369 34104 0 _0741_
rlabel metal3 17920 30184 17920 30184 0 _0742_
rlabel metal2 17752 29316 17752 29316 0 _0743_
rlabel metal3 17136 34216 17136 34216 0 _0744_
rlabel metal2 13272 32431 13272 32431 0 _0745_
rlabel via2 12824 33312 12824 33312 0 _0746_
rlabel metal3 12049 31752 12049 31752 0 _0747_
rlabel metal2 11032 32368 11032 32368 0 _0748_
rlabel metal2 11704 30800 11704 30800 0 _0749_
rlabel metal2 9688 29478 9688 29478 0 _0750_
rlabel metal2 11704 28840 11704 28840 0 _0751_
rlabel metal2 8139 28028 8139 28028 0 _0752_
rlabel metal2 12152 29064 12152 29064 0 _0753_
rlabel metal2 12712 29372 12712 29372 0 _0754_
rlabel metal2 7896 28448 7896 28448 0 _0755_
rlabel metal2 9688 27328 9688 27328 0 _0756_
rlabel metal2 18368 23212 18368 23212 0 _0757_
rlabel metal2 18200 23968 18200 23968 0 _0758_
rlabel metal3 17668 24136 17668 24136 0 _0759_
rlabel metal2 18984 23408 18984 23408 0 _0760_
rlabel metal2 24976 42588 24976 42588 0 _0761_
rlabel metal2 27944 41426 27944 41426 0 _0762_
rlabel via1 30072 41958 30072 41958 0 _0763_
rlabel metal2 24584 41048 24584 41048 0 _0764_
rlabel metal2 29008 40544 29008 40544 0 _0765_
rlabel metal3 29120 40488 29120 40488 0 _0766_
rlabel metal2 31080 40712 31080 40712 0 _0767_
rlabel metal2 29400 37940 29400 37940 0 _0768_
rlabel metal2 30632 37744 30632 37744 0 _0769_
rlabel metal2 30464 39592 30464 39592 0 _0770_
rlabel metal2 30912 39592 30912 39592 0 _0771_
rlabel metal3 30352 39592 30352 39592 0 _0772_
rlabel metal2 26656 40460 26656 40460 0 _0773_
rlabel metal2 27720 39760 27720 39760 0 _0774_
rlabel metal3 29176 39592 29176 39592 0 _0775_
rlabel via1 29792 41961 29792 41961 0 _0776_
rlabel metal2 29568 42224 29568 42224 0 _0777_
rlabel metal2 30184 43232 30184 43232 0 _0778_
rlabel metal2 24584 46928 24584 46928 0 _0779_
rlabel metal3 30044 44296 30044 44296 0 _0780_
rlabel metal2 27720 44156 27720 44156 0 _0781_
rlabel metal3 29624 43512 29624 43512 0 _0782_
rlabel metal2 33264 43428 33264 43428 0 _0783_
rlabel metal2 32648 45360 32648 45360 0 _0784_
rlabel metal3 32480 43624 32480 43624 0 _0785_
rlabel metal2 31136 43512 31136 43512 0 _0786_
rlabel metal2 31416 43764 31416 43764 0 _0787_
rlabel metal2 32256 43960 32256 43960 0 _0788_
rlabel metal2 32816 42812 32816 42812 0 _0789_
rlabel metal2 32648 42112 32648 42112 0 _0790_
rlabel metal2 35000 43414 35000 43414 0 _0791_
rlabel metal2 35672 42784 35672 42784 0 _0792_
rlabel metal2 34804 42168 34804 42168 0 _0793_
rlabel metal2 35448 42776 35448 42776 0 _0794_
rlabel metal2 32536 42616 32536 42616 0 _0795_
rlabel metal2 36120 43064 36120 43064 0 _0796_
rlabel metal3 33544 42728 33544 42728 0 _0797_
rlabel metal2 32872 40432 32872 40432 0 _0798_
rlabel metal2 26040 37800 26040 37800 0 _0799_
rlabel metal2 31808 38360 31808 38360 0 _0800_
rlabel metal2 31248 39060 31248 39060 0 _0801_
rlabel metal2 31472 38696 31472 38696 0 _0802_
rlabel metal2 31360 40264 31360 40264 0 _0803_
rlabel metal2 30296 40572 30296 40572 0 _0804_
rlabel metal2 30632 44044 30632 44044 0 _0805_
rlabel metal3 33936 43512 33936 43512 0 _0806_
rlabel metal2 30968 42700 30968 42700 0 _0807_
rlabel metal2 31192 42840 31192 42840 0 _0808_
rlabel metal2 31304 41860 31304 41860 0 _0809_
rlabel metal2 31416 41356 31416 41356 0 _0810_
rlabel metal2 32760 40320 32760 40320 0 _0811_
rlabel metal2 22680 36568 22680 36568 0 _0812_
rlabel metal3 25480 38808 25480 38808 0 _0813_
rlabel metal2 23576 41216 23576 41216 0 _0814_
rlabel metal2 26712 38192 26712 38192 0 _0815_
rlabel metal2 27132 38808 27132 38808 0 _0816_
rlabel metal2 23296 45864 23296 45864 0 _0817_
rlabel metal2 24640 39592 24640 39592 0 _0818_
rlabel metal2 23436 36680 23436 36680 0 _0819_
rlabel metal2 22988 38864 22988 38864 0 _0820_
rlabel metal2 26152 40488 26152 40488 0 _0821_
rlabel metal3 24752 38696 24752 38696 0 _0822_
rlabel metal2 24976 40096 24976 40096 0 _0823_
rlabel metal2 25816 40068 25816 40068 0 _0824_
rlabel metal2 24444 43568 24444 43568 0 _0825_
rlabel metal2 22456 38780 22456 38780 0 _0826_
rlabel metal2 23464 40964 23464 40964 0 _0827_
rlabel metal2 21896 43596 21896 43596 0 _0828_
rlabel metal3 23184 43512 23184 43512 0 _0829_
rlabel metal2 22008 42812 22008 42812 0 _0830_
rlabel metal3 22792 45024 22792 45024 0 _0831_
rlabel metal3 24304 44408 24304 44408 0 _0832_
rlabel metal2 23464 47208 23464 47208 0 _0833_
rlabel via1 25611 46663 25611 46663 0 _0834_
rlabel metal2 25368 46928 25368 46928 0 _0835_
rlabel metal2 30576 46648 30576 46648 0 _0836_
rlabel via1 29456 45849 29456 45849 0 _0837_
rlabel metal2 31500 46677 31500 46677 0 _0838_
rlabel metal3 31668 45080 31668 45080 0 _0839_
rlabel metal2 31304 45248 31304 45248 0 _0840_
rlabel metal2 30856 47208 30856 47208 0 _0841_
rlabel metal2 34776 44520 34776 44520 0 _0842_
rlabel metal2 35784 45416 35784 45416 0 _0843_
rlabel metal3 29736 23912 29736 23912 0 _0844_
rlabel metal2 28560 24304 28560 24304 0 _0845_
rlabel metal2 40292 19208 40292 19208 0 _0846_
rlabel metal2 39704 21336 39704 21336 0 _0847_
rlabel metal2 41776 17612 41776 17612 0 _0848_
rlabel metal2 42336 16856 42336 16856 0 _0849_
rlabel metal2 40488 17024 40488 17024 0 _0850_
rlabel metal3 42196 16632 42196 16632 0 _0851_
rlabel metal2 42840 15960 42840 15960 0 _0852_
rlabel via2 42280 15295 42280 15295 0 _0853_
rlabel metal3 46200 16856 46200 16856 0 _0854_
rlabel metal3 45192 15176 45192 15176 0 _0855_
rlabel metal2 46928 15960 46928 15960 0 _0856_
rlabel metal2 45686 18424 45686 18424 0 _0857_
rlabel metal2 46088 16716 46088 16716 0 _0858_
rlabel metal2 46340 16968 46340 16968 0 _0859_
rlabel metal3 47012 18424 47012 18424 0 _0860_
rlabel metal2 42616 18312 42616 18312 0 _0861_
rlabel metal2 43176 17920 43176 17920 0 _0862_
rlabel metal2 38472 28532 38472 28532 0 _0863_
rlabel metal3 37716 27608 37716 27608 0 _0864_
rlabel metal2 38388 27272 38388 27272 0 _0865_
rlabel metal2 39178 27907 39178 27907 0 _0866_
rlabel metal2 39144 27328 39144 27328 0 _0867_
rlabel metal2 39424 27328 39424 27328 0 _0868_
rlabel metal3 32256 27048 32256 27048 0 _0869_
rlabel metal2 28616 27104 28616 27104 0 _0870_
rlabel metal2 28056 25984 28056 25984 0 _0871_
rlabel via2 31752 26283 31752 26283 0 _0872_
rlabel metal2 28336 27048 28336 27048 0 _0873_
rlabel metal3 28588 27048 28588 27048 0 _0874_
rlabel metal2 31444 27048 31444 27048 0 _0875_
rlabel metal2 31640 26124 31640 26124 0 _0876_
rlabel metal3 31696 26376 31696 26376 0 _0877_
rlabel metal3 30268 27272 30268 27272 0 _0878_
rlabel metal2 35112 25760 35112 25760 0 _0879_
rlabel metal2 34300 24920 34300 24920 0 _0880_
rlabel metal3 35056 25480 35056 25480 0 _0881_
rlabel metal3 35756 25480 35756 25480 0 _0882_
rlabel metal3 34636 27048 34636 27048 0 _0883_
rlabel metal2 33852 25256 33852 25256 0 _0884_
rlabel metal2 34664 26432 34664 26432 0 _0885_
rlabel metal2 35420 27048 35420 27048 0 _0886_
rlabel metal2 12600 7728 12600 7728 0 _0887_
rlabel metal2 39032 29232 39032 29232 0 _0888_
rlabel metal2 39032 30926 39032 30926 0 _0889_
rlabel metal2 42560 30968 42560 30968 0 _0890_
rlabel via1 39256 30982 39256 30982 0 _0891_
rlabel metal2 39704 32760 39704 32760 0 _0892_
rlabel metal2 39760 31360 39760 31360 0 _0893_
rlabel metal2 40488 29680 40488 29680 0 _0894_
rlabel metal3 40572 32536 40572 32536 0 _0895_
rlabel metal2 42672 29960 42672 29960 0 _0896_
rlabel via2 43624 30170 43624 30170 0 _0897_
rlabel metal2 43372 28504 43372 28504 0 _0898_
rlabel metal2 45388 29400 45388 29400 0 _0899_
rlabel metal2 45696 30688 45696 30688 0 _0900_
rlabel metal2 43988 30408 43988 30408 0 _0901_
rlabel metal2 34888 20880 34888 20880 0 _0902_
rlabel metal2 33880 19894 33880 19894 0 _0903_
rlabel metal2 34384 20160 34384 20160 0 _0904_
rlabel metal2 33936 18536 33936 18536 0 _0905_
rlabel metal2 28168 23318 28168 23318 0 _0906_
rlabel metal2 28168 22036 28168 22036 0 _0907_
rlabel metal2 26600 21896 26600 21896 0 _0908_
rlabel metal3 28980 20776 28980 20776 0 _0909_
rlabel via1 39872 24735 39872 24735 0 _0910_
rlabel metal2 40320 25032 40320 25032 0 _0911_
rlabel metal3 39284 25704 39284 25704 0 _0912_
rlabel metal2 39032 23464 39032 23464 0 _0913_
rlabel metal2 40208 26628 40208 26628 0 _0914_
rlabel metal2 22960 6188 22960 6188 0 _0915_
rlabel metal2 14392 4424 14392 4424 0 _0916_
rlabel metal2 15736 4368 15736 4368 0 _0917_
rlabel metal3 20655 5880 20655 5880 0 _0918_
rlabel metal2 26170 4480 26170 4480 0 _0919_
rlabel metal2 43176 20832 43176 20832 0 _0920_
rlabel metal2 30184 16660 30184 16660 0 _0921_
rlabel via2 31976 18437 31976 18437 0 _0922_
rlabel metal3 33684 17864 33684 17864 0 _0923_
rlabel metal2 31752 18732 31752 18732 0 _0924_
rlabel metal2 31528 8743 31528 8743 0 _0925_
rlabel metal2 30968 21672 30968 21672 0 _0926_
rlabel metal2 31304 21644 31304 21644 0 _0927_
rlabel metal2 24808 17584 24808 17584 0 _0928_
rlabel metal3 32312 21560 32312 21560 0 _0929_
rlabel metal3 31864 21448 31864 21448 0 _0930_
rlabel metal2 31752 14552 31752 14552 0 _0931_
rlabel metal3 33572 19992 33572 19992 0 _0932_
rlabel metal2 31528 21476 31528 21476 0 _0933_
rlabel metal2 31080 19684 31080 19684 0 _0934_
rlabel metal2 30800 19908 30800 19908 0 _0935_
rlabel via2 31864 11360 31864 11360 0 _0936_
rlabel metal2 33300 8316 33300 8316 0 _0937_
rlabel metal3 37912 8232 37912 8232 0 _0938_
rlabel metal2 33880 8316 33880 8316 0 _0939_
rlabel metal2 5320 30520 5320 30520 0 _0940_
rlabel metal3 11088 12152 11088 12152 0 _0941_
rlabel metal3 7560 12208 7560 12208 0 _0942_
rlabel metal2 7560 13328 7560 13328 0 _0943_
rlabel metal2 7756 21000 7756 21000 0 _0944_
rlabel metal2 6272 18788 6272 18788 0 _0945_
rlabel metal2 6048 20300 6048 20300 0 _0946_
rlabel metal2 7336 20104 7336 20104 0 _0947_
rlabel metal2 6720 16324 6720 16324 0 _0948_
rlabel metal3 6664 15176 6664 15176 0 _0949_
rlabel metal2 7112 17416 7112 17416 0 _0950_
rlabel metal2 7168 14504 7168 14504 0 _0951_
rlabel metal2 7224 13272 7224 13272 0 _0952_
rlabel metal2 7336 12236 7336 12236 0 _0953_
rlabel metal2 7336 10175 7336 10175 0 _0954_
rlabel metal2 9744 5488 9744 5488 0 _0955_
rlabel metal2 7784 8988 7784 8988 0 _0956_
rlabel metal2 6328 10080 6328 10080 0 _0957_
rlabel metal2 6440 9660 6440 9660 0 _0958_
rlabel metal2 8232 9296 8232 9296 0 _0959_
rlabel metal2 7896 11256 7896 11256 0 _0960_
rlabel metal2 5656 29904 5656 29904 0 _0961_
rlabel metal2 5936 30156 5936 30156 0 _0962_
rlabel metal2 7112 30044 7112 30044 0 _0963_
rlabel metal3 4312 30184 4312 30184 0 _0964_
rlabel metal2 8120 6160 8120 6160 0 _0965_
rlabel metal3 11172 7560 11172 7560 0 _0966_
rlabel metal2 2744 26208 2744 26208 0 _0967_
rlabel metal2 7392 31080 7392 31080 0 _0968_
rlabel metal2 6328 27804 6328 27804 0 _0969_
rlabel metal3 5236 31080 5236 31080 0 _0970_
rlabel metal2 3528 31674 3528 31674 0 _0971_
rlabel metal2 5992 28728 5992 28728 0 _0972_
rlabel metal2 4424 13048 4424 13048 0 _0973_
rlabel metal2 2987 27720 2987 27720 0 _0974_
rlabel metal2 5936 27160 5936 27160 0 _0975_
rlabel metal2 2744 27888 2744 27888 0 _0976_
rlabel metal3 5236 27048 5236 27048 0 _0977_
rlabel metal2 6440 26740 6440 26740 0 _0978_
rlabel metal2 6216 25802 6216 25802 0 _0979_
rlabel metal3 5236 24808 5236 24808 0 _0980_
rlabel metal2 5992 25788 5992 25788 0 _0981_
rlabel metal2 3416 20888 3416 20888 0 _0982_
rlabel metal2 2408 22288 2408 22288 0 _0983_
rlabel metal2 4200 22792 4200 22792 0 _0984_
rlabel metal2 3640 23212 3640 23212 0 _0985_
rlabel metal2 3080 26047 3080 26047 0 _0986_
rlabel metal2 2744 20992 2744 20992 0 _0987_
rlabel metal2 3752 20818 3752 20818 0 _0988_
rlabel metal2 4088 20384 4088 20384 0 _0989_
rlabel metal2 3528 20692 3528 20692 0 _0990_
rlabel metal2 3864 18592 3864 18592 0 _0991_
rlabel metal3 4284 22568 4284 22568 0 _0992_
rlabel metal3 6020 23240 6020 23240 0 _0993_
rlabel metal3 6608 19992 6608 19992 0 _0994_
rlabel metal2 2408 19320 2408 19320 0 _0995_
rlabel metal2 6683 21504 6683 21504 0 _0996_
rlabel metal2 6272 21672 6272 21672 0 _0997_
rlabel metal2 7280 17640 7280 17640 0 _0998_
rlabel metal2 7112 18331 7112 18331 0 _0999_
rlabel metal2 7336 18984 7336 18984 0 _1000_
rlabel metal2 7448 18508 7448 18508 0 _1001_
rlabel metal2 4872 14224 4872 14224 0 _1002_
rlabel metal2 4760 18900 4760 18900 0 _1003_
rlabel metal2 4424 18312 4424 18312 0 _1004_
rlabel metal2 3080 18480 3080 18480 0 _1005_
rlabel via2 5096 16869 5096 16869 0 _1006_
rlabel metal2 6216 17584 6216 17584 0 _1007_
rlabel metal2 5432 17192 5432 17192 0 _1008_
rlabel metal2 5320 16548 5320 16548 0 _1009_
rlabel metal2 3528 15960 3528 15960 0 _1010_
rlabel metal2 5040 16352 5040 16352 0 _1011_
rlabel metal2 4648 15372 4648 15372 0 _1012_
rlabel metal2 7000 14770 7000 14770 0 _1013_
rlabel metal2 8344 17688 8344 17688 0 _1014_
rlabel metal2 8456 17164 8456 17164 0 _1015_
rlabel metal2 9464 16912 9464 16912 0 _1016_
rlabel metal2 6440 14672 6440 14672 0 _1017_
rlabel metal2 7616 14812 7616 14812 0 _1018_
rlabel metal2 5992 13258 5992 13258 0 _1019_
rlabel metal2 7672 12264 7672 12264 0 _1020_
rlabel metal2 8120 12880 8120 12880 0 _1021_
rlabel metal3 4760 12936 4760 12936 0 _1022_
rlabel metal2 10472 10920 10472 10920 0 _1023_
rlabel metal2 9016 12656 9016 12656 0 _1024_
rlabel metal2 7840 13328 7840 13328 0 _1025_
rlabel metal3 9408 13720 9408 13720 0 _1026_
rlabel metal2 12152 13622 12152 13622 0 _1027_
rlabel metal2 13216 12320 13216 12320 0 _1028_
rlabel metal2 11928 14504 11928 14504 0 _1029_
rlabel metal2 12376 11404 12376 11404 0 _1030_
rlabel metal2 12600 11088 12600 11088 0 _1031_
rlabel metal2 12488 8316 12488 8316 0 _1032_
rlabel metal2 10136 10261 10136 10261 0 _1033_
rlabel metal2 5096 11172 5096 11172 0 _1034_
rlabel metal3 9072 10584 9072 10584 0 _1035_
rlabel metal2 5656 6552 5656 6552 0 _1036_
rlabel metal2 4312 11572 4312 11572 0 _1037_
rlabel metal3 5348 10584 5348 10584 0 _1038_
rlabel metal3 3360 11368 3360 11368 0 _1039_
rlabel metal2 3528 11032 3528 11032 0 _1040_
rlabel metal2 4424 8297 4424 8297 0 _1041_
rlabel metal3 3192 9800 3192 9800 0 _1042_
rlabel metal3 5516 9016 5516 9016 0 _1043_
rlabel metal2 6328 8316 6328 8316 0 _1044_
rlabel metal2 5152 8344 5152 8344 0 _1045_
rlabel metal2 5992 6580 5992 6580 0 _1046_
rlabel metal2 6944 6580 6944 6580 0 _1047_
rlabel metal2 6272 5880 6272 5880 0 _1048_
rlabel metal2 6328 6720 6328 6720 0 _1049_
rlabel metal3 4312 6664 4312 6664 0 _1050_
rlabel metal2 6104 5824 6104 5824 0 _1051_
rlabel metal2 5096 6664 5096 6664 0 _1052_
rlabel via2 7896 5088 7896 5088 0 _1053_
rlabel metal2 4760 5992 4760 5992 0 _1054_
rlabel metal2 7336 5824 7336 5824 0 _1055_
rlabel metal2 8680 5152 8680 5152 0 _1056_
rlabel metal2 8456 5368 8456 5368 0 _1057_
rlabel metal2 8288 6132 8288 6132 0 _1058_
rlabel metal2 8008 7588 8008 7588 0 _1059_
rlabel metal2 8120 7243 8120 7243 0 _1060_
rlabel metal2 8820 5992 8820 5992 0 _1061_
rlabel metal2 10808 7125 10808 7125 0 _1062_
rlabel metal2 10024 7007 10024 7007 0 _1063_
rlabel metal2 11256 7448 11256 7448 0 _1064_
rlabel metal2 11088 5880 11088 5880 0 _1065_
rlabel metal3 20496 26152 20496 26152 0 _1066_
rlabel metal2 12908 34328 12908 34328 0 _1067_
rlabel metal2 31976 28616 31976 28616 0 _1068_
rlabel metal2 32536 28258 32536 28258 0 _1069_
rlabel metal2 31080 28196 31080 28196 0 _1070_
rlabel metal2 34328 29876 34328 29876 0 _1071_
rlabel metal2 37800 28876 37800 28876 0 _1072_
rlabel metal2 35896 29456 35896 29456 0 _1073_
rlabel metal2 34216 29652 34216 29652 0 _1074_
rlabel metal2 25452 23352 25452 23352 0 _1075_
rlabel metal2 15848 21924 15848 21924 0 _1076_
rlabel metal2 42224 19992 42224 19992 0 _1077_
rlabel metal2 41888 19992 41888 19992 0 _1078_
rlabel metal2 23128 21112 23128 21112 0 _1079_
rlabel metal3 23856 18424 23856 18424 0 _1080_
rlabel metal2 21896 20986 21896 20986 0 _1081_
rlabel metal2 16072 21868 16072 21868 0 _1082_
rlabel metal2 16576 21896 16576 21896 0 _1083_
rlabel metal2 10528 29064 10528 29064 0 _1084_
rlabel metal2 10248 21840 10248 21840 0 _1085_
rlabel metal2 13216 31192 13216 31192 0 _1086_
rlabel metal2 13552 22848 13552 22848 0 _1087_
rlabel metal3 11760 29064 11760 29064 0 _1088_
rlabel metal2 10920 22232 10920 22232 0 _1089_
rlabel metal2 37576 21504 37576 21504 0 _1090_
rlabel metal2 20552 39508 20552 39508 0 _1091_
rlabel metal2 21420 21000 21420 21000 0 _1092_
rlabel metal2 31752 30072 31752 30072 0 _1093_
rlabel metal2 10388 31192 10388 31192 0 _1094_
rlabel metal2 10920 33012 10920 33012 0 _1095_
rlabel metal2 42504 24136 42504 24136 0 _1096_
rlabel metal2 10780 31528 10780 31528 0 _1097_
rlabel metal2 10696 32732 10696 32732 0 _1098_
rlabel metal3 9660 33544 9660 33544 0 _1099_
rlabel metal2 9380 35672 9380 35672 0 _1100_
rlabel metal2 6216 34664 6216 34664 0 _1101_
rlabel metal2 10836 34104 10836 34104 0 _1102_
rlabel metal2 24808 21056 24808 21056 0 _1103_
rlabel metal2 37464 5768 37464 5768 0 _1104_
rlabel metal2 37912 4620 37912 4620 0 _1105_
rlabel metal2 38136 5152 38136 5152 0 _1106_
rlabel metal2 38248 4788 38248 4788 0 _1107_
rlabel metal2 37184 7168 37184 7168 0 _1108_
rlabel metal2 38248 8176 38248 8176 0 _1109_
rlabel metal3 35308 8232 35308 8232 0 _1110_
rlabel metal2 37072 7112 37072 7112 0 _1111_
rlabel metal2 39704 6160 39704 6160 0 _1112_
rlabel metal2 39312 5628 39312 5628 0 _1113_
rlabel metal2 37968 6944 37968 6944 0 _1114_
rlabel metal2 38444 8232 38444 8232 0 _1115_
rlabel metal3 37968 13048 37968 13048 0 _1116_
rlabel metal2 38584 11648 38584 11648 0 _1117_
rlabel metal2 37576 8456 37576 8456 0 _1118_
rlabel metal2 39368 10541 39368 10541 0 _1119_
rlabel metal2 39256 12488 39256 12488 0 _1120_
rlabel metal2 39592 10948 39592 10948 0 _1121_
rlabel metal2 36568 11648 36568 11648 0 _1122_
rlabel metal2 36092 8232 36092 8232 0 _1123_
rlabel metal2 36316 10024 36316 10024 0 _1124_
rlabel metal2 36092 11256 36092 11256 0 _1125_
rlabel metal2 35840 8232 35840 8232 0 _1126_
rlabel metal2 34832 7448 34832 7448 0 _1127_
rlabel metal2 34384 10864 34384 10864 0 _1128_
rlabel metal2 35000 10311 35000 10311 0 _1129_
rlabel metal2 34832 5880 34832 5880 0 _1130_
rlabel metal2 35980 7448 35980 7448 0 _1131_
rlabel metal2 35000 6350 35000 6350 0 _1132_
rlabel metal2 25592 18480 25592 18480 0 _1133_
rlabel metal2 28952 8176 28952 8176 0 _1134_
rlabel metal2 30296 5824 30296 5824 0 _1135_
rlabel metal3 33208 5768 33208 5768 0 _1136_
rlabel metal2 32732 5880 32732 5880 0 _1137_
rlabel metal2 31416 4480 31416 4480 0 _1138_
rlabel metal2 35448 3640 35448 3640 0 _1139_
rlabel metal3 32116 6664 32116 6664 0 _1140_
rlabel metal2 22792 21392 22792 21392 0 _1141_
rlabel metal2 22904 19656 22904 19656 0 _1142_
rlabel metal2 43624 13216 43624 13216 0 _1143_
rlabel metal3 39312 9016 39312 9016 0 _1144_
rlabel metal2 44968 11200 44968 11200 0 _1145_
rlabel metal3 42084 12824 42084 12824 0 _1146_
rlabel metal2 44744 8918 44744 8918 0 _1147_
rlabel metal2 48720 9016 48720 9016 0 _1148_
rlabel metal3 42196 9800 42196 9800 0 _1149_
rlabel metal2 41944 9856 41944 9856 0 _1150_
rlabel metal2 45528 8148 45528 8148 0 _1151_
rlabel metal3 42140 9016 42140 9016 0 _1152_
rlabel metal2 39536 9352 39536 9352 0 _1153_
rlabel metal2 43176 3528 43176 3528 0 _1154_
rlabel metal2 44128 6104 44128 6104 0 _1155_
rlabel metal3 45892 3528 45892 3528 0 _1156_
rlabel metal2 45304 7532 45304 7532 0 _1157_
rlabel metal2 48216 5138 48216 5138 0 _1158_
rlabel metal2 48608 3528 48608 3528 0 _1159_
rlabel metal2 48664 15204 48664 15204 0 _1160_
rlabel metal2 48664 4648 48664 4648 0 _1161_
rlabel metal2 47432 4872 47432 4872 0 _1162_
rlabel metal2 46116 8120 46116 8120 0 _1163_
rlabel metal2 31248 7224 31248 7224 0 _1164_
rlabel metal3 31276 7448 31276 7448 0 _1165_
rlabel metal2 31024 9016 31024 9016 0 _1166_
rlabel metal2 30296 6552 30296 6552 0 _1167_
rlabel metal2 30968 6216 30968 6216 0 _1168_
rlabel metal2 29624 6384 29624 6384 0 _1169_
rlabel metal3 30072 3640 30072 3640 0 _1170_
rlabel metal2 28224 4984 28224 4984 0 _1171_
rlabel metal2 27944 5040 27944 5040 0 _1172_
rlabel metal2 19096 6440 19096 6440 0 _1173_
rlabel metal2 20776 5152 20776 5152 0 _1174_
rlabel metal3 17948 4200 17948 4200 0 _1175_
rlabel metal2 18536 4396 18536 4396 0 _1176_
rlabel metal2 16240 4396 16240 4396 0 _1177_
rlabel metal2 16828 5656 16828 5656 0 _1178_
rlabel metal2 15400 5656 15400 5656 0 _1179_
rlabel metal2 17416 6048 17416 6048 0 _1180_
rlabel metal3 17668 6552 17668 6552 0 _1181_
rlabel metal2 17304 7756 17304 7756 0 _1182_
rlabel metal2 19432 6700 19432 6700 0 _1183_
rlabel metal3 20104 6664 20104 6664 0 _1184_
rlabel metal2 19544 7084 19544 7084 0 _1185_
rlabel metal2 21168 5096 21168 5096 0 _1186_
rlabel metal3 30240 14504 30240 14504 0 _1187_
rlabel metal2 31584 14616 31584 14616 0 _1188_
rlabel metal3 30072 15624 30072 15624 0 _1189_
rlabel metal3 31864 14504 31864 14504 0 _1190_
rlabel metal2 29680 16184 29680 16184 0 _1191_
rlabel metal2 30520 13208 30520 13208 0 _1192_
rlabel metal2 29736 16856 29736 16856 0 _1193_
rlabel metal2 29736 12978 29736 12978 0 _1194_
rlabel metal2 29400 12824 29400 12824 0 _1195_
rlabel metal3 28784 12936 28784 12936 0 _1196_
rlabel metal2 29624 11404 29624 11404 0 _1197_
rlabel metal2 29148 10696 29148 10696 0 _1198_
rlabel metal3 28728 10584 28728 10584 0 _1199_
rlabel metal3 29344 9016 29344 9016 0 _1200_
rlabel metal2 27832 8036 27832 8036 0 _1201_
rlabel metal3 28952 7448 28952 7448 0 _1202_
rlabel metal2 27776 9800 27776 9800 0 _1203_
rlabel metal2 27496 6720 27496 6720 0 _1204_
rlabel metal2 28672 7000 28672 7000 0 _1205_
rlabel metal2 26600 7952 26600 7952 0 _1206_
rlabel metal2 25480 6720 25480 6720 0 _1207_
rlabel metal2 24024 7392 24024 7392 0 _1208_
rlabel metal3 23688 6664 23688 6664 0 _1209_
rlabel metal2 24248 4984 24248 4984 0 _1210_
rlabel metal3 28224 30968 28224 30968 0 _1211_
rlabel metal2 21000 38942 21000 38942 0 _1212_
rlabel metal2 12712 35532 12712 35532 0 _1213_
rlabel metal2 21336 39032 21336 39032 0 _1214_
rlabel metal2 20328 39144 20328 39144 0 _1215_
rlabel metal2 14952 35042 14952 35042 0 _1216_
rlabel metal2 14476 35112 14476 35112 0 _1217_
rlabel metal2 18872 35728 18872 35728 0 _1218_
rlabel metal2 11956 36456 11956 36456 0 _1219_
rlabel metal2 11984 34104 11984 34104 0 _1220_
rlabel metal2 20440 39452 20440 39452 0 _1221_
rlabel metal2 20216 39508 20216 39508 0 _1222_
rlabel metal2 19628 39816 19628 39816 0 _1223_
rlabel metal3 21952 43736 21952 43736 0 _1224_
rlabel metal2 19600 45640 19600 45640 0 _1225_
rlabel metal2 20552 44334 20552 44334 0 _1226_
rlabel metal2 19572 44296 19572 44296 0 _1227_
rlabel via1 20757 42000 20757 42000 0 _1228_
rlabel metal2 19824 42112 19824 42112 0 _1229_
rlabel metal3 33600 27832 33600 27832 0 _1230_
rlabel metal2 31864 30016 31864 30016 0 _1231_
rlabel metal2 15624 24752 15624 24752 0 _1232_
rlabel metal2 15288 24976 15288 24976 0 _1233_
rlabel metal2 14280 24584 14280 24584 0 _1234_
rlabel metal2 14700 26264 14700 26264 0 _1235_
rlabel metal2 12124 24136 12124 24136 0 _1236_
rlabel metal2 11536 25984 11536 25984 0 _1237_
rlabel metal3 9660 24696 9660 24696 0 _1238_
rlabel metal2 26152 29540 26152 29540 0 _1239_
rlabel metal2 25648 32536 25648 32536 0 _1240_
rlabel metal3 25648 26600 25648 26600 0 _1241_
rlabel metal2 24304 30968 24304 30968 0 _1242_
rlabel metal2 25984 26152 25984 26152 0 _1243_
rlabel metal2 26824 30240 26824 30240 0 _1244_
rlabel metal2 26675 23212 26675 23212 0 _1245_
rlabel metal2 24808 30072 24808 30072 0 _1246_
rlabel via2 25256 26281 25256 26281 0 _1247_
rlabel metal2 26096 26628 26096 26628 0 _1248_
rlabel metal2 26600 28878 26600 28878 0 _1249_
rlabel metal2 26824 28672 26824 28672 0 _1250_
rlabel metal3 24976 32760 24976 32760 0 _1251_
rlabel metal2 22904 33418 22904 33418 0 _1252_
rlabel metal3 22652 31976 22652 31976 0 _1253_
rlabel metal2 22372 33544 22372 33544 0 _1254_
rlabel metal2 25144 34440 25144 34440 0 _1255_
rlabel metal2 26124 31752 26124 31752 0 _1256_
rlabel metal2 47208 12936 47208 12936 0 _1257_
rlabel metal2 47432 12109 47432 12109 0 _1258_
rlabel metal2 48888 14336 48888 14336 0 _1259_
rlabel metal2 47880 12236 47880 12236 0 _1260_
rlabel metal3 47488 14840 47488 14840 0 _1261_
rlabel metal2 45211 14420 45211 14420 0 _1262_
rlabel metal2 47656 16296 47656 16296 0 _1263_
rlabel metal2 43960 12984 43960 12984 0 _1264_
rlabel via2 41944 12928 41944 12928 0 _1265_
rlabel metal2 30968 11404 30968 11404 0 _1266_
rlabel metal2 31192 11312 31192 11312 0 _1267_
rlabel metal2 31080 9800 31080 9800 0 _1268_
rlabel metal2 26658 17444 26658 17444 0 _1269_
rlabel metal2 35168 14504 35168 14504 0 _1270_
rlabel metal3 12376 8176 12376 8176 0 blink.LED
rlabel metal2 4760 30044 4760 30044 0 blink.counter\[0\]
rlabel metal3 3192 21224 3192 21224 0 blink.counter\[10\]
rlabel metal3 8232 20776 8232 20776 0 blink.counter\[11\]
rlabel metal2 9016 19656 9016 19656 0 blink.counter\[12\]
rlabel metal2 5768 15680 5768 15680 0 blink.counter\[13\]
rlabel metal2 5880 16576 5880 16576 0 blink.counter\[14\]
rlabel metal2 3192 16016 3192 16016 0 blink.counter\[15\]
rlabel metal2 8568 16632 8568 16632 0 blink.counter\[16\]
rlabel metal3 10192 14616 10192 14616 0 blink.counter\[17\]
rlabel metal3 7168 13720 7168 13720 0 blink.counter\[18\]
rlabel metal2 8344 12544 8344 12544 0 blink.counter\[19\]
rlabel metal2 5096 30016 5096 30016 0 blink.counter\[1\]
rlabel metal2 13832 14168 13832 14168 0 blink.counter\[20\]
rlabel metal2 11928 11885 11928 11885 0 blink.counter\[21\]
rlabel metal2 11256 11200 11256 11200 0 blink.counter\[22\]
rlabel metal2 5320 10640 5320 10640 0 blink.counter\[23\]
rlabel metal2 4312 10752 4312 10752 0 blink.counter\[24\]
rlabel metal2 4760 8316 4760 8316 0 blink.counter\[25\]
rlabel metal2 7112 6776 7112 6776 0 blink.counter\[26\]
rlabel metal2 5824 5096 5824 5096 0 blink.counter\[27\]
rlabel metal2 7896 5656 7896 5656 0 blink.counter\[28\]
rlabel metal3 10528 8120 10528 8120 0 blink.counter\[29\]
rlabel metal3 4760 30968 4760 30968 0 blink.counter\[2\]
rlabel metal3 9912 5880 9912 5880 0 blink.counter\[30\]
rlabel metal3 9619 9800 9619 9800 0 blink.counter\[31\]
rlabel metal2 4984 31080 4984 31080 0 blink.counter\[3\]
rlabel metal3 6944 27832 6944 27832 0 blink.counter\[4\]
rlabel metal2 4312 27496 4312 27496 0 blink.counter\[5\]
rlabel metal2 5432 25032 5432 25032 0 blink.counter\[6\]
rlabel metal2 4312 23632 4312 23632 0 blink.counter\[7\]
rlabel metal3 2352 24696 2352 24696 0 blink.counter\[8\]
rlabel metal2 3080 20888 3080 20888 0 blink.counter\[9\]
rlabel metal2 17836 19320 17836 19320 0 clknet_0_wb_clk_i
rlabel metal2 7252 8344 7252 8344 0 clknet_2_0__leaf_wb_clk_i
rlabel metal2 7560 29357 7560 29357 0 clknet_2_1__leaf_wb_clk_i
rlabel metal2 29176 12277 29176 12277 0 clknet_2_2__leaf_wb_clk_i
rlabel metal2 45864 46522 45864 46522 0 clknet_2_3__leaf_wb_clk_i
rlabel metal3 10640 15064 10640 15064 0 clknet_leaf_0_wb_clk_i
rlabel metal2 16072 43232 16072 43232 0 clknet_leaf_10_wb_clk_i
rlabel metal3 24360 44296 24360 44296 0 clknet_leaf_11_wb_clk_i
rlabel metal3 23968 40376 23968 40376 0 clknet_leaf_12_wb_clk_i
rlabel metal2 21784 32480 21784 32480 0 clknet_leaf_13_wb_clk_i
rlabel metal3 26152 33320 26152 33320 0 clknet_leaf_14_wb_clk_i
rlabel metal3 33992 35896 33992 35896 0 clknet_leaf_15_wb_clk_i
rlabel metal2 26488 41440 26488 41440 0 clknet_leaf_16_wb_clk_i
rlabel metal2 36344 46256 36344 46256 0 clknet_leaf_17_wb_clk_i
rlabel metal2 36624 41944 36624 41944 0 clknet_leaf_18_wb_clk_i
rlabel metal2 43848 47712 43848 47712 0 clknet_leaf_19_wb_clk_i
rlabel metal2 1624 22736 1624 22736 0 clknet_leaf_1_wb_clk_i
rlabel metal2 46368 44744 46368 44744 0 clknet_leaf_20_wb_clk_i
rlabel metal3 41608 37240 41608 37240 0 clknet_leaf_21_wb_clk_i
rlabel metal2 49392 33320 49392 33320 0 clknet_leaf_22_wb_clk_i
rlabel metal2 41384 27440 41384 27440 0 clknet_leaf_23_wb_clk_i
rlabel metal2 38136 34216 38136 34216 0 clknet_leaf_24_wb_clk_i
rlabel metal3 26264 25480 26264 25480 0 clknet_leaf_25_wb_clk_i
rlabel metal3 35000 21560 35000 21560 0 clknet_leaf_26_wb_clk_i
rlabel metal2 41496 20776 41496 20776 0 clknet_leaf_27_wb_clk_i
rlabel metal2 49000 22512 49000 22512 0 clknet_leaf_28_wb_clk_i
rlabel metal3 46200 15512 46200 15512 0 clknet_leaf_29_wb_clk_i
rlabel metal3 6272 25480 6272 25480 0 clknet_leaf_2_wb_clk_i
rlabel metal3 48776 9800 48776 9800 0 clknet_leaf_30_wb_clk_i
rlabel metal2 41104 6664 41104 6664 0 clknet_leaf_31_wb_clk_i
rlabel metal2 38584 5376 38584 5376 0 clknet_leaf_32_wb_clk_i
rlabel metal3 37464 11368 37464 11368 0 clknet_leaf_33_wb_clk_i
rlabel metal2 31192 4816 31192 4816 0 clknet_leaf_34_wb_clk_i
rlabel metal2 29288 8316 29288 8316 0 clknet_leaf_35_wb_clk_i
rlabel via2 28280 16072 28280 16072 0 clknet_leaf_36_wb_clk_i
rlabel metal2 25144 22736 25144 22736 0 clknet_leaf_37_wb_clk_i
rlabel metal2 19880 15960 19880 15960 0 clknet_leaf_38_wb_clk_i
rlabel metal3 20776 7448 20776 7448 0 clknet_leaf_39_wb_clk_i
rlabel metal2 14056 17640 14056 17640 0 clknet_leaf_3_wb_clk_i
rlabel metal2 14056 6272 14056 6272 0 clknet_leaf_40_wb_clk_i
rlabel metal2 13384 6944 13384 6944 0 clknet_leaf_41_wb_clk_i
rlabel metal3 6664 7672 6664 7672 0 clknet_leaf_42_wb_clk_i
rlabel metal2 2744 12656 2744 12656 0 clknet_leaf_43_wb_clk_i
rlabel metal2 20440 23016 20440 23016 0 clknet_leaf_4_wb_clk_i
rlabel metal2 9352 29792 9352 29792 0 clknet_leaf_5_wb_clk_i
rlabel metal2 1960 29456 1960 29456 0 clknet_leaf_6_wb_clk_i
rlabel metal2 5544 33320 5544 33320 0 clknet_leaf_7_wb_clk_i
rlabel metal2 10304 38584 10304 38584 0 clknet_leaf_8_wb_clk_i
rlabel metal3 9352 44296 9352 44296 0 clknet_leaf_9_wb_clk_i
rlabel metal2 44380 39368 44380 39368 0 custom_settings[0]
rlabel metal2 47208 43512 47208 43512 0 custom_settings[1]
rlabel metal2 49336 47544 49336 47544 0 custom_settings[3]
rlabel metal3 47474 2072 47474 2072 0 io_in_1[0]
rlabel metal2 21840 23912 21840 23912 0 io_in_1[1]
rlabel metal2 44016 21336 44016 21336 0 io_in_1[2]
rlabel metal2 39200 24360 39200 24360 0 io_in_1[3]
rlabel metal2 49392 16856 49392 16856 0 io_in_1[4]
rlabel metal3 49826 23352 49826 23352 0 io_in_1[5]
rlabel metal2 49336 27720 49336 27720 0 io_in_1[6]
rlabel metal3 46508 34104 46508 34104 0 io_in_1[7]
rlabel metal2 31976 46648 31976 46648 0 io_in_2[0]
rlabel metal2 47320 47768 47320 47768 0 io_in_2[1]
rlabel metal3 19712 5656 19712 5656 0 io_out[10]
rlabel metal3 21504 3640 21504 3640 0 io_out[11]
rlabel metal2 31640 2142 31640 2142 0 io_out[17]
rlabel metal2 33432 2198 33432 2198 0 io_out[18]
rlabel metal2 35224 2254 35224 2254 0 io_out[19]
rlabel metal2 37016 2086 37016 2086 0 io_out[20]
rlabel metal2 38808 1638 38808 1638 0 io_out[21]
rlabel metal2 15512 2030 15512 2030 0 io_out[8]
rlabel metal3 17920 5096 17920 5096 0 io_out[9]
rlabel metal2 45472 19376 45472 19376 0 net1
rlabel metal2 19040 47208 19040 47208 0 net10
rlabel metal2 19040 6104 19040 6104 0 net11
rlabel metal2 21448 3626 21448 3626 0 net12
rlabel metal2 34664 3738 34664 3738 0 net13
rlabel metal2 36232 4970 36232 4970 0 net14
rlabel metal2 37912 5557 37912 5557 0 net15
rlabel metal2 41720 6832 41720 6832 0 net16
rlabel metal2 37688 6832 37688 6832 0 net17
rlabel metal2 14056 3794 14056 3794 0 net18
rlabel metal2 15400 4704 15400 4704 0 net19
rlabel metal3 46480 43288 46480 43288 0 net2
rlabel metal2 1176 2086 1176 2086 0 net20
rlabel metal2 2968 2030 2968 2030 0 net21
rlabel metal2 4760 2086 4760 2086 0 net22
rlabel metal2 6552 2030 6552 2030 0 net23
rlabel metal2 8344 2030 8344 2030 0 net24
rlabel metal2 10136 2030 10136 2030 0 net25
rlabel metal2 11928 2030 11928 2030 0 net26
rlabel metal2 13720 2030 13720 2030 0 net27
rlabel metal2 20160 3388 20160 3388 0 net28
rlabel metal2 24472 1750 24472 1750 0 net29
rlabel metal2 49000 47152 49000 47152 0 net3
rlabel metal2 26432 2968 26432 2968 0 net30
rlabel metal2 28056 2030 28056 2030 0 net31
rlabel metal2 29848 2086 29848 2086 0 net32
rlabel metal3 43960 4760 43960 4760 0 net33
rlabel metal3 46676 4872 46676 4872 0 net34
rlabel metal3 44968 3976 44968 3976 0 net35
rlabel metal2 48160 8876 48160 8876 0 net36
rlabel metal2 49364 9576 49364 9576 0 net37
rlabel metal2 40768 2184 40768 2184 0 net38
rlabel metal2 40432 18088 40432 18088 0 net4
rlabel metal2 44408 29484 44408 29484 0 net5
rlabel metal2 44856 29988 44856 29988 0 net6
rlabel metal2 40264 34048 40264 34048 0 net7
rlabel metal2 33040 42504 33040 42504 0 net8
rlabel metal3 45164 28056 45164 28056 0 net9
rlabel metal2 19068 47544 19068 47544 0 rst_n
rlabel metal2 47264 3528 47264 3528 0 tt_um_rejunity_ay8913.DAC_clk
rlabel metal2 43736 10696 43736 10696 0 tt_um_rejunity_ay8913.DAC_dat
rlabel metal2 36344 5936 36344 5936 0 tt_um_rejunity_ay8913.DAC_le
rlabel metal2 38920 28224 38920 28224 0 tt_um_rejunity_ay8913.active
rlabel metal2 28392 19782 28392 19782 0 tt_um_rejunity_ay8913.amplitude_A\[0\]
rlabel via2 27944 22330 27944 22330 0 tt_um_rejunity_ay8913.amplitude_B\[0\]
rlabel metal2 33824 19096 33824 19096 0 tt_um_rejunity_ay8913.amplitude_C\[0\]
rlabel metal2 39816 19432 39816 19432 0 tt_um_rejunity_ay8913.clk_counter\[0\]
rlabel metal2 40656 20664 40656 20664 0 tt_um_rejunity_ay8913.clk_counter\[1\]
rlabel metal2 41048 18088 41048 18088 0 tt_um_rejunity_ay8913.clk_counter\[2\]
rlabel metal3 41888 16856 41888 16856 0 tt_um_rejunity_ay8913.clk_counter\[3\]
rlabel metal2 44072 16632 44072 16632 0 tt_um_rejunity_ay8913.clk_counter\[4\]
rlabel metal3 45976 17640 45976 17640 0 tt_um_rejunity_ay8913.clk_counter\[5\]
rlabel via1 44072 18431 44072 18431 0 tt_um_rejunity_ay8913.clk_counter\[6\]
rlabel metal2 30408 19880 30408 19880 0 tt_um_rejunity_ay8913.envelope_A
rlabel metal2 30520 21392 30520 21392 0 tt_um_rejunity_ay8913.envelope_B
rlabel via2 33656 18438 33656 18438 0 tt_um_rejunity_ay8913.envelope_C
rlabel metal3 40320 25480 40320 25480 0 tt_um_rejunity_ay8913.envelope_alternate
rlabel metal3 39928 22456 39928 22456 0 tt_um_rejunity_ay8913.envelope_attack
rlabel metal3 41888 26376 41888 26376 0 tt_um_rejunity_ay8913.envelope_continue
rlabel metal2 48664 21448 48664 21448 0 tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[0\]
rlabel metal3 47880 19992 47880 19992 0 tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[1\]
rlabel metal2 48104 24024 48104 24024 0 tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[2\]
rlabel metal2 47712 26264 47712 26264 0 tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[3\]
rlabel metal2 42616 25424 42616 25424 0 tt_um_rejunity_ay8913.envelope_generator.hold
rlabel metal3 43792 22232 43792 22232 0 tt_um_rejunity_ay8913.envelope_generator.invert_output
rlabel metal2 38472 32984 38472 32984 0 tt_um_rejunity_ay8913.envelope_generator.period\[0\]
rlabel metal2 41812 42028 41812 42028 0 tt_um_rejunity_ay8913.envelope_generator.period\[10\]
rlabel metal2 40264 40656 40264 40656 0 tt_um_rejunity_ay8913.envelope_generator.period\[11\]
rlabel metal2 44968 44128 44968 44128 0 tt_um_rejunity_ay8913.envelope_generator.period\[12\]
rlabel metal2 44744 44548 44744 44548 0 tt_um_rejunity_ay8913.envelope_generator.period\[13\]
rlabel metal2 44744 42742 44744 42742 0 tt_um_rejunity_ay8913.envelope_generator.period\[14\]
rlabel via2 44520 40390 44520 40390 0 tt_um_rejunity_ay8913.envelope_generator.period\[15\]
rlabel metal2 39032 32760 39032 32760 0 tt_um_rejunity_ay8913.envelope_generator.period\[1\]
rlabel via1 41534 30976 41534 30976 0 tt_um_rejunity_ay8913.envelope_generator.period\[2\]
rlabel metal2 42056 32648 42056 32648 0 tt_um_rejunity_ay8913.envelope_generator.period\[3\]
rlabel via2 43176 28602 43176 28602 0 tt_um_rejunity_ay8913.envelope_generator.period\[4\]
rlabel metal3 45528 32536 45528 32536 0 tt_um_rejunity_ay8913.envelope_generator.period\[5\]
rlabel metal2 45416 30954 45416 30954 0 tt_um_rejunity_ay8913.envelope_generator.period\[6\]
rlabel metal3 44632 30856 44632 30856 0 tt_um_rejunity_ay8913.envelope_generator.period\[7\]
rlabel metal2 41832 40432 41832 40432 0 tt_um_rejunity_ay8913.envelope_generator.period\[8\]
rlabel metal2 40824 40040 40824 40040 0 tt_um_rejunity_ay8913.envelope_generator.period\[9\]
rlabel metal3 48608 29400 48608 29400 0 tt_um_rejunity_ay8913.envelope_generator.signal_edge.previous_signal_state_0
rlabel metal2 47096 38741 47096 38741 0 tt_um_rejunity_ay8913.envelope_generator.signal_edge.signal
rlabel metal2 46312 26544 46312 26544 0 tt_um_rejunity_ay8913.envelope_generator.stop
rlabel metal2 34104 34804 34104 34804 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[0\]
rlabel metal2 40936 42224 40936 42224 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[10\]
rlabel metal2 41272 45696 41272 45696 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[11\]
rlabel metal2 48104 46480 48104 46480 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[12\]
rlabel via2 45752 45097 45752 45097 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[13\]
rlabel metal2 45192 44072 45192 44072 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[14\]
rlabel metal3 47768 41048 47768 41048 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[15\]
rlabel metal2 39088 34188 39088 34188 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[1\]
rlabel metal3 41664 34888 41664 34888 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[2\]
rlabel metal2 39928 36008 39928 36008 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[3\]
rlabel metal2 46648 35392 46648 35392 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[4\]
rlabel metal2 49168 34776 49168 34776 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[5\]
rlabel metal2 45640 34720 45640 34720 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[6\]
rlabel metal2 45080 39200 45080 39200 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[7\]
rlabel metal2 43568 38696 43568 38696 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[8\]
rlabel metal2 43176 44744 43176 44744 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[9\]
rlabel metal2 30352 26376 30352 26376 0 tt_um_rejunity_ay8913.latched_register\[0\]
rlabel metal2 31304 28616 31304 28616 0 tt_um_rejunity_ay8913.latched_register\[1\]
rlabel metal2 33208 25760 33208 25760 0 tt_um_rejunity_ay8913.latched_register\[2\]
rlabel metal2 35336 26628 35336 26628 0 tt_um_rejunity_ay8913.latched_register\[3\]
rlabel metal2 29624 23324 29624 23324 0 tt_um_rejunity_ay8913.noise_disable_A
rlabel metal2 33432 21728 33432 21728 0 tt_um_rejunity_ay8913.noise_disable_B
rlabel metal2 35896 21812 35896 21812 0 tt_um_rejunity_ay8913.noise_disable_C
rlabel metal3 29512 16856 29512 16856 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[0\]
rlabel metal3 17248 9800 17248 9800 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[10\]
rlabel metal2 18088 9380 18088 9380 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[11\]
rlabel metal2 18312 8232 18312 8232 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[12\]
rlabel metal2 22120 8400 22120 8400 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[13\]
rlabel metal3 25928 10584 25928 10584 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[14\]
rlabel metal3 25816 11480 25816 11480 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[15\]
rlabel metal2 26600 11928 26600 11928 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[16\]
rlabel metal3 25088 15288 25088 15288 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[1\]
rlabel metal2 23688 15251 23688 15251 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[2\]
rlabel metal2 22792 16128 22792 16128 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[3\]
rlabel metal3 21672 15512 21672 15512 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[4\]
rlabel via2 19992 16061 19992 16061 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[5\]
rlabel metal2 16520 15736 16520 15736 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[6\]
rlabel metal2 16968 14420 16968 14420 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[7\]
rlabel metal2 16520 13860 16520 13860 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[8\]
rlabel metal2 16800 11368 16800 11368 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[9\]
rlabel metal2 16296 21644 16296 21644 0 tt_um_rejunity_ay8913.noise_generator.period\[0\]
rlabel via2 12376 22330 12376 22330 0 tt_um_rejunity_ay8913.noise_generator.period\[1\]
rlabel metal2 15176 21784 15176 21784 0 tt_um_rejunity_ay8913.noise_generator.period\[2\]
rlabel metal2 11984 20664 11984 20664 0 tt_um_rejunity_ay8913.noise_generator.period\[3\]
rlabel metal2 20944 20776 20944 20776 0 tt_um_rejunity_ay8913.noise_generator.period\[4\]
rlabel metal2 23240 18760 23240 18760 0 tt_um_rejunity_ay8913.noise_generator.signal_edge.previous_signal_state_0
rlabel metal2 22568 18648 22568 18648 0 tt_um_rejunity_ay8913.noise_generator.signal_edge.signal
rlabel metal2 16856 20160 16856 20160 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[0\]
rlabel metal2 12376 19432 12376 19432 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[1\]
rlabel metal2 16520 18256 16520 18256 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[2\]
rlabel metal2 15288 18872 15288 18872 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[3\]
rlabel metal2 16744 18200 16744 18200 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[4\]
rlabel metal2 32536 10584 32536 10584 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[2\]
rlabel metal2 34328 11592 34328 11592 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[3\]
rlabel metal2 33880 13776 33880 13776 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[4\]
rlabel metal2 35448 13832 35448 13832 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[5\]
rlabel metal2 36120 16016 36120 16016 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[6\]
rlabel metal2 39256 16520 39256 16520 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[7\]
rlabel metal2 39592 15204 39592 15204 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[8\]
rlabel metal3 23632 3640 23632 3640 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[9\]
rlabel metal3 32816 15288 32816 15288 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[2\]
rlabel metal2 30520 15456 30520 15456 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[3\]
rlabel metal3 30184 12936 30184 12936 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[4\]
rlabel metal2 28448 11256 28448 11256 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[5\]
rlabel metal2 28672 9128 28672 9128 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[6\]
rlabel metal2 28000 7448 28000 7448 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[7\]
rlabel metal2 24472 7896 24472 7896 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[8\]
rlabel metal2 23184 4312 23184 4312 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[9\]
rlabel metal2 31864 8680 31864 8680 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[2\]
rlabel metal3 30240 6664 30240 6664 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[3\]
rlabel metal2 29624 4480 29624 4480 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[4\]
rlabel metal3 19992 3640 19992 3640 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[5\]
rlabel metal2 16408 5600 16408 5600 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[6\]
rlabel metal3 17192 6664 17192 6664 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[7\]
rlabel metal2 20328 7784 20328 7784 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[8\]
rlabel metal2 22344 5152 22344 5152 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[9\]
rlabel metal3 29568 4312 29568 4312 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[10\]
rlabel metal2 38472 6384 38472 6384 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[2\]
rlabel metal3 38080 6664 38080 6664 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[3\]
rlabel metal2 37016 11536 37016 11536 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[4\]
rlabel metal2 38248 10920 38248 10920 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[5\]
rlabel metal2 38024 10472 38024 10472 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[6\]
rlabel metal2 33432 9352 33432 9352 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[7\]
rlabel metal2 35000 7280 35000 7280 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[8\]
rlabel metal2 33544 5544 33544 5544 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[9\]
rlabel metal2 42168 22960 42168 22960 0 tt_um_rejunity_ay8913.restart_envelope
rlabel metal2 47880 10864 47880 10864 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[0\]
rlabel metal2 46648 11767 46648 11767 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[1\]
rlabel metal2 49112 14728 49112 14728 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[2\]
rlabel metal2 45472 13608 45472 13608 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[3\]
rlabel metal2 45696 13020 45696 13020 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[4\]
rlabel metal2 45491 7532 45491 7532 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[10\]
rlabel metal2 45528 9968 45528 9968 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[11\]
rlabel metal2 44296 9100 44296 9100 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[2\]
rlabel metal3 43960 8344 43960 8344 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[3\]
rlabel metal2 43680 5992 43680 5992 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[4\]
rlabel metal2 44072 4928 44072 4928 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[5\]
rlabel metal2 44632 4592 44632 4592 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[6\]
rlabel metal3 45360 5208 45360 5208 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[7\]
rlabel via1 46256 3520 46256 3520 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[8\]
rlabel metal3 45640 6552 45640 6552 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[9\]
rlabel metal3 31808 24696 31808 24696 0 tt_um_rejunity_ay8913.tone_A
rlabel metal2 28840 38724 28840 38724 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[0\]
rlabel metal2 33432 44296 33432 44296 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[10\]
rlabel metal2 35952 44100 35952 44100 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[11\]
rlabel metal2 24024 37912 24024 37912 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[1\]
rlabel metal2 27104 40376 27104 40376 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[2\]
rlabel metal3 20776 40544 20776 40544 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[3\]
rlabel metal2 24360 42280 24360 42280 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[4\]
rlabel metal2 25032 44632 25032 44632 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[5\]
rlabel metal2 22904 47096 22904 47096 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[6\]
rlabel metal2 26600 46648 26600 46648 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[7\]
rlabel metal3 31696 46648 31696 46648 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[8\]
rlabel metal2 31752 44968 31752 44968 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[9\]
rlabel metal2 30688 38836 30688 38836 0 tt_um_rejunity_ay8913.tone_A_generator.period\[0\]
rlabel metal2 35784 31528 35784 31528 0 tt_um_rejunity_ay8913.tone_A_generator.period\[10\]
rlabel metal2 34944 41944 34944 41944 0 tt_um_rejunity_ay8913.tone_A_generator.period\[11\]
rlabel metal2 29848 36904 29848 36904 0 tt_um_rejunity_ay8913.tone_A_generator.period\[1\]
rlabel metal2 27990 40376 27990 40376 0 tt_um_rejunity_ay8913.tone_A_generator.period\[2\]
rlabel metal2 28672 40376 28672 40376 0 tt_um_rejunity_ay8913.tone_A_generator.period\[3\]
rlabel metal2 29288 41104 29288 41104 0 tt_um_rejunity_ay8913.tone_A_generator.period\[4\]
rlabel via2 32200 38822 32200 38822 0 tt_um_rejunity_ay8913.tone_A_generator.period\[5\]
rlabel metal2 28056 44506 28056 44506 0 tt_um_rejunity_ay8913.tone_A_generator.period\[6\]
rlabel via2 27720 42714 27720 42714 0 tt_um_rejunity_ay8913.tone_A_generator.period\[7\]
rlabel metal2 32760 43680 32760 43680 0 tt_um_rejunity_ay8913.tone_A_generator.period\[8\]
rlabel metal2 31752 41832 31752 41832 0 tt_um_rejunity_ay8913.tone_A_generator.period\[9\]
rlabel metal2 21112 23072 21112 23072 0 tt_um_rejunity_ay8913.tone_B
rlabel metal2 20552 31920 20552 31920 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[0\]
rlabel metal2 10136 27104 10136 27104 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[10\]
rlabel metal2 9800 27552 9800 27552 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[11\]
rlabel metal2 20888 31052 20888 31052 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[1\]
rlabel metal2 21840 26376 21840 26376 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[2\]
rlabel metal3 19432 25592 19432 25592 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[3\]
rlabel metal2 21336 29876 21336 29876 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[4\]
rlabel metal3 18592 33432 18592 33432 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[5\]
rlabel metal2 15736 33488 15736 33488 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[6\]
rlabel metal2 12320 30968 12320 30968 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[7\]
rlabel metal3 11648 30184 11648 30184 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[8\]
rlabel metal2 12488 27216 12488 27216 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[9\]
rlabel metal2 18984 31024 18984 31024 0 tt_um_rejunity_ay8913.tone_B_generator.period\[0\]
rlabel metal2 11816 26432 11816 26432 0 tt_um_rejunity_ay8913.tone_B_generator.period\[10\]
rlabel metal2 11144 26342 11144 26342 0 tt_um_rejunity_ay8913.tone_B_generator.period\[11\]
rlabel metal2 25312 30072 25312 30072 0 tt_um_rejunity_ay8913.tone_B_generator.period\[1\]
rlabel metal3 23128 25592 23128 25592 0 tt_um_rejunity_ay8913.tone_B_generator.period\[2\]
rlabel metal2 23106 26600 23106 26600 0 tt_um_rejunity_ay8913.tone_B_generator.period\[3\]
rlabel metal2 22680 31920 22680 31920 0 tt_um_rejunity_ay8913.tone_B_generator.period\[4\]
rlabel metal2 22680 33418 22680 33418 0 tt_um_rejunity_ay8913.tone_B_generator.period\[5\]
rlabel metal2 23800 33488 23800 33488 0 tt_um_rejunity_ay8913.tone_B_generator.period\[6\]
rlabel metal2 14616 30688 14616 30688 0 tt_um_rejunity_ay8913.tone_B_generator.period\[7\]
rlabel metal2 14000 30968 14000 30968 0 tt_um_rejunity_ay8913.tone_B_generator.period\[8\]
rlabel metal2 13944 24472 13944 24472 0 tt_um_rejunity_ay8913.tone_B_generator.period\[9\]
rlabel metal2 23688 23912 23688 23912 0 tt_um_rejunity_ay8913.tone_C
rlabel metal3 16744 38024 16744 38024 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[0\]
rlabel metal2 10136 38080 10136 38080 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[10\]
rlabel metal2 8680 38080 8680 38080 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[11\]
rlabel metal3 21056 38024 21056 38024 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[1\]
rlabel metal2 10976 41944 10976 41944 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[2\]
rlabel metal2 13048 44296 13048 44296 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[3\]
rlabel metal2 13720 44707 13720 44707 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[4\]
rlabel metal2 17864 45808 17864 45808 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[5\]
rlabel metal3 18032 45752 18032 45752 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[6\]
rlabel metal3 17024 43512 17024 43512 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[7\]
rlabel metal2 16184 42644 16184 42644 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[8\]
rlabel metal3 8456 41048 8456 41048 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[9\]
rlabel metal2 14280 35168 14280 35168 0 tt_um_rejunity_ay8913.tone_C_generator.period\[0\]
rlabel metal2 9912 34300 9912 34300 0 tt_um_rejunity_ay8913.tone_C_generator.period\[10\]
rlabel metal2 7896 36344 7896 36344 0 tt_um_rejunity_ay8913.tone_C_generator.period\[11\]
rlabel metal2 16968 36834 16968 36834 0 tt_um_rejunity_ay8913.tone_C_generator.period\[1\]
rlabel metal2 12936 37408 12936 37408 0 tt_um_rejunity_ay8913.tone_C_generator.period\[2\]
rlabel metal2 12264 35980 12264 35980 0 tt_um_rejunity_ay8913.tone_C_generator.period\[3\]
rlabel metal3 18872 40376 18872 40376 0 tt_um_rejunity_ay8913.tone_C_generator.period\[4\]
rlabel metal2 20664 44912 20664 44912 0 tt_um_rejunity_ay8913.tone_C_generator.period\[5\]
rlabel metal2 21112 44632 21112 44632 0 tt_um_rejunity_ay8913.tone_C_generator.period\[6\]
rlabel metal2 20664 42392 20664 42392 0 tt_um_rejunity_ay8913.tone_C_generator.period\[7\]
rlabel via2 10472 33306 10472 33306 0 tt_um_rejunity_ay8913.tone_C_generator.period\[8\]
rlabel metal2 10024 37520 10024 37520 0 tt_um_rejunity_ay8913.tone_C_generator.period\[9\]
rlabel metal2 31192 22792 31192 22792 0 tt_um_rejunity_ay8913.tone_disable_A
rlabel via2 26040 23142 26040 23142 0 tt_um_rejunity_ay8913.tone_disable_B
rlabel via2 26600 23898 26600 23898 0 tt_um_rejunity_ay8913.tone_disable_C
rlabel metal2 6104 31192 6104 31192 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 51000 51000
<< end >>
