VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_tholin_riscv
  CLASS BLOCK ;
  FOREIGN wrapped_tholin_riscv ;
  ORIGIN 0.000 0.000 ;
  SIZE 1150.000 BY 1150.000 ;
  PIN custom_settings[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 90.720 4.000 91.280 ;
    END
  END custom_settings[0]
  PIN custom_settings[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.960 4.000 121.520 ;
    END
  END custom_settings[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 151.200 4.000 151.760 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 453.600 4.000 454.160 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 483.840 4.000 484.400 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 514.080 4.000 514.640 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 544.320 4.000 544.880 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 574.560 4.000 575.120 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 604.800 4.000 605.360 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 635.040 4.000 635.600 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 665.280 4.000 665.840 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 695.520 4.000 696.080 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 725.760 4.000 726.320 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 181.440 4.000 182.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 756.000 4.000 756.560 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 786.240 4.000 786.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 816.480 4.000 817.040 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 846.720 4.000 847.280 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 876.960 4.000 877.520 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 907.200 4.000 907.760 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 937.440 4.000 938.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 967.680 4.000 968.240 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 997.920 4.000 998.480 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1028.160 4.000 1028.720 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 211.680 4.000 212.240 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1058.400 4.000 1058.960 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1088.640 4.000 1089.200 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1118.880 4.000 1119.440 ;
    END
  END io_in[32]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 241.920 4.000 242.480 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 272.160 4.000 272.720 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 302.400 4.000 302.960 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 332.640 4.000 333.200 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 362.880 4.000 363.440 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 393.120 4.000 393.680 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 423.360 4.000 423.920 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 19.040 1146.000 19.600 1150.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 1146.000 366.800 1150.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 400.960 1146.000 401.520 1150.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 435.680 1146.000 436.240 1150.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 470.400 1146.000 470.960 1150.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 505.120 1146.000 505.680 1150.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 539.840 1146.000 540.400 1150.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 574.560 1146.000 575.120 1150.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 609.280 1146.000 609.840 1150.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 644.000 1146.000 644.560 1150.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 1146.000 679.280 1150.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 1146.000 54.320 1150.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 713.440 1146.000 714.000 1150.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 748.160 1146.000 748.720 1150.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 782.880 1146.000 783.440 1150.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 817.600 1146.000 818.160 1150.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 852.320 1146.000 852.880 1150.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 887.040 1146.000 887.600 1150.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 921.760 1146.000 922.320 1150.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 956.480 1146.000 957.040 1150.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 991.200 1146.000 991.760 1150.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1025.920 1146.000 1026.480 1150.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 88.480 1146.000 89.040 1150.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1060.640 1146.000 1061.200 1150.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1095.360 1146.000 1095.920 1150.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1130.080 1146.000 1130.640 1150.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 123.200 1146.000 123.760 1150.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 1146.000 158.480 1150.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 192.640 1146.000 193.200 1150.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 227.360 1146.000 227.920 1150.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 1146.000 262.640 1150.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 296.800 1146.000 297.360 1150.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 331.520 1146.000 332.080 1150.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 19.040 0.000 19.600 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 0.000 366.800 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 400.960 0.000 401.520 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 435.680 0.000 436.240 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 470.400 0.000 470.960 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 505.120 0.000 505.680 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 539.840 0.000 540.400 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 574.560 0.000 575.120 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 609.280 0.000 609.840 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 644.000 0.000 644.560 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 0.000 679.280 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 0.000 54.320 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 713.440 0.000 714.000 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 748.160 0.000 748.720 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 782.880 0.000 783.440 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 817.600 0.000 818.160 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 852.320 0.000 852.880 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 887.040 0.000 887.600 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 921.760 0.000 922.320 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 956.480 0.000 957.040 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 991.200 0.000 991.760 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1025.920 0.000 1026.480 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 88.480 0.000 89.040 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1060.640 0.000 1061.200 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1095.360 0.000 1095.920 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1130.080 0.000 1130.640 4.000 ;
    END
  END io_out[32]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 123.200 0.000 123.760 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 0.000 158.480 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 192.640 0.000 193.200 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 227.360 0.000 227.920 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 0.000 262.640 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 296.800 0.000 297.360 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 331.520 0.000 332.080 4.000 ;
    END
  END io_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 60.480 4.000 61.040 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 1133.180 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 1133.180 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 30.240 4.000 30.800 ;
    END
  END wb_clk_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 1142.960 1134.410 ;
      LAYER Metal2 ;
        RECT 6.860 1145.700 18.740 1146.740 ;
        RECT 19.900 1145.700 53.460 1146.740 ;
        RECT 54.620 1145.700 88.180 1146.740 ;
        RECT 89.340 1145.700 122.900 1146.740 ;
        RECT 124.060 1145.700 157.620 1146.740 ;
        RECT 158.780 1145.700 192.340 1146.740 ;
        RECT 193.500 1145.700 227.060 1146.740 ;
        RECT 228.220 1145.700 261.780 1146.740 ;
        RECT 262.940 1145.700 296.500 1146.740 ;
        RECT 297.660 1145.700 331.220 1146.740 ;
        RECT 332.380 1145.700 365.940 1146.740 ;
        RECT 367.100 1145.700 400.660 1146.740 ;
        RECT 401.820 1145.700 435.380 1146.740 ;
        RECT 436.540 1145.700 470.100 1146.740 ;
        RECT 471.260 1145.700 504.820 1146.740 ;
        RECT 505.980 1145.700 539.540 1146.740 ;
        RECT 540.700 1145.700 574.260 1146.740 ;
        RECT 575.420 1145.700 608.980 1146.740 ;
        RECT 610.140 1145.700 643.700 1146.740 ;
        RECT 644.860 1145.700 678.420 1146.740 ;
        RECT 679.580 1145.700 713.140 1146.740 ;
        RECT 714.300 1145.700 747.860 1146.740 ;
        RECT 749.020 1145.700 782.580 1146.740 ;
        RECT 783.740 1145.700 817.300 1146.740 ;
        RECT 818.460 1145.700 852.020 1146.740 ;
        RECT 853.180 1145.700 886.740 1146.740 ;
        RECT 887.900 1145.700 921.460 1146.740 ;
        RECT 922.620 1145.700 956.180 1146.740 ;
        RECT 957.340 1145.700 990.900 1146.740 ;
        RECT 992.060 1145.700 1025.620 1146.740 ;
        RECT 1026.780 1145.700 1060.340 1146.740 ;
        RECT 1061.500 1145.700 1095.060 1146.740 ;
        RECT 1096.220 1145.700 1129.780 1146.740 ;
        RECT 1130.940 1145.700 1142.260 1146.740 ;
        RECT 6.860 4.300 1142.260 1145.700 ;
        RECT 6.860 3.500 18.740 4.300 ;
        RECT 19.900 3.500 53.460 4.300 ;
        RECT 54.620 3.500 88.180 4.300 ;
        RECT 89.340 3.500 122.900 4.300 ;
        RECT 124.060 3.500 157.620 4.300 ;
        RECT 158.780 3.500 192.340 4.300 ;
        RECT 193.500 3.500 227.060 4.300 ;
        RECT 228.220 3.500 261.780 4.300 ;
        RECT 262.940 3.500 296.500 4.300 ;
        RECT 297.660 3.500 331.220 4.300 ;
        RECT 332.380 3.500 365.940 4.300 ;
        RECT 367.100 3.500 400.660 4.300 ;
        RECT 401.820 3.500 435.380 4.300 ;
        RECT 436.540 3.500 470.100 4.300 ;
        RECT 471.260 3.500 504.820 4.300 ;
        RECT 505.980 3.500 539.540 4.300 ;
        RECT 540.700 3.500 574.260 4.300 ;
        RECT 575.420 3.500 608.980 4.300 ;
        RECT 610.140 3.500 643.700 4.300 ;
        RECT 644.860 3.500 678.420 4.300 ;
        RECT 679.580 3.500 713.140 4.300 ;
        RECT 714.300 3.500 747.860 4.300 ;
        RECT 749.020 3.500 782.580 4.300 ;
        RECT 783.740 3.500 817.300 4.300 ;
        RECT 818.460 3.500 852.020 4.300 ;
        RECT 853.180 3.500 886.740 4.300 ;
        RECT 887.900 3.500 921.460 4.300 ;
        RECT 922.620 3.500 956.180 4.300 ;
        RECT 957.340 3.500 990.900 4.300 ;
        RECT 992.060 3.500 1025.620 4.300 ;
        RECT 1026.780 3.500 1060.340 4.300 ;
        RECT 1061.500 3.500 1095.060 4.300 ;
        RECT 1096.220 3.500 1129.780 4.300 ;
        RECT 1130.940 3.500 1142.260 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 1119.740 1142.310 1138.340 ;
        RECT 4.300 1118.580 1142.310 1119.740 ;
        RECT 4.000 1089.500 1142.310 1118.580 ;
        RECT 4.300 1088.340 1142.310 1089.500 ;
        RECT 4.000 1059.260 1142.310 1088.340 ;
        RECT 4.300 1058.100 1142.310 1059.260 ;
        RECT 4.000 1029.020 1142.310 1058.100 ;
        RECT 4.300 1027.860 1142.310 1029.020 ;
        RECT 4.000 998.780 1142.310 1027.860 ;
        RECT 4.300 997.620 1142.310 998.780 ;
        RECT 4.000 968.540 1142.310 997.620 ;
        RECT 4.300 967.380 1142.310 968.540 ;
        RECT 4.000 938.300 1142.310 967.380 ;
        RECT 4.300 937.140 1142.310 938.300 ;
        RECT 4.000 908.060 1142.310 937.140 ;
        RECT 4.300 906.900 1142.310 908.060 ;
        RECT 4.000 877.820 1142.310 906.900 ;
        RECT 4.300 876.660 1142.310 877.820 ;
        RECT 4.000 847.580 1142.310 876.660 ;
        RECT 4.300 846.420 1142.310 847.580 ;
        RECT 4.000 817.340 1142.310 846.420 ;
        RECT 4.300 816.180 1142.310 817.340 ;
        RECT 4.000 787.100 1142.310 816.180 ;
        RECT 4.300 785.940 1142.310 787.100 ;
        RECT 4.000 756.860 1142.310 785.940 ;
        RECT 4.300 755.700 1142.310 756.860 ;
        RECT 4.000 726.620 1142.310 755.700 ;
        RECT 4.300 725.460 1142.310 726.620 ;
        RECT 4.000 696.380 1142.310 725.460 ;
        RECT 4.300 695.220 1142.310 696.380 ;
        RECT 4.000 666.140 1142.310 695.220 ;
        RECT 4.300 664.980 1142.310 666.140 ;
        RECT 4.000 635.900 1142.310 664.980 ;
        RECT 4.300 634.740 1142.310 635.900 ;
        RECT 4.000 605.660 1142.310 634.740 ;
        RECT 4.300 604.500 1142.310 605.660 ;
        RECT 4.000 575.420 1142.310 604.500 ;
        RECT 4.300 574.260 1142.310 575.420 ;
        RECT 4.000 545.180 1142.310 574.260 ;
        RECT 4.300 544.020 1142.310 545.180 ;
        RECT 4.000 514.940 1142.310 544.020 ;
        RECT 4.300 513.780 1142.310 514.940 ;
        RECT 4.000 484.700 1142.310 513.780 ;
        RECT 4.300 483.540 1142.310 484.700 ;
        RECT 4.000 454.460 1142.310 483.540 ;
        RECT 4.300 453.300 1142.310 454.460 ;
        RECT 4.000 424.220 1142.310 453.300 ;
        RECT 4.300 423.060 1142.310 424.220 ;
        RECT 4.000 393.980 1142.310 423.060 ;
        RECT 4.300 392.820 1142.310 393.980 ;
        RECT 4.000 363.740 1142.310 392.820 ;
        RECT 4.300 362.580 1142.310 363.740 ;
        RECT 4.000 333.500 1142.310 362.580 ;
        RECT 4.300 332.340 1142.310 333.500 ;
        RECT 4.000 303.260 1142.310 332.340 ;
        RECT 4.300 302.100 1142.310 303.260 ;
        RECT 4.000 273.020 1142.310 302.100 ;
        RECT 4.300 271.860 1142.310 273.020 ;
        RECT 4.000 242.780 1142.310 271.860 ;
        RECT 4.300 241.620 1142.310 242.780 ;
        RECT 4.000 212.540 1142.310 241.620 ;
        RECT 4.300 211.380 1142.310 212.540 ;
        RECT 4.000 182.300 1142.310 211.380 ;
        RECT 4.300 181.140 1142.310 182.300 ;
        RECT 4.000 152.060 1142.310 181.140 ;
        RECT 4.300 150.900 1142.310 152.060 ;
        RECT 4.000 121.820 1142.310 150.900 ;
        RECT 4.300 120.660 1142.310 121.820 ;
        RECT 4.000 91.580 1142.310 120.660 ;
        RECT 4.300 90.420 1142.310 91.580 ;
        RECT 4.000 61.340 1142.310 90.420 ;
        RECT 4.300 60.180 1142.310 61.340 ;
        RECT 4.000 31.100 1142.310 60.180 ;
        RECT 4.300 29.940 1142.310 31.100 ;
        RECT 4.000 6.860 1142.310 29.940 ;
      LAYER Metal4 ;
        RECT 9.660 1133.480 1133.300 1137.270 ;
        RECT 9.660 15.080 21.940 1133.480 ;
        RECT 24.140 15.080 98.740 1133.480 ;
        RECT 100.940 15.080 175.540 1133.480 ;
        RECT 177.740 15.080 252.340 1133.480 ;
        RECT 254.540 15.080 329.140 1133.480 ;
        RECT 331.340 15.080 405.940 1133.480 ;
        RECT 408.140 15.080 482.740 1133.480 ;
        RECT 484.940 15.080 559.540 1133.480 ;
        RECT 561.740 15.080 636.340 1133.480 ;
        RECT 638.540 15.080 713.140 1133.480 ;
        RECT 715.340 15.080 789.940 1133.480 ;
        RECT 792.140 15.080 866.740 1133.480 ;
        RECT 868.940 15.080 943.540 1133.480 ;
        RECT 945.740 15.080 1020.340 1133.480 ;
        RECT 1022.540 15.080 1097.140 1133.480 ;
        RECT 1099.340 15.080 1133.300 1133.480 ;
        RECT 9.660 6.810 1133.300 15.080 ;
  END
END wrapped_tholin_riscv
END LIBRARY

