* NGSPICE file created from tholin_avalonsemi_tbb1143.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 D RN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 D SETN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_1 D CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

.subckt tholin_avalonsemi_tbb1143 clk io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] rst_n vdd vss
XFILLER_0_49_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1270_ CIRCUIT_2223.tone_generator_2_2.MEMORY_32.d _0048_ CIRCUIT_2223.MEMORY_18.s_currentState
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_32.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_0985_ _0165_ CIRCUIT_2223.tone_generator_2_2.GATES_8.input2 _0446_ _0447_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_9_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0770_ _0164_ _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1253_ CIRCUIT_2223.tone_generator_2_1.MEMORY_28.clock _0043_ CIRCUIT_2223.tone_generator_2_1.MEMORY_37.s_currentState
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_38.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_1184_ CIRCUIT_2223.tone_generator_1.MEMORY_11.s_currentState _0002_ net19 CIRCUIT_2223.tone_generator_1.MEMORY_12.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XTAP_TAPCELL_ROW_34_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0968_ _0434_ _0436_ _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_19_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0899_ _0193_ _0387_ _0390_ _0104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_25_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0822_ CIRCUIT_2223.GATES_3.input2 CIRCUIT_2223.GATES_2.input2 CIRCUIT_2223.tone_generator_2_2.MEMORY_39.s_currentState
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_39.s_currentState _0338_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and4_1
X_0753_ spi_dac_i_2.spi_dat_buff\[4\] _0073_ _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0684_ CIRCUIT_2223.tone_generator_2_1.MEMORY_36.s_currentState CIRCUIT_2223.tone_generator_2_1.GATES_15.input2
+ _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_39_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1236_ _0115_ net26 CIRCUIT_2223.triangle_wave_generator_1.GATES_12.input2 vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1167_ _0093_ net59 slow_clock\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1098_ _0373_ _0172_ _0462_ _0516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_19_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_8_Left_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0780__A1 _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1021_ _0469_ _0035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0805_ _0319_ _0322_ _0323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0736_ _0267_ spi_dac_i_2.counter\[1\] _0271_ _0069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0598_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.s_currentState CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0667_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_38.s_currentState _0205_ _0206_
+ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.s_currentState _0207_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1219_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.d _0024_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.s_currentState
+ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.s_currentState vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1004_ _0456_ _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0719_ CIRCUIT_2223.tone_generator_2_2.GATES_11.input2 _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_37_Left_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0984_ _0154_ _0445_ _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1124__A1 net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1221__CLK net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1252_ CIRCUIT_2223.tone_generator_2_1.MEMORY_37.d _0042_ CIRCUIT_2223.tone_generator_2_1.MEMORY_36.s_currentState
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_37.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_1183_ CIRCUIT_2223.tone_generator_1.MEMORY_10.s_currentState net19 CIRCUIT_2223.tone_generator_1.MEMORY_11.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0967_ _0428_ _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0898_ _0389_ _0386_ _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_25_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_48_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0752_ spi_dac_i_2.spi_dat_buff\[3\] _0068_ _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0821_ _0337_ _0088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0683_ CIRCUIT_2223.tone_generator_2_1.MEMORY_37.s_currentState _0220_ CIRCUIT_2223.tone_generator_2_1.GATES_8.input2
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_29.d _0221_ _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_19_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_24_Left_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1166_ _0092_ net51 slow_clock\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1235_ _0114_ net26 CIRCUIT_2223.triangle_wave_generator_1.GATES_11.input2 vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1097_ _0515_ _0054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_30_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1020_ _0422_ _0466_ _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_44_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0804_ _0320_ CIRCUIT_2223.GATES_4.input1\[2\] CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState
+ _0321_ _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_0735_ _0267_ spi_dac_i_2.counter\[1\] _0269_ _0270_ _0271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_21_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0597_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.s_currentState CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0666_ CIRCUIT_2223.triangle_wave_generator_1.GATES_9.input2 _0206_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1149_ _0075_ net57 spi_dac_i_2.spi_dat_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1218_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.d _0023_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.s_currentState
+ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.s_currentState vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_0_30_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1002__I0 _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0577__I CIRCUIT_2223.MEMORY_18.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1003_ _0457_ _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0718_ CIRCUIT_2223.tone_generator_2_2.MEMORY_35.s_currentState _0248_ _0252_ CIRCUIT_2223.tone_generator_2_2.MEMORY_30.s_currentState
+ _0256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_0649_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_15.input2 _0190_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_11_Left_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput10 net10 io_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input3_I io_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_17_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_8_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0983_ _0151_ _0424_ _0445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_1_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout61_I net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1182_ CIRCUIT_2223.tone_generator_1.GATES_3.result net19 CIRCUIT_2223.tone_generator_1.MEMORY_10.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1251_ CIRCUIT_2223.tone_generator_2_1.MEMORY_36.d _0041_ CIRCUIT_2223.tone_generator_2_1.MEMORY_35.s_currentState
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_36.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_0_27_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0897_ _0161_ _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0966_ _0435_ _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0751_ _0279_ _0280_ _0075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0820_ _0293_ _0336_ _0337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_36_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1303_ CIRCUIT_2223.MEMORY_18.d _0067_ CIRCUIT_2223.MEMORY_26.s_currentState CIRCUIT_2223.MEMORY_18.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_0682_ CIRCUIT_2223.tone_generator_2_1.MEMORY_33.d CIRCUIT_2223.tone_generator_2_1.GATES_12.input2
+ _0220_ CIRCUIT_2223.tone_generator_2_1.MEMORY_37.s_currentState _0221_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1165_ _0091_ net51 slow_clock\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1096_ _0367_ _0500_ _0515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1234_ _0113_ net45 CIRCUIT_2223.tone_generator_2_2.GATES_10.input2 vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout24_I net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0949_ _0423_ _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_41_Left_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1024__I _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0863__I _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0803_ CIRCUIT_2223.GATES_5.input2 _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0734_ _0263_ _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0665_ CIRCUIT_2223.triangle_wave_generator_1.GATES_17.input2 _0205_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0596_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.s_currentState CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1148_ _0074_ net56 spi_dac_i_2.spi_dat_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1079_ _0505_ _0046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1217_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.d _0022_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_38.s_currentState
+ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.s_currentState vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XTAP_TAPCELL_ROW_41_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1002_ _0165_ CIRCUIT_2223.triangle_wave_generator_1.GATES_15.input2 _0456_ _0457_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_29_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0648_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.d CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_11.input2
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_12.input2 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.d
+ _0189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0717_ CIRCUIT_2223.tone_generator_2_2.MEMORY_28.clock CIRCUIT_2223.tone_generator_2_2.GATES_17.input2
+ _0251_ CIRCUIT_2223.tone_generator_2_2.MEMORY_28.s_currentState _0255_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0579_ _0174_ CIRCUIT_2223.GATES_11.result vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput11 net11 io_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput9 net9 io_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_17_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0982_ _0444_ _0032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_38_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1181_ CIRCUIT_2223.tone_generator_1.MEMORY_8.s_currentState net17 CIRCUIT_2223.tone_generator_1.MEMORY_9.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1250_ CIRCUIT_2223.tone_generator_2_1.MEMORY_35.d _0040_ CIRCUIT_2223.tone_generator_2_1.MEMORY_34.s_currentState
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_35.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XTAP_TAPCELL_ROW_19_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0896_ _0196_ _0387_ _0388_ _0103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0965_ _0434_ _0430_ _0435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0750_ spi_dac_i_2.spi_dat_buff\[3\] _0073_ _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0681_ CIRCUIT_2223.tone_generator_2_1.GATES_16.input2 _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_24_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1302_ CIRCUIT_2223.MEMORY_19.d _0066_ CIRCUIT_2223.MEMORY_18.s_currentState CIRCUIT_2223.MEMORY_19.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_1233_ _0112_ net45 CIRCUIT_2223.tone_generator_2_2.GATES_9.input2 vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1164_ _0090_ net50 spi_dac_i_2.spi_dat_buff\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1095_ _0514_ _0053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1163__CLK net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0948_ _0422_ _0407_ _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_22_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0879_ net4 _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_33_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0802_ CIRCUIT_2223.s_logisimNet48 _0320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0733_ _0268_ _0269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0664_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.d CIRCUIT_2223.triangle_wave_generator_1.GATES_15.input2
+ _0203_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.s_currentState _0204_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_0595_ net14 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.clock vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1216_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.d _0021_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_38.s_currentState
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.s_currentState vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1147_ _0073_ net58 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1078_ _0504_ _0501_ _0505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_47_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0995__A1 _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0964__I _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0910__A1 _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1001_ _0297_ _0403_ _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_32_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0578_ CIRCUIT_2223.GATES_11.input2 net53 _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_0647_ _0182_ _0185_ _0186_ _0187_ _0188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_12_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0716_ _0246_ _0247_ _0250_ _0253_ _0254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput12 net12 io_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_27_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1247__CLK CIRCUIT_2223.MEMORY_18.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0981_ _0440_ _0429_ _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout47_I net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1180_ CIRCUIT_2223.tone_generator_1.GATES_2.result net17 CIRCUIT_2223.tone_generator_1.MEMORY_8.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_19_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0964_ _0367_ _0434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0895_ _0376_ _0387_ _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_33_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0680_ _0219_ CIRCUIT_2223.triangle_wave_generator_1.GATES_27.result vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1301_ CIRCUIT_2223.MEMORY_20.d _0065_ CIRCUIT_2223.MEMORY_19.s_currentState CIRCUIT_2223.MEMORY_20.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_0_19_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1232_ _0111_ net44 CIRCUIT_2223.tone_generator_2_2.GATES_8.input2 vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_47_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1163_ _0089_ net53 spi_dac_i_2.spi_dat_buff\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1094_ _0510_ _0500_ _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_0947_ _0401_ _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0878_ _0374_ _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_33_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Left_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0801_ CIRCUIT_2223.s_logisimNet48 CIRCUIT_2223.GATES_5.input2 CIRCUIT_2223.GATES_4.input1\[2\]
+ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState _0319_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_21_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0594_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.clock
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0732_ _0264_ _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0663_ CIRCUIT_2223.triangle_wave_generator_1.GATES_16.input2 _0203_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1146_ _0072_ net55 spi_dac_i_2.counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1215_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.d _0020_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.s_currentState
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_0_47_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1077_ _0471_ _0504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_30_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1000_ _0455_ _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0715_ CIRCUIT_2223.tone_generator_2_2.MEMORY_28.s_currentState _0251_ _0252_ CIRCUIT_2223.tone_generator_2_2.MEMORY_30.s_currentState
+ _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_0577_ CIRCUIT_2223.MEMORY_18.s_currentState CIRCUIT_2223.MEMORY_18.d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0646_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.d CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_13.input2
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_16.input2 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.d
+ _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1129_ _0533_ _0534_ _0056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput13 net13 io_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_43_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0895__A1 _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_15_Left_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0629_ CIRCUIT_2223.tone_generator_2_2.MEMORY_37.s_currentState CIRCUIT_2223.tone_generator_2_2.MEMORY_37.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1063__A1 _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_14_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0980_ _0443_ _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input1_I clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1045__A1 _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0894_ _0386_ _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0963_ _0433_ _0024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_33_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1231_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.clock CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState
+ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_42.s_currentState vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_1162_ _0088_ net54 spi_dac_i_2.spi_dat_buff\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1300_ CIRCUIT_2223.MEMORY_21.d _0064_ CIRCUIT_2223.MEMORY_20.s_currentState CIRCUIT_2223.MEMORY_21.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XTAP_TAPCELL_ROW_47_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1093_ _0513_ _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1099__I1 _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0946_ _0421_ _0020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0877_ _0373_ _0168_ _0297_ _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_15_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_3_Left_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0731_ spi_dac_i_2.counter\[0\] _0267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0800_ _0294_ _0316_ _0318_ _0086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_21_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0593_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.s_currentState CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0662_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.d CIRCUIT_2223.triangle_wave_generator_1.GATES_13.input2
+ CIRCUIT_2223.triangle_wave_generator_1.GATES_10.input2 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.d
+ _0201_ _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_1145_ _0071_ net54 spi_dac_i_2.counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1214_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.d _0019_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.s_currentState vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_0_1_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1076_ _0503_ _0045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0929_ _0411_ _0408_ _0412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__0999__S _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_45_Left_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_41_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0645_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.d CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_14.input2
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_9.input2 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.d
+ _0186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0714_ CIRCUIT_2223.tone_generator_2_2.GATES_9.input2 _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__0985__I0 _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0576_ CIRCUIT_2223.MEMORY_19.s_currentState CIRCUIT_2223.MEMORY_19.d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1128_ _0533_ _0534_ _0055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1059_ _0168_ _0170_ _0462_ _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_35_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1270__CLK CIRCUIT_2223.MEMORY_18.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0628_ CIRCUIT_2223.tone_generator_2_2.MEMORY_36.s_currentState CIRCUIT_2223.tone_generator_2_2.MEMORY_36.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0559_ _0166_ _0144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_32_Left_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1117__I0 _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1289__D net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_19_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0962_ _0002_ _0430_ _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_0893_ _0373_ _0385_ _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_10_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout52_I net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_33_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0777__A1 _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout60 net61 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_47_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1230_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.clock net14 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_1161_ _0087_ net50 spi_dac_i_2.spi_dat_buff\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1092_ _0510_ _0500_ _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_19_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0945_ _0417_ _0407_ _0421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_0876_ _0169_ _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0730_ _0266_ _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0661_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.clock CIRCUIT_2223.triangle_wave_generator_1.GATES_17.input2
+ CIRCUIT_2223.triangle_wave_generator_1.GATES_7.input2 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.d
+ _0201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_24_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0592_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1213_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.d _0018_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.s_currentState
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.s_currentState vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_1144_ _0070_ net54 spi_dac_i_2.counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1075_ _0478_ _0501_ _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_7_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0859_ _0291_ _0365_ _0098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0928_ _0401_ _0411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_38_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0644_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_38.s_currentState
+ _0183_ _0184_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.s_currentState
+ _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0713_ CIRCUIT_2223.tone_generator_2_2.GATES_7.input2 _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0575_ CIRCUIT_2223.MEMORY_20.s_currentState CIRCUIT_2223.MEMORY_20.d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1127_ _0363_ _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1058_ _0227_ _0487_ _0491_ _0128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0900__I1 _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0558_ _0165_ CIRCUIT_2223.GATES_2.input2 _0155_ _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_0627_ CIRCUIT_2223.tone_generator_2_2.MEMORY_35.s_currentState CIRCUIT_2223.tone_generator_2_2.MEMORY_35.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1053__I0 _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0961_ _0432_ _0023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0892_ _0167_ _0296_ _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_2_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout50 net61 net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout61 net1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_47_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1160_ _0086_ net50 spi_dac_i_2.spi_dat_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1091_ _0512_ _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0944_ _0420_ _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0875_ _0371_ _0372_ _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1289_ net4 _0001_ net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_21_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0591_ net15 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.d vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_21_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0660_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.s_currentState CIRCUIT_2223.triangle_wave_generator_1.GATES_8.input2
+ _0200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1212_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.d _0017_ net25
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_1143_ _0069_ net54 spi_dac_i_2.counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1074_ _0502_ _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0927_ _0410_ _0012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0789_ CIRCUIT_2223.s_logisimNet48 CIRCUIT_2223.GATES_5.input2 CIRCUIT_2223.GATES_4.input1\[0\]
+ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState _0309_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_0858_ _0363_ _0364_ _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0574_ CIRCUIT_2223.MEMORY_21.s_currentState CIRCUIT_2223.MEMORY_21.d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0643_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_9.input2 _0184_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__0898__A1 _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0712_ CIRCUIT_2223.tone_generator_2_2.MEMORY_35.s_currentState _0248_ _0249_ CIRCUIT_2223.tone_generator_2_2.MEMORY_31.s_currentState
+ _0250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1126_ _0354_ _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1057_ _0383_ _0486_ _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1057__A1 _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0557_ _0164_ _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0626_ CIRCUIT_2223.tone_generator_2_2.MEMORY_34.s_currentState CIRCUIT_2223.tone_generator_2_2.MEMORY_34.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1109_ _0257_ _0522_ _0523_ _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_19_Left_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0609_ CIRCUIT_2223.tone_generator_2_1.MEMORY_29.s_currentState CIRCUIT_2223.tone_generator_2_1.MEMORY_29.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_36_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0960_ _0002_ _0430_ _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_6_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0891_ _0191_ _0375_ _0384_ _0102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_2_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout51 net52 net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout40 net41 net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1090_ _0510_ _0507_ _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_0874_ _0371_ _0372_ _0009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_30_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0943_ _0417_ _0407_ _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_2_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1288_ _0143_ net46 CIRCUIT_2223.tone_generator_2_2.GATES_7.input2 vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0590_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.s_currentState
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1142_ _0068_ net58 spi_dac_i_2.counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1211_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.d _0016_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.s_currentState vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_0_47_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1073_ _0402_ _0501_ _0502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_0857_ slow_clock\[6\] _0360_ _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0926_ _0402_ _0408_ _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_15_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0788_ _0308_ _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_7_Left_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0711_ CIRCUIT_2223.tone_generator_2_2.GATES_10.input2 _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0573_ CIRCUIT_2223.MEMORY_22.s_currentState CIRCUIT_2223.MEMORY_22.d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0642_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_17.input2 _0183_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1125_ _0251_ _0529_ _0532_ _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_49_Left_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1056_ _0224_ _0487_ _0490_ _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0909_ _0394_ _0397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_27_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0625_ CIRCUIT_2223.tone_generator_2_2.MEMORY_33.s_currentState CIRCUIT_2223.tone_generator_2_2.MEMORY_33.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0556_ net4 _0164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1039_ _0480_ _0042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1108_ _0164_ _0522_ _0523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_31_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0608_ CIRCUIT_2223.tone_generator_2_1.MEMORY_28.s_currentState CIRCUIT_2223.tone_generator_2_1.MEMORY_28.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0539_ CIRCUIT_2223.GATES_1.input1\[2\] _0150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_36_Left_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0890_ _0383_ _0377_ _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_35_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1120__A1 _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout52 net53 net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout30 net31 net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout41 net48 net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1102__A1 _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0873_ _0371_ _0372_ _0008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_30_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0942_ _0419_ _0018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1287_ _0142_ net44 CIRCUIT_2223.tone_generator_2_2.GATES_17.input2 vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0997__I1 _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1141_ _0536_ _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1210_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.d _0015_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.s_currentState
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.s_currentState vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_1072_ _0500_ _0501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_23_Left_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0787_ spi_dac_i_2.spi_dat_buff\[0\] _0288_ _0306_ spi_dac_i_2.spi_dat_buff\[1\]
+ _0307_ _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_0856_ net46 _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0925_ _0409_ _0011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0641_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.d CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_15.input2
+ _0181_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.s_currentState
+ _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0710_ CIRCUIT_2223.tone_generator_2_2.GATES_14.input2 _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0572_ CIRCUIT_2223.MEMORY_23.s_currentState CIRCUIT_2223.GATES_11.input2 vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1055_ _0157_ _0486_ _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1124_ net7 _0529_ _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0839_ _0293_ _0350_ _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0908_ _0167_ _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0537__I net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0624_ CIRCUIT_2223.tone_generator_2_2.MEMORY_32.s_currentState CIRCUIT_2223.tone_generator_2_2.MEMORY_32.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0555_ _0163_ _0145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1038_ _0478_ _0465_ _0480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1107_ _0521_ _0522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_16_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_10_Left_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1047__I0 _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0538_ CIRCUIT_2223.s_logisimNet48 _0149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0607_ CIRCUIT_2223.tone_generator_2_1.MEMORY_39.s_currentState CIRCUIT_2223.tone_generator_2_1.MEMORY_39.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout20 net22 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout53 net61 net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout42 net43 net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout31 net35 net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0941_ _0417_ _0414_ _0419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_0872_ _0371_ _0372_ _0007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_30_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1286_ _0141_ net46 CIRCUIT_2223.tone_generator_2_2.GATES_16.input2 vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_21_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1096__A1 _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1140_ _0536_ _0066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1071_ _0499_ _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0924_ _0402_ _0408_ _0409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_0786_ _0292_ _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0855_ slow_clock\[6\] _0360_ _0362_ _0097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1269_ CIRCUIT_2223.tone_generator_2_2.MEMORY_31.d _0047_ CIRCUIT_2223.tone_generator_2_2.MEMORY_30.s_currentState
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_31.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XPHY_EDGE_ROW_40_Left_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0640_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_16.input2 _0181_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0571_ net24 CIRCUIT_2223.MEMORY_24.d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1054_ _0489_ _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1123_ _0531_ _0142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0907_ _0395_ _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0838_ _0347_ slow_clock\[1\] slow_clock\[2\] _0350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_0769_ _0293_ _0294_ _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1065__I1 _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0553__I _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0554_ _0162_ CIRCUIT_2223.GATES_3.input2 _0155_ _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_0623_ CIRCUIT_2223.tone_generator_2_2.MEMORY_31.s_currentState CIRCUIT_2223.tone_generator_2_2.MEMORY_31.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1106_ _0171_ _0445_ _0521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_48_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1037_ _0479_ _0041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0558__I0 _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0537_ net7 _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0606_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_38.s_currentState CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.clock
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_36_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout21 net22 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0916__I _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout54 net60 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout43 net44 net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout32 net33 net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0940_ _0418_ _0017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1110__I0 _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0871_ _0369_ _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_30_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1285_ _0140_ net42 CIRCUIT_2223.tone_generator_2_2.GATES_15.input2 vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0540__A1 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0906__I0 _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0556__I net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1070_ _0174_ CIRCUIT_2223.tone_generator_2_2.GATES_27.result _0445_ _0498_ _0499_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_0854_ slow_clock\[6\] _0360_ _0307_ _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0923_ _0407_ _0408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0785_ _0305_ _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1268_ CIRCUIT_2223.tone_generator_2_2.MEMORY_30.d _0046_ CIRCUIT_2223.tone_generator_2_2.MEMORY_29.s_currentState
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_30.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_0_36_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1199_ _0105_ net27 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_13.input2
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_40_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0570_ CIRCUIT_2223.MEMORY_25.s_currentState CIRCUIT_2223.MEMORY_25.d vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1122_ _0158_ CIRCUIT_2223.tone_generator_2_2.GATES_17.input2 _0527_ _0531_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1053_ _0162_ CIRCUIT_2223.tone_generator_2_1.GATES_12.input2 _0486_ _0489_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_0837_ _0347_ slow_clock\[1\] slow_clock\[2\] _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0906_ _0165_ _0373_ _0394_ _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_22_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0768_ _0286_ _0294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0699_ CIRCUIT_2223.tone_generator_2_1.MEMORY_32.d CIRCUIT_2223.tone_generator_2_1.GATES_11.input2
+ _0228_ CIRCUIT_2223.tone_generator_2_1.MEMORY_31.s_currentState _0238_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_11_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input8_I rst_n vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0553_ _0161_ _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0622_ CIRCUIT_2223.tone_generator_2_2.MEMORY_30.s_currentState CIRCUIT_2223.tone_generator_2_2.MEMORY_30.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1105_ _0228_ _0518_ _0520_ _0135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1036_ _0478_ _0465_ _0479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_16_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0605_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.s_currentState CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1019_ _0468_ _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1114__A1 net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout22 net23 net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout55 net60 net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout44 net47 net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout33 net34 net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0870_ _0354_ _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1284_ _0139_ net39 CIRCUIT_2223.tone_generator_2_2.GATES_14.input2 vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0999_ CIRCUIT_2223.triangle_wave_generator_1.GATES_14.input2 _0148_ _0426_ _0455_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__0540__A2 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0853_ _0360_ _0361_ _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0922_ _0406_ _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0784_ _0262_ _0268_ _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1198_ _0104_ net28 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_12.input2
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput1 clk net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1267_ CIRCUIT_2223.tone_generator_2_2.MEMORY_29.d _0045_ CIRCUIT_2223.tone_generator_2_2.MEMORY_28.s_currentState
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_29.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XPHY_EDGE_ROW_27_Left_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1052_ _0236_ _0487_ _0488_ _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1121_ _0241_ _0529_ _0530_ _0141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0767_ _0292_ _0293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0836_ _0291_ _0348_ _0092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0905_ net3 _0393_ _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0698_ CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState _0236_ CIRCUIT_2223.tone_generator_2_1.GATES_12.input2
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_33.d _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0621_ CIRCUIT_2223.tone_generator_2_2.MEMORY_29.s_currentState CIRCUIT_2223.tone_generator_2_2.MEMORY_29.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0552_ net5 _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1104_ _0302_ _0518_ _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1035_ _0471_ _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0819_ _0329_ _0287_ _0334_ _0269_ _0335_ _0336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_39_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0604_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.s_currentState CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_36_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1018_ _0422_ _0466_ _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_14_Left_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1172__CLK net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout56 net59 net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout23 net24 net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout45 net47 net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout34 net35 net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1283_ _0138_ net45 CIRCUIT_2223.tone_generator_2_2.GATES_13.input2 vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0998_ _0454_ _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1005__A1 _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0921_ _0174_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_27.result _0405_
+ net30 _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_0783_ _0304_ _0083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0852_ slow_clock\[5\] _0358_ _0307_ _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput2 io_in[0] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1197_ _0103_ net28 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_11.input2
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1266_ CIRCUIT_2223.tone_generator_2_2.MEMORY_28.d _0044_ CIRCUIT_2223.tone_generator_2_2.MEMORY_38.s_currentState
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_28.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XANTENNA_fanout41_I net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0763__I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_2_Left_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1051_ _0164_ _0487_ _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1120_ _0161_ _0529_ _0530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0904_ net2 _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0835_ _0347_ slow_clock\[1\] _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_43_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0766_ _0263_ _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0697_ CIRCUIT_2223.tone_generator_2_1.GATES_11.input2 _0236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1249_ CIRCUIT_2223.tone_generator_2_1.MEMORY_34.d _0039_ CIRCUIT_2223.tone_generator_2_1.MEMORY_33.s_currentState
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_34.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XPHY_EDGE_ROW_44_Left_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0551_ _0160_ _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0620_ CIRCUIT_2223.tone_generator_2_2.MEMORY_28.s_currentState CIRCUIT_2223.tone_generator_2_2.MEMORY_28.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1103_ _0231_ _0518_ _0519_ _0134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1034_ _0477_ _0040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0749_ spi_dac_i_2.spi_dat_buff\[2\] _0068_ _0279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0818_ spi_dac_i_2.spi_dat_buff\[9\] _0267_ _0268_ _0335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_3_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0861__I _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0603_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.s_currentState CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1017_ _0467_ _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1122__I0 _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_31_Left_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout57 net58 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout46 net47 net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_32_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout24 net25 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_24_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout35 net49 net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1282_ _0137_ net45 CIRCUIT_2223.tone_generator_2_2.GATES_12.input2 vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0997_ CIRCUIT_2223.triangle_wave_generator_1.GATES_13.input2 _0302_ _0426_ _0454_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_20_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_43_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0920_ _0385_ _0404_ _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0851_ slow_clock\[5\] _0358_ _0360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_0782_ spi_dac_i_2.spi_dat_buff\[0\] _0286_ _0288_ _0293_ _0304_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_11_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1265_ _0132_ net38 CIRCUIT_2223.tone_generator_2_1.GATES_7.input2 vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1196_ _0102_ net36 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_7.input2
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput3 io_in[1] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1050_ _0486_ _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0834_ _0291_ _0347_ _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0903_ _0194_ _0387_ _0392_ _0106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_22_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0765_ _0285_ _0288_ _0289_ _0291_ _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_0696_ CIRCUIT_2223.tone_generator_2_1.MEMORY_35.s_currentState _0227_ _0231_ CIRCUIT_2223.tone_generator_2_1.MEMORY_30.s_currentState
+ _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_11_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1248_ CIRCUIT_2223.tone_generator_2_1.MEMORY_33.d _0038_ CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_33.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_1179_ CIRCUIT_2223.tone_generator_1.GATES_1.result net17 CIRCUIT_2223.tone_generator_1.MEMORY_7.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0550_ _0158_ _0159_ _0155_ _0160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1102_ _0389_ _0518_ _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1033_ _0472_ _0473_ _0477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_0817_ _0332_ _0333_ _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0748_ _0277_ _0278_ _0074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0679_ _0200_ _0202_ _0210_ _0218_ _0219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0602_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.s_currentState CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input6_I io_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1016_ _0402_ _0466_ _0467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_8_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout14 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_42.s_currentState net14 vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout58 net59 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout47 net48 net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout36 net41 net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_24_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout25 CIRCUIT_2223.MEMORY_24.s_currentState net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1281_ _0136_ net39 CIRCUIT_2223.tone_generator_2_2.GATES_11.input2 vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0996_ _0212_ _0451_ _0453_ _0115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0850_ _0358_ _0359_ _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_43_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0781_ _0216_ _0300_ _0303_ _0082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_23_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1264_ _0131_ net37 CIRCUIT_2223.tone_generator_2_1.GATES_17.input2 vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput4 io_in[2] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1195_ _0101_ net36 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_17.input2
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0979_ _0440_ _0429_ _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0833_ slow_clock\[0\] _0347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0902_ _0383_ _0386_ _0392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0764_ _0290_ _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0695_ CIRCUIT_2223.tone_generator_2_1.MEMORY_28.clock CIRCUIT_2223.tone_generator_2_1.GATES_17.input2
+ _0230_ CIRCUIT_2223.tone_generator_2_1.MEMORY_28.s_currentState _0234_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1178_ CIRCUIT_2223.tone_generator_1.MEMORY_4.s_currentState net17 CIRCUIT_2223.tone_generator_1.MEMORY_6.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1247_ CIRCUIT_2223.tone_generator_2_1.MEMORY_32.d _0037_ CIRCUIT_2223.MEMORY_18.s_currentState
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_19_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1126__I _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1101_ _0516_ _0518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1032_ _0476_ _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0747_ spi_dac_i_2.spi_dat_buff\[2\] _0073_ _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0816_ _0323_ _0326_ _0319_ _0333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0678_ _0213_ _0214_ _0215_ _0217_ _0218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_30_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_7_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0601_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1015_ _0465_ _0466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_29_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_18_Left_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout15 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState
+ net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout37 net40 net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout26 net31 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_24_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout59 net60 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout48 net49 net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1280_ _0135_ net37 CIRCUIT_2223.tone_generator_2_1.GATES_10.input2 vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0995_ _0389_ _0451_ _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0780_ _0302_ _0300_ _0303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1263_ _0130_ net38 CIRCUIT_2223.tone_generator_2_1.GATES_16.input2 vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1194_ _0100_ net29 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_16.input2
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput5 io_in[3] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0978_ _0442_ _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0832_ _0345_ _0346_ _0090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0763_ net8 _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0901_ _0391_ _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0694_ _0225_ _0226_ _0229_ _0232_ _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_1177_ CIRCUIT_2223.tone_generator_1.MEMORY_14.s_currentState net15 CIRCUIT_2223.GATES_4.input1\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1246_ CIRCUIT_2223.tone_generator_2_1.MEMORY_31.d _0036_ CIRCUIT_2223.tone_generator_2_1.MEMORY_30.s_currentState
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_31.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_0_19_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_6_Left_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1100_ _0517_ _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1031_ _0472_ _0473_ _0476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_16_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0746_ spi_dac_i_2.spi_dat_buff\[1\] _0068_ _0277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0815_ _0330_ _0331_ _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_48_Left_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0677_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.d CIRCUIT_2223.triangle_wave_generator_1.GATES_11.input2
+ _0216_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.s_currentState _0217_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1229_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.d CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState
+ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.s_currentState vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0600_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.s_currentState CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_21_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1014_ _0464_ _0465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0729_ _0262_ _0265_ _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0997__S _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout16 CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState net16 vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout49 CIRCUIT_2223.CLK net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout38 net40 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout27 net28 net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_24_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Left_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0994_ _0211_ _0451_ _0452_ _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_20_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0921__A1 _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0988__A1 _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0912__A1 _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1193_ _0099_ net29 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_15.input2
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1262_ _0129_ net37 CIRCUIT_2223.tone_generator_2_1.GATES_15.input2 vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput6 io_in[4] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0977_ _0440_ _0429_ _0442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0900_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_13.input2 _0158_ _0386_
+ _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0762_ spi_dac_i_2.spi_dat_buff\[11\] _0287_ _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0831_ spi_dac_i_2.spi_dat_buff\[10\] _0317_ _0306_ spi_dac_i_2.spi_dat_buff\[11\]
+ _0270_ _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_0693_ CIRCUIT_2223.tone_generator_2_1.MEMORY_28.s_currentState _0230_ _0231_ CIRCUIT_2223.tone_generator_2_1.MEMORY_30.s_currentState
+ _0232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_11_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0889__I net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_22_Left_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1176_ CIRCUIT_2223.tone_generator_1.MEMORY_17.s_currentState net15 CIRCUIT_2223.GATES_4.input1\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1245_ CIRCUIT_2223.tone_generator_2_1.MEMORY_30.d _0035_ CIRCUIT_2223.tone_generator_2_1.MEMORY_29.s_currentState
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_30.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_0_42_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1030_ _0475_ _0038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0814_ _0149_ CIRCUIT_2223.GATES_4.input1\[3\] CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.s_currentState
+ _0159_ _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_16_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0745_ _0276_ _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0676_ CIRCUIT_2223.triangle_wave_generator_1.GATES_10.input2 _0216_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1228_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.d CIRCUIT_2223.triangle_wave_generator_1.GATES_27.result
+ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1159_ _0085_ net50 spi_dac_i_2.spi_dat_buff\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0992__I _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1013_ _0174_ CIRCUIT_2223.tone_generator_2_1.GATES_27.result _0463_ net39 _0464_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_12_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0728_ _0263_ _0264_ _0265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0659_ _0199_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_27.result vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_35_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1043__I0 _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0897__I _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input4_I io_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout17 net18 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout28 net31 net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout39 net40 net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0993_ _0376_ _0451_ _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0921__A2 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_27.result
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1261_ _0128_ net38 CIRCUIT_2223.tone_generator_2_1.GATES_14.input2 vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1192_ CIRCUIT_2223.tone_generator_1.MEMORY_19.s_currentState _0010_ net20 CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput7 io_in[5] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0976_ _0441_ _0029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_40_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0830_ _0340_ _0342_ _0269_ _0338_ _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_22_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0761_ _0287_ _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0692_ CIRCUIT_2223.tone_generator_2_1.GATES_9.input2 _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1244_ CIRCUIT_2223.tone_generator_2_1.MEMORY_29.d _0034_ CIRCUIT_2223.tone_generator_2_1.MEMORY_28.s_currentState
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_29.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1175_ CIRCUIT_2223.tone_generator_1.MEMORY_19.s_currentState net15 CIRCUIT_2223.GATES_4.input1\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0959_ _0431_ _0022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0813_ _0320_ _0321_ CIRCUIT_2223.GATES_4.input1\[3\] CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.s_currentState
+ _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_3_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0744_ _0262_ _0263_ _0268_ _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_0675_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.d CIRCUIT_2223.triangle_wave_generator_1.GATES_12.input2
+ CIRCUIT_2223.triangle_wave_generator_1.GATES_14.input2 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.d
+ _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_24_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1158_ _0084_ net56 spi_dac_i_2.spi_dat_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1227_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.clock _0032_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.s_currentState
+ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_38.s_currentState vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_1089_ _0511_ _0050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_7_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1012_ _0154_ _0462_ _0463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0727_ spi_dac_i_2.counter\[3\] spi_dac_i_2.counter\[4\] _0264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0658_ _0178_ _0180_ _0188_ _0198_ _0199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_TAPCELL_ROW_4_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0589_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0554__I0 _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_49_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0545__I0 _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout18 net23 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout29 net31 net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0992_ _0426_ _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1191_ CIRCUIT_2223.tone_generator_1.MEMORY_18.s_currentState _0009_ net21 CIRCUIT_2223.tone_generator_1.MEMORY_19.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_0_36_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput8 rst_n net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1260_ _0127_ net38 CIRCUIT_2223.tone_generator_2_1.GATES_13.input2 vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0975_ _0440_ _0436_ _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0760_ spi_dac_i_2.counter\[0\] _0286_ _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_36_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0691_ CIRCUIT_2223.tone_generator_2_1.GATES_7.input2 _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1174_ CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState
+ CIRCUIT_2223.GATES_4.input1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1243_ CIRCUIT_2223.tone_generator_2_1.MEMORY_28.d _0033_ CIRCUIT_2223.tone_generator_2_1.MEMORY_38.s_currentState
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_28.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_0958_ _0002_ _0430_ _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_0889_ net7 _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0812_ spi_dac_i_2.spi_dat_buff\[8\] _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0743_ _0265_ _0275_ _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0674_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.d CIRCUIT_2223.triangle_wave_generator_1.GATES_15.input2
+ CIRCUIT_2223.triangle_wave_generator_1.GATES_7.input2 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.d
+ _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1157_ _0083_ net56 spi_dac_i_2.spi_dat_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1226_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.d _0031_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.s_currentState
+ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.s_currentState vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_0_47_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1088_ _0510_ _0507_ _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_30_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1011_ CIRCUIT_2223.GATES_1.input1\[3\] _0424_ _0462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_28_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0726_ net8 _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0657_ _0189_ _0192_ _0195_ _0197_ _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_0588_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.s_currentState
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_4_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1209_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.d _0014_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.s_currentState
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.s_currentState vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_35_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_26_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout19 net23 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0709_ CIRCUIT_2223.tone_generator_2_2.MEMORY_34.d CIRCUIT_2223.tone_generator_2_2.GATES_13.input2
+ CIRCUIT_2223.tone_generator_2_2.GATES_8.input2 CIRCUIT_2223.tone_generator_2_2.MEMORY_29.d
+ _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_35_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0924__A1 _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0991_ _0249_ _0448_ _0450_ _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_26_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_39_Left_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1190_ CIRCUIT_2223.tone_generator_1.MEMORY_17.s_currentState _0008_ net20 CIRCUIT_2223.tone_generator_1.MEMORY_18.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_0974_ _0367_ _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_40_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0690_ CIRCUIT_2223.tone_generator_2_1.MEMORY_35.s_currentState _0227_ _0228_ CIRCUIT_2223.tone_generator_2_1.MEMORY_31.s_currentState
+ _0229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1173_ net16 net18 CIRCUIT_2223.tone_generator_1.MEMORY_4.s_currentState vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1242_ _0121_ net32 CIRCUIT_2223.triangle_wave_generator_1.GATES_7.input2 vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0888_ _0183_ _0375_ _0382_ _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0957_ _0429_ _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_26_Left_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0811_ _0294_ _0327_ _0328_ _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0742_ spi_dac_i_2.counter\[3\] _0273_ spi_dac_i_2.counter\[4\] _0275_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0673_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.s_currentState _0211_ _0212_
+ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState _0213_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_24_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1156_ _0082_ net27 CIRCUIT_2223.triangle_wave_generator_1.GATES_10.input2 vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1225_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.d _0030_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.s_currentState
+ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.s_currentState vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_1087_ _0471_ _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_38_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1010_ _0461_ _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0725_ spi_dac_i_2.counter\[0\] _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0656_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState
+ _0196_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_10.input2 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.d
+ _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_4_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0587_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.s_currentState
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1208_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.d _0013_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.s_currentState
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.s_currentState vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XTAP_TAPCELL_ROW_35_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1139_ _0536_ _0065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_32_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0639_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.d CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_13.input2
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_10.input2 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.d
+ _0179_ _0180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XPHY_EDGE_ROW_13_Left_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0708_ CIRCUIT_2223.tone_generator_2_2.MEMORY_34.s_currentState _0245_ CIRCUIT_2223.tone_generator_2_2.GATES_17.input2
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_28.clock _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_23_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_46_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0990_ _0381_ _0448_ _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I io_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0973_ _0439_ _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1241_ _0120_ net32 CIRCUIT_2223.triangle_wave_generator_1.GATES_17.input2 vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1172_ _0098_ net53 CIRCUIT_2223.CLK vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0956_ _0428_ _0429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0887_ _0381_ _0377_ _0382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_1_Left_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0810_ spi_dac_i_2.spi_dat_buff\[7\] _0317_ _0305_ spi_dac_i_2.spi_dat_buff\[8\]
+ _0292_ _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_0741_ _0265_ _0274_ _0071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0672_ CIRCUIT_2223.triangle_wave_generator_1.GATES_12.input2 _0212_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1224_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.d _0029_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.s_currentState
+ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.s_currentState vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_1155_ _0081_ net34 CIRCUIT_2223.triangle_wave_generator_1.GATES_9.input2 vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1086_ _0509_ _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0939_ _0417_ _0414_ _0418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_43_Left_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0655_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_11.input2 _0196_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0586_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0724_ _0261_ CIRCUIT_2223.tone_generator_2_2.GATES_27.result vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_4_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1207_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.d _0012_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.s_currentState
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.s_currentState vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_1138_ _0536_ _0064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1069_ _0059_ _0403_ _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_38_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0707_ CIRCUIT_2223.tone_generator_2_2.GATES_13.input2 _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0569_ CIRCUIT_2223.MEMORY_26.s_currentState CIRCUIT_2223.MEMORY_18.clock vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0638_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.clock CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_17.input2
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_7.input2 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.d
+ _0179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_0_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_23_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_30_Left_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0726__I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0914__I0 _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0972_ _0434_ _0436_ _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_14_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1171_ _0097_ net52 slow_clock\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1240_ _0119_ net32 CIRCUIT_2223.triangle_wave_generator_1.GATES_16.input2 vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0886_ net6 _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0955_ CIRCUIT_2223.GATES_11.result _0219_ _0427_ _0059_ _0428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__0990__A1 _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0740_ spi_dac_i_2.counter\[3\] _0273_ _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_0671_ CIRCUIT_2223.triangle_wave_generator_1.GATES_11.input2 _0211_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1223_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.d _0028_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState
+ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.s_currentState vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_1154_ _0080_ net32 CIRCUIT_2223.triangle_wave_generator_1.GATES_8.input2 vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1085_ _0504_ _0507_ _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_0869_ _0368_ _0370_ _0006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0938_ _0401_ _0417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_15_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_29_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0723_ _0243_ _0244_ _0254_ _0260_ _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_0654_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.s_currentState
+ _0193_ _0194_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.s_currentState
+ _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_0585_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.s_currentState
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1137_ _0369_ _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1206_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.clock _0011_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.s_currentState
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_38.s_currentState vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_0_28_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1068_ _0230_ _0494_ _0497_ _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1104__A1 _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0706_ CIRCUIT_2223.tone_generator_2_2.MEMORY_36.s_currentState CIRCUIT_2223.tone_generator_2_2.GATES_15.input2
+ _0244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_0637_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_8.input2 _0178_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_0568_ _0152_ _0173_ _0001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0999__I1 _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0971_ _0438_ _0027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1170_ _0096_ net52 slow_clock\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0885_ _0181_ _0375_ _0380_ _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0954_ net42 _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1299_ CIRCUIT_2223.MEMORY_22.d _0063_ CIRCUIT_2223.MEMORY_21.s_currentState CIRCUIT_2223.MEMORY_22.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_0_18_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0670_ _0204_ _0207_ _0208_ _0209_ _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_24_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1153_ _0079_ net55 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1222_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.d _0027_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.s_currentState
+ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_1084_ _0508_ _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_15_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0799_ spi_dac_i_2.spi_dat_buff\[6\] _0317_ _0306_ spi_dac_i_2.spi_dat_buff\[7\]
+ _0270_ _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_0868_ _0368_ _0370_ _0005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0937_ _0416_ _0016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0890__A1 _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0653_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_14.input2 _0194_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0722_ _0255_ _0256_ _0258_ _0259_ _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_0584_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.s_currentState
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1205_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.d CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_27.result
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1136_ _0535_ _0063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1067_ _0383_ _0494_ _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__0881__A1 _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0636_ _0177_ CIRCUIT_2223.tone_generator_1.GATES_3.result vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0705_ CIRCUIT_2223.tone_generator_2_2.MEMORY_37.s_currentState _0241_ CIRCUIT_2223.tone_generator_2_2.GATES_8.input2
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_29.d _0242_ _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_0_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0567_ _0169_ _0172_ _0173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_23_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1119_ _0527_ _0529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_46_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0845__A1 _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1013__A1 _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_17_Left_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_20_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0619_ CIRCUIT_2223.tone_generator_2_2.MEMORY_39.s_currentState CIRCUIT_2223.tone_generator_2_2.MEMORY_39.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_42_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0970_ _0434_ _0436_ _0438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_26_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0884_ _0379_ _0377_ _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0953_ _0396_ _0297_ _0426_ _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1298_ CIRCUIT_2223.GATES_11.input2 _0062_ CIRCUIT_2223.MEMORY_22.s_currentState
+ CIRCUIT_2223.MEMORY_23.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_0_33_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1221_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.d _0026_ net25 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_1152_ _0078_ net56 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1083_ _0504_ _0507_ _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_0936_ _0411_ _0414_ _0416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_15_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0798_ _0287_ _0317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0867_ _0368_ _0370_ _0004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_38_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_5_Left_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0652_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_12.input2 _0193_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0583_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.s_currentState
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0721_ CIRCUIT_2223.tone_generator_2_2.MEMORY_32.d CIRCUIT_2223.tone_generator_2_2.GATES_11.input2
+ _0249_ CIRCUIT_2223.tone_generator_2_2.MEMORY_31.s_currentState _0259_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1204_ _0110_ net36 CIRCUIT_2223.GATES_1.input1\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1066_ _0496_ _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1135_ _0535_ _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_47_Left_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0919_ _0152_ _0403_ _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_3_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0635_ net16 CIRCUIT_2223.tone_generator_1.MEMORY_9.s_currentState _0177_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0566_ _0168_ _0153_ _0172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0704_ CIRCUIT_2223.tone_generator_2_2.MEMORY_33.d CIRCUIT_2223.tone_generator_2_2.GATES_12.input2
+ _0241_ CIRCUIT_2223.tone_generator_2_2.MEMORY_37.s_currentState _0242_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1118_ _0528_ _0140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1049_ _0403_ _0425_ _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_35_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0542__A1 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_20_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0549_ CIRCUIT_2223.GATES_5.input2 _0159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0618_ CIRCUIT_2223.tone_generator_2_1.MEMORY_38.s_currentState CIRCUIT_2223.tone_generator_2_1.MEMORY_28.clock
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_34_Left_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0993__A1 _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0952_ _0154_ _0425_ _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_12_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0883_ net5 _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1297_ CIRCUIT_2223.MEMORY_24.d _0061_ CIRCUIT_2223.GATES_11.result CIRCUIT_2223.MEMORY_24.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_18_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1151_ _0077_ net58 spi_dac_i_2.spi_dat_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1220_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.d _0025_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.s_currentState
+ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.s_currentState vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_1082_ _0499_ _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0866_ _0368_ _0370_ _0003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0935_ _0415_ _0015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_15_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_21_Left_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0797_ _0309_ _0314_ _0315_ _0316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_46_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0720_ CIRCUIT_2223.tone_generator_2_2.MEMORY_32.s_currentState _0257_ CIRCUIT_2223.tone_generator_2_2.GATES_12.input2
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_33.d _0258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_0582_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.s_currentState
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0651_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.s_currentState
+ _0190_ _0191_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.s_currentState
+ _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__0579__I _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1203_ _0109_ net29 CIRCUIT_2223.GATES_1.input1\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1134_ _0535_ _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1065_ CIRCUIT_2223.tone_generator_2_1.GATES_17.input2 _0302_ _0492_ _0496_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0849_ slow_clock\[4\] _0355_ _0307_ _0359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0918_ _0169_ _0167_ _0153_ _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_38_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0862__I _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0703_ CIRCUIT_2223.tone_generator_2_2.GATES_16.input2 _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0634_ _0176_ CIRCUIT_2223.tone_generator_1.GATES_2.result vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0565_ _0152_ _0171_ _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1117_ _0295_ CIRCUIT_2223.tone_generator_2_2.GATES_15.input2 _0527_ _0528_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_0_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1048_ _0485_ _0124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0542__A2 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0617_ CIRCUIT_2223.tone_generator_2_1.MEMORY_37.s_currentState CIRCUIT_2223.tone_generator_2_1.MEMORY_37.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0548_ _0157_ _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0870__I _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0882_ _0190_ _0375_ _0378_ _0099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0951_ CIRCUIT_2223.GATES_1.input1\[3\] _0424_ _0425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1296_ CIRCUIT_2223.MEMORY_25.d _0060_ net24 CIRCUIT_2223.MEMORY_25.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_0_24_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1150_ _0076_ net57 spi_dac_i_2.spi_dat_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1081_ _0506_ _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0865_ _0369_ _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0934_ _0411_ _0414_ _0415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_15_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1070__A1 _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0796_ _0159_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_42.s_currentState _0315_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1279_ _0134_ net37 CIRCUIT_2223.tone_generator_2_1.GATES_9.input2 vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0884__A1 _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0581_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.s_currentState
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.d vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0650_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_7.input2 _0191_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1133_ _0535_ _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1064_ _0220_ _0494_ _0495_ _0130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1202_ _0108_ net30 CIRCUIT_2223.GATES_1.input1\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0848_ slow_clock\[4\] _0355_ _0358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_43_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0917_ _0401_ _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0779_ _0157_ _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_3_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0633_ net16 CIRCUIT_2223.tone_generator_1.MEMORY_7.s_currentState _0176_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_0702_ _0240_ CIRCUIT_2223.tone_generator_2_1.GATES_27.result vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0564_ _0168_ _0170_ _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_48_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1212__CLK net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1047_ _0158_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_10.input2 _0482_
+ _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1116_ _0173_ _0445_ _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_31_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1016__A1 _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0550__I0 _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1007__A1 _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_20_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0616_ CIRCUIT_2223.tone_generator_2_1.MEMORY_36.s_currentState CIRCUIT_2223.tone_generator_2_1.MEMORY_36.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0547_ net6 _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0881_ _0376_ _0377_ _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0950_ net3 net2 CIRCUIT_2223.GATES_1.input1\[2\] _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1295_ CIRCUIT_2223.MEMORY_18.clock _0059_ CIRCUIT_2223.MEMORY_25.s_currentState
+ CIRCUIT_2223.MEMORY_26.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1080_ _0504_ _0501_ _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1290__CLKN _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0795_ _0149_ CIRCUIT_2223.GATES_4.input1\[1\] _0314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0864_ _0363_ _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0933_ _0406_ _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_23_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1278_ _0133_ net36 CIRCUIT_2223.tone_generator_2_1.GATES_8.input2 vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0580_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_38.s_currentState
+ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.clock vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1201_ _0107_ net41 CIRCUIT_2223.GATES_1.input1\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1132_ _0369_ _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1063_ _0389_ _0494_ _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0916_ _0366_ _0401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0847_ _0357_ _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0778_ _0206_ _0300_ _0301_ _0081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_3_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_9_Left_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_26_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0632_ _0175_ CIRCUIT_2223.tone_generator_1.GATES_1.result vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0701_ _0222_ _0223_ _0233_ _0239_ _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_0563_ _0169_ _0153_ _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_20_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1046_ _0184_ _0482_ _0484_ _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1115_ _0248_ _0522_ _0526_ _0139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_31_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0546_ _0156_ _0147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0615_ CIRCUIT_2223.tone_generator_2_1.MEMORY_35.s_currentState CIRCUIT_2223.tone_generator_2_1.MEMORY_35.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1029_ _0472_ _0473_ _0475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_31_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0974__I _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0902__A1 _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_38_Left_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0880_ _0374_ _0377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0879__I net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1294_ _0147_ _0058_ net42 CIRCUIT_2223.s_logisimNet48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_32_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0932_ _0413_ _0014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0794_ _0312_ _0313_ _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0863_ _0354_ _0368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_23_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1277_ CIRCUIT_2223.tone_generator_2_2.MEMORY_39.d CIRCUIT_2223.tone_generator_2_2.GATES_27.result
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_39.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1290__D net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1200_ _0106_ net28 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_14.input2
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1131_ _0533_ _0534_ _0058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1062_ _0492_ _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_25_Left_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0915_ _0400_ _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0846_ _0353_ _0356_ _0357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_11_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0777_ _0162_ _0300_ _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_3_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0700_ _0234_ _0235_ _0237_ _0238_ _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_0631_ CIRCUIT_2223.tone_generator_1.MEMORY_6.s_currentState net16 _0175_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_0562_ CIRCUIT_2223.GATES_1.input1\[0\] _0169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_20_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1114_ net7 _0521_ _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1045_ _0161_ _0482_ _0484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0829_ _0294_ _0343_ _0344_ _0089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_31_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0545_ _0148_ _0149_ _0155_ _0156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0614_ CIRCUIT_2223.tone_generator_2_1.MEMORY_34.s_currentState CIRCUIT_2223.tone_generator_2_1.MEMORY_34.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1028_ _0474_ _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Left_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1293_ _0146_ _0057_ net42 CIRCUIT_2223.GATES_5.input2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_10_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1073__A1 _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0887__A1 _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_9_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0862_ _0367_ _0002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0931_ _0411_ _0408_ _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_23_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0793_ spi_dac_i_2.spi_dat_buff\[5\] _0288_ _0306_ spi_dac_i_2.spi_dat_buff\[6\]
+ _0270_ _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_2_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1276_ CIRCUIT_2223.tone_generator_2_2.MEMORY_28.clock _0054_ CIRCUIT_2223.tone_generator_2_2.MEMORY_37.s_currentState
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_38.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_0_3_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_0_Left_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1060__I1 _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1130_ _0533_ _0534_ _0057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1061_ _0493_ _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0845_ _0354_ _0355_ _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0914_ _0148_ CIRCUIT_2223.GATES_1.input1\[3\] _0394_ _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_11_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0776_ _0298_ _0300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1259_ _0126_ net39 CIRCUIT_2223.tone_generator_2_1.GATES_12.input2 vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_42_Left_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0561_ _0167_ _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0630_ CIRCUIT_2223.tone_generator_2_2.MEMORY_38.s_currentState CIRCUIT_2223.tone_generator_2_2.MEMORY_28.clock
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1044_ _0483_ _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1113_ _0245_ _0522_ _0525_ _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0828_ spi_dac_i_2.spi_dat_buff\[9\] _0317_ _0305_ spi_dac_i_2.spi_dat_buff\[10\]
+ _0292_ _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_0759_ spi_dac_i_2.counter\[3\] spi_dac_i_2.counter\[4\] _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_31_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1302__CLKN CIRCUIT_2223.MEMORY_18.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0613_ CIRCUIT_2223.tone_generator_2_1.MEMORY_33.s_currentState CIRCUIT_2223.tone_generator_2_1.MEMORY_33.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0544_ _0152_ _0154_ _0155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1027_ _0472_ _0473_ _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_48_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1292_ _0145_ _0056_ net43 CIRCUIT_2223.GATES_3.input2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_18_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_9_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0792_ _0309_ _0311_ _0269_ _0312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0861_ _0366_ _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0930_ _0412_ _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1275_ CIRCUIT_2223.tone_generator_2_2.MEMORY_37.d _0053_ CIRCUIT_2223.tone_generator_2_2.MEMORY_36.s_currentState
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_37.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XTAP_TAPCELL_ROW_37_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1060_ CIRCUIT_2223.tone_generator_2_1.GATES_15.input2 _0295_ _0492_ _0493_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0844_ slow_clock\[0\] slow_clock\[1\] slow_clock\[2\] slow_clock\[3\] _0355_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0913_ _0150_ _0397_ _0399_ _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0775_ _0299_ _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1189_ CIRCUIT_2223.tone_generator_1.MEMORY_16.s_currentState _0007_ net21 CIRCUIT_2223.tone_generator_1.MEMORY_17.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_1258_ _0125_ net40 CIRCUIT_2223.tone_generator_2_1.GATES_11.input2 vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0950__A1 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1205__CLK CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_27.result
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0560_ CIRCUIT_2223.GATES_1.input1\[1\] _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_45_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1043_ _0295_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_8.input2 _0482_
+ _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1112_ _0157_ _0521_ _0525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_31_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0758_ net11 _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0827_ _0340_ _0342_ _0343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_3_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0689_ CIRCUIT_2223.tone_generator_2_1.GATES_10.input2 _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0774__I1 _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0953__B _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0612_ CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState CIRCUIT_2223.tone_generator_2_1.MEMORY_32.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input7_I io_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0543_ CIRCUIT_2223.GATES_1.input1\[0\] CIRCUIT_2223.GATES_1.input1\[1\] _0153_ _0154_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_48_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1026_ _0464_ _0473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_31_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0905__A1 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1009_ _0148_ CIRCUIT_2223.triangle_wave_generator_1.GATES_7.input2 _0456_ _0461_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_12_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1291_ _0144_ _0055_ net43 CIRCUIT_2223.GATES_2.input2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_18_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0791_ _0310_ _0311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0860_ _0290_ _0363_ _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_23_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1274_ CIRCUIT_2223.tone_generator_2_2.MEMORY_36.d _0052_ CIRCUIT_2223.tone_generator_2_2.MEMORY_35.s_currentState
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_36.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_0_46_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0989_ _0252_ _0448_ _0449_ _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_6_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0912_ _0381_ _0397_ _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0843_ _0290_ _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0774_ CIRCUIT_2223.triangle_wave_generator_1.GATES_8.input2 _0295_ _0298_ _0299_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1188_ CIRCUIT_2223.tone_generator_1.MEMORY_15.s_currentState _0006_ net20 CIRCUIT_2223.tone_generator_1.MEMORY_16.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_1257_ _0124_ net26 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_10.input2
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0950__A2 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_29_Left_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1042_ _0404_ _0482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1111_ _0524_ _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1009__I0 _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0757_ _0283_ _0284_ _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0826_ _0331_ _0341_ _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0688_ CIRCUIT_2223.tone_generator_2_1.GATES_14.input2 _0227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0611_ CIRCUIT_2223.tone_generator_2_1.MEMORY_31.s_currentState CIRCUIT_2223.tone_generator_2_1.MEMORY_31.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0542_ net3 net2 _0153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_1025_ _0471_ _0472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0809_ _0323_ _0326_ _0327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_31_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_16_Left_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1008_ _0205_ _0458_ _0460_ _0120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1067__A1 _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1290_ net4 _0000_ net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XTAP_TAPCELL_ROW_18_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0790_ _0149_ CIRCUIT_2223.GATES_4.input1\[0\] CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState
+ _0159_ _0310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_2_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1273_ CIRCUIT_2223.tone_generator_2_2.MEMORY_35.d _0051_ CIRCUIT_2223.tone_generator_2_2.MEMORY_34.s_currentState
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_35.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XTAP_TAPCELL_ROW_14_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0988_ _0379_ _0448_ _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0842_ _0352_ _0350_ _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0911_ _0396_ _0397_ _0398_ _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_11_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0773_ _0171_ _0297_ _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1256_ _0123_ net29 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_9.input2
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1187_ CIRCUIT_2223.tone_generator_1.MEMORY_14.s_currentState _0005_ net18 CIRCUIT_2223.tone_generator_1.MEMORY_15.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_46_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_4_Left_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_25_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1110_ _0162_ CIRCUIT_2223.tone_generator_2_2.GATES_12.input2 _0521_ _0524_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1041_ _0481_ _0043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0825_ _0323_ _0326_ _0330_ _0319_ _0341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0756_ spi_dac_i_2.spi_dat_buff\[5\] _0276_ _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0687_ CIRCUIT_2223.tone_generator_2_1.MEMORY_34.d CIRCUIT_2223.tone_generator_2_1.GATES_13.input2
+ CIRCUIT_2223.tone_generator_2_1.GATES_8.input2 CIRCUIT_2223.tone_generator_2_1.MEMORY_29.d
+ _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Left_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_39_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1239_ _0118_ net33 CIRCUIT_2223.triangle_wave_generator_1.GATES_15.input2 vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0610_ CIRCUIT_2223.tone_generator_2_1.MEMORY_30.s_currentState CIRCUIT_2223.tone_generator_2_1.MEMORY_30.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0541_ _0150_ _0151_ _0152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1024_ _0366_ _0471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0808_ _0309_ _0324_ _0325_ _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_21_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0739_ _0265_ _0272_ _0273_ _0070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1007_ _0381_ _0458_ _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Left_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0904__I net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1272_ CIRCUIT_2223.tone_generator_2_2.MEMORY_34.d _0050_ CIRCUIT_2223.tone_generator_2_2.MEMORY_33.s_currentState
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_34.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_0987_ _0446_ _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_6_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0841_ slow_clock\[3\] _0352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0772_ _0296_ _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0910_ _0379_ _0397_ _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1186_ CIRCUIT_2223.tone_generator_1.MEMORY_13.s_currentState _0004_ net20 CIRCUIT_2223.tone_generator_1.MEMORY_14.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1255_ _0122_ net27 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_8.input2
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_20_Left_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_25_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0926__A1 _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1040_ _0478_ _0465_ _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_28_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0755_ spi_dac_i_2.spi_dat_buff\[4\] _0266_ _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0824_ _0338_ _0339_ _0340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0686_ CIRCUIT_2223.tone_generator_2_1.MEMORY_34.s_currentState _0224_ CIRCUIT_2223.tone_generator_2_1.GATES_17.input2
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_28.clock _0225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1169_ _0095_ net52 slow_clock\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1238_ _0117_ net26 CIRCUIT_2223.triangle_wave_generator_1.GATES_14.input2 vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0540_ net3 net2 CIRCUIT_2223.GATES_1.input1\[3\] _0151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_21_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1023_ _0470_ _0036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0807_ _0320_ _0321_ CIRCUIT_2223.GATES_4.input1\[1\] net14 _0325_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_0738_ _0262_ spi_dac_i_2.counter\[1\] spi_dac_i_2.counter\[2\] _0273_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_24_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0669_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.d CIRCUIT_2223.triangle_wave_generator_1.GATES_13.input2
+ CIRCUIT_2223.triangle_wave_generator_1.GATES_16.input2 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.d
+ _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_42_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input5_I io_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1006_ _0203_ _0458_ _0459_ _0119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__0578__A2 net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1271_ CIRCUIT_2223.tone_generator_2_2.MEMORY_33.d _0049_ CIRCUIT_2223.tone_generator_2_2.MEMORY_32.s_currentState
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_33.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0986_ _0447_ _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_6_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0840_ _0349_ _0351_ _0093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_11_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0771_ CIRCUIT_2223.GATES_1.input1\[2\] _0151_ _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1185_ CIRCUIT_2223.tone_generator_1.MEMORY_12.s_currentState _0003_ net19 CIRCUIT_2223.tone_generator_1.MEMORY_13.s_currentState
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_1254_ CIRCUIT_2223.tone_generator_2_1.MEMORY_39.d CIRCUIT_2223.tone_generator_2_1.GATES_27.result
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_39.s_currentState vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_34_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0969_ _0437_ _0026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_2_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0754_ _0281_ _0282_ _0076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0823_ CIRCUIT_2223.GATES_2.input2 CIRCUIT_2223.tone_generator_2_2.MEMORY_39.s_currentState
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_39.s_currentState CIRCUIT_2223.GATES_3.input2
+ _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_3_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0685_ CIRCUIT_2223.tone_generator_2_1.GATES_13.input2 _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1168_ _0094_ net51 slow_clock\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1099_ CIRCUIT_2223.tone_generator_2_1.GATES_8.input2 _0376_ _0516_ _0517_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1237_ _0116_ net27 CIRCUIT_2223.triangle_wave_generator_1.GATES_13.input2 vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1022_ _0422_ _0466_ _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_8_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0806_ _0320_ CIRCUIT_2223.GATES_4.input1\[1\] net14 _0321_ _0324_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_0737_ _0267_ spi_dac_i_2.counter\[1\] spi_dac_i_2.counter\[2\] _0272_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0668_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.d CIRCUIT_2223.triangle_wave_generator_1.GATES_14.input2
+ CIRCUIT_2223.triangle_wave_generator_1.GATES_9.input2 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.d
+ _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0599_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.s_currentState CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.d
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1005_ _0379_ _0458_ _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
.ends

