magic
tech gf180mcuD
magscale 1 10
timestamp 1698715248
<< nwell >>
rect 1258 146176 228678 146694
rect 1258 145447 19910 145472
rect 1258 144633 228678 145447
rect 1258 144608 17726 144633
rect 1258 143879 30326 143904
rect 1258 143065 228678 143879
rect 1258 143040 26406 143065
rect 1258 142311 12517 142336
rect 1258 141497 228678 142311
rect 1258 141472 29671 141497
rect 1258 140743 11566 140768
rect 1258 139929 228678 140743
rect 1258 139904 26863 139929
rect 1258 139175 13974 139200
rect 1258 138361 228678 139175
rect 1258 138336 9942 138361
rect 1258 137607 56758 137632
rect 1258 136793 228678 137607
rect 1258 136768 8654 136793
rect 1258 136039 25398 136064
rect 1258 135225 228678 136039
rect 1258 135200 31222 135225
rect 1258 134471 9718 134496
rect 1258 133657 228678 134471
rect 1258 133632 72801 133657
rect 1258 132903 41087 132928
rect 1258 132089 228678 132903
rect 1258 132064 7487 132089
rect 1258 131335 9727 131360
rect 1258 130521 228678 131335
rect 1258 130496 15878 130521
rect 1258 129767 12182 129792
rect 1258 128953 228678 129767
rect 1258 128928 10626 128953
rect 1258 128199 9718 128224
rect 1258 127385 228678 128199
rect 1258 127360 35959 127385
rect 1258 126631 12462 126656
rect 1258 125817 228678 126631
rect 1258 125792 7478 125817
rect 1258 125063 11286 125088
rect 1258 124249 228678 125063
rect 1258 124224 9494 124249
rect 1258 123495 36542 123520
rect 1258 122681 228678 123495
rect 1258 122656 11398 122681
rect 1258 121927 8162 121952
rect 1258 121113 228678 121927
rect 1258 121088 7814 121113
rect 1258 120359 17558 120384
rect 1258 119545 228678 120359
rect 1258 119520 7982 119545
rect 1258 118791 10175 118816
rect 1258 117977 228678 118791
rect 1258 117952 21814 117977
rect 1258 117223 15430 117248
rect 1258 116409 228678 117223
rect 1258 116384 24726 116409
rect 1258 115655 18575 115680
rect 1258 114841 228678 115655
rect 1258 114816 15542 114841
rect 1258 114087 13918 114112
rect 1258 113273 228678 114087
rect 1258 113248 22934 113273
rect 1258 112519 8206 112544
rect 1258 111705 228678 112519
rect 1258 111680 14775 111705
rect 1258 110951 9952 110976
rect 1258 110137 228678 110951
rect 1258 110112 22108 110137
rect 1258 109383 43822 109408
rect 1258 108569 228678 109383
rect 1258 108544 18109 108569
rect 1258 107815 6461 107840
rect 1258 107001 228678 107815
rect 1258 106976 9933 107001
rect 1258 106247 3437 106272
rect 1258 105433 228678 106247
rect 1258 105408 24157 105433
rect 1258 104679 2541 104704
rect 1258 103865 228678 104679
rect 1258 103840 34526 103865
rect 1258 103111 2765 103136
rect 1258 102297 228678 103111
rect 1258 102272 9973 102297
rect 1258 101543 10061 101568
rect 1258 100729 228678 101543
rect 1258 100704 2541 100729
rect 1258 99975 7366 100000
rect 1258 99161 228678 99975
rect 1258 99136 32333 99161
rect 1258 98407 20540 98432
rect 1258 97593 228678 98407
rect 1258 97568 10278 97593
rect 1258 96839 9727 96864
rect 1258 96025 228678 96839
rect 1258 96000 6836 96025
rect 1258 95271 2541 95296
rect 1258 94457 228678 95271
rect 1258 94432 18252 94457
rect 1258 93703 20380 93728
rect 1258 92889 228678 93703
rect 1258 92864 32109 92889
rect 1258 92135 2541 92160
rect 1258 91321 228678 92135
rect 1258 91296 47341 91321
rect 1258 90567 27741 90592
rect 1258 89753 228678 90567
rect 1258 89728 32333 89753
rect 1258 88999 46109 89024
rect 1258 88185 228678 88999
rect 1258 88160 16773 88185
rect 1258 87431 2541 87456
rect 1258 86617 228678 87431
rect 1258 86592 16681 86617
rect 1258 85863 2765 85888
rect 1258 85049 228678 85863
rect 1258 85024 111965 85049
rect 1258 84295 19966 84320
rect 1258 83481 228678 84295
rect 1258 83456 2541 83481
rect 1258 82727 17567 82752
rect 1258 81913 228678 82727
rect 1258 81888 29322 81913
rect 1258 81159 17901 81184
rect 1258 80345 228678 81159
rect 1258 80320 38605 80345
rect 1258 79591 19272 79616
rect 1258 78777 228678 79591
rect 1258 78752 11880 78777
rect 1258 78023 14749 78048
rect 1258 77209 228678 78023
rect 1258 77184 24157 77209
rect 1258 76455 20255 76480
rect 1258 75641 228678 76455
rect 1258 75616 18230 75641
rect 1258 74887 12406 74912
rect 1258 74073 228678 74887
rect 1258 74048 9277 74073
rect 1258 73319 3343 73344
rect 1258 72505 228678 73319
rect 1258 72480 4175 72505
rect 1258 71751 19518 71776
rect 1258 70937 228678 71751
rect 1258 70912 6134 70937
rect 1258 70183 9942 70208
rect 1258 69369 228678 70183
rect 1258 69344 9162 69369
rect 1258 68615 13694 68640
rect 1258 67801 228678 68615
rect 1258 67776 7254 67801
rect 1258 67047 3343 67072
rect 1258 66233 228678 67047
rect 1258 66208 9718 66233
rect 1258 65479 2606 65504
rect 1258 64665 228678 65479
rect 1258 64640 9942 64665
rect 1258 63911 13918 63936
rect 1258 63097 228678 63911
rect 1258 63072 7030 63097
rect 1258 62343 5014 62368
rect 1258 61529 228678 62343
rect 1258 61504 54417 61529
rect 1258 60775 17567 60800
rect 1258 59961 228678 60775
rect 1258 59936 1888 59961
rect 1258 59207 26759 59232
rect 1258 58393 228678 59207
rect 1258 58368 3390 58393
rect 1258 57639 17916 57664
rect 1258 56825 228678 57639
rect 1258 56800 2662 56825
rect 1258 56071 20156 56096
rect 1258 55257 228678 56071
rect 1258 55232 4242 55257
rect 1258 54503 15878 54528
rect 1258 53689 228678 54503
rect 1258 53664 13638 53689
rect 1258 52935 18252 52960
rect 1258 52121 228678 52935
rect 1258 52096 18286 52121
rect 1258 51367 28077 51392
rect 1258 50553 228678 51367
rect 1258 50528 2718 50553
rect 1258 49799 3567 49824
rect 1258 48985 228678 49799
rect 1258 48960 24977 48985
rect 1258 48231 10061 48256
rect 1258 47417 228678 48231
rect 1258 47392 80760 47417
rect 1258 46663 6255 46688
rect 1258 45849 228678 46663
rect 1258 45824 3816 45849
rect 1258 45095 6685 45120
rect 1258 44281 228678 45095
rect 1258 44256 15421 44281
rect 1258 43527 3592 43552
rect 1258 42713 228678 43527
rect 1258 42688 14330 42713
rect 1258 41959 10747 41984
rect 1258 41145 228678 41959
rect 1258 41120 2989 41145
rect 1258 40391 4669 40416
rect 1258 39577 228678 40391
rect 1258 39552 22141 39577
rect 1258 38823 2541 38848
rect 1258 38009 228678 38823
rect 1258 37984 8701 38009
rect 1258 37255 2541 37280
rect 1258 36441 228678 37255
rect 1258 36416 6461 36441
rect 1258 35687 6909 35712
rect 1258 34873 228678 35687
rect 1258 34848 2541 34873
rect 1258 34119 13112 34144
rect 1258 33305 228678 34119
rect 1258 33280 7917 33305
rect 1258 32551 2541 32576
rect 1258 31737 228678 32551
rect 1258 31712 10641 31737
rect 1258 30983 6685 31008
rect 1258 30169 228678 30983
rect 1258 30144 2653 30169
rect 1258 29415 12397 29440
rect 1258 28601 228678 29415
rect 1258 28576 2877 28601
rect 1258 27847 11316 27872
rect 1258 27033 228678 27847
rect 1258 27008 9149 27033
rect 1258 26279 5677 26304
rect 1258 25465 228678 26279
rect 1258 25440 2765 25465
rect 1258 24711 6939 24736
rect 1258 23897 228678 24711
rect 1258 23872 2653 23897
rect 1258 23143 6573 23168
rect 1258 22329 228678 23143
rect 1258 22304 2877 22329
rect 1258 21575 22141 21600
rect 1258 20761 228678 21575
rect 1258 20736 14301 20761
rect 1258 20007 2653 20032
rect 1258 19193 228678 20007
rect 1258 19168 10847 19193
rect 1258 18439 14749 18464
rect 1258 17625 228678 18439
rect 1258 17600 2541 17625
rect 1258 16871 5229 16896
rect 1258 16057 228678 16871
rect 1258 16032 10177 16057
rect 1258 15303 5341 15328
rect 1258 14489 228678 15303
rect 1258 14464 2541 14489
rect 1258 13735 35713 13760
rect 1258 12921 228678 13735
rect 1258 12896 16765 12921
rect 1258 12167 4109 12192
rect 1258 11353 228678 12167
rect 1258 11328 2541 11353
rect 1258 10599 3661 10624
rect 1258 9785 228678 10599
rect 1258 9760 17905 9785
rect 1258 9031 6013 9056
rect 1258 8217 228678 9031
rect 1258 8192 16225 8217
rect 1258 7463 26845 7488
rect 1258 6649 228678 7463
rect 1258 6624 7581 6649
rect 1258 5895 13629 5920
rect 1258 5081 228678 5895
rect 1258 5056 15757 5081
rect 1258 4327 11725 4352
rect 1258 3513 228678 4327
rect 1258 3488 59997 3513
<< pwell >>
rect 1258 145472 228678 146176
rect 1258 143904 228678 144608
rect 1258 142336 228678 143040
rect 1258 140768 228678 141472
rect 1258 139200 228678 139904
rect 1258 137632 228678 138336
rect 1258 136064 228678 136768
rect 1258 134496 228678 135200
rect 1258 132928 228678 133632
rect 1258 131360 228678 132064
rect 1258 129792 228678 130496
rect 1258 128224 228678 128928
rect 1258 126656 228678 127360
rect 1258 125088 228678 125792
rect 1258 123520 228678 124224
rect 1258 121952 228678 122656
rect 1258 120384 228678 121088
rect 1258 118816 228678 119520
rect 1258 117248 228678 117952
rect 1258 115680 228678 116384
rect 1258 114112 228678 114816
rect 1258 112544 228678 113248
rect 1258 110976 228678 111680
rect 1258 109408 228678 110112
rect 1258 107840 228678 108544
rect 1258 106272 228678 106976
rect 1258 104704 228678 105408
rect 1258 103136 228678 103840
rect 1258 101568 228678 102272
rect 1258 100000 228678 100704
rect 1258 98432 228678 99136
rect 1258 96864 228678 97568
rect 1258 95296 228678 96000
rect 1258 93728 228678 94432
rect 1258 92160 228678 92864
rect 1258 90592 228678 91296
rect 1258 89024 228678 89728
rect 1258 87456 228678 88160
rect 1258 85888 228678 86592
rect 1258 84320 228678 85024
rect 1258 82752 228678 83456
rect 1258 81184 228678 81888
rect 1258 79616 228678 80320
rect 1258 78048 228678 78752
rect 1258 76480 228678 77184
rect 1258 74912 228678 75616
rect 1258 73344 228678 74048
rect 1258 71776 228678 72480
rect 1258 70208 228678 70912
rect 1258 68640 228678 69344
rect 1258 67072 228678 67776
rect 1258 65504 228678 66208
rect 1258 63936 228678 64640
rect 1258 62368 228678 63072
rect 1258 60800 228678 61504
rect 1258 59232 228678 59936
rect 1258 57664 228678 58368
rect 1258 56096 228678 56800
rect 1258 54528 228678 55232
rect 1258 52960 228678 53664
rect 1258 51392 228678 52096
rect 1258 49824 228678 50528
rect 1258 48256 228678 48960
rect 1258 46688 228678 47392
rect 1258 45120 228678 45824
rect 1258 43552 228678 44256
rect 1258 41984 228678 42688
rect 1258 40416 228678 41120
rect 1258 38848 228678 39552
rect 1258 37280 228678 37984
rect 1258 35712 228678 36416
rect 1258 34144 228678 34848
rect 1258 32576 228678 33280
rect 1258 31008 228678 31712
rect 1258 29440 228678 30144
rect 1258 27872 228678 28576
rect 1258 26304 228678 27008
rect 1258 24736 228678 25440
rect 1258 23168 228678 23872
rect 1258 21600 228678 22304
rect 1258 20032 228678 20736
rect 1258 18464 228678 19168
rect 1258 16896 228678 17600
rect 1258 15328 228678 16032
rect 1258 13760 228678 14464
rect 1258 12192 228678 12896
rect 1258 10624 228678 11328
rect 1258 9056 228678 9760
rect 1258 7488 228678 8192
rect 1258 5920 228678 6624
rect 1258 4352 228678 5056
rect 1258 3050 228678 3488
<< obsm1 >>
rect 1344 3076 228592 146802
<< metal2 >>
rect 114912 149200 115024 150000
rect 57344 0 57456 800
rect 172256 0 172368 800
<< obsm2 >>
rect 1708 149140 114852 149200
rect 115084 149140 228452 149200
rect 1708 860 228452 149140
rect 1708 800 57284 860
rect 57516 800 172196 860
rect 172428 800 228452 860
<< metal3 >>
rect 229200 146048 230000 146160
rect 229200 143360 230000 143472
rect 229200 140672 230000 140784
rect 229200 137984 230000 138096
rect 229200 135296 230000 135408
rect 229200 132608 230000 132720
rect 229200 129920 230000 130032
rect 229200 127232 230000 127344
rect 229200 124544 230000 124656
rect 229200 121856 230000 121968
rect 229200 119168 230000 119280
rect 229200 116480 230000 116592
rect 229200 113792 230000 113904
rect 229200 111104 230000 111216
rect 229200 108416 230000 108528
rect 229200 105728 230000 105840
rect 229200 103040 230000 103152
rect 229200 100352 230000 100464
rect 229200 97664 230000 97776
rect 229200 94976 230000 95088
rect 229200 92288 230000 92400
rect 229200 89600 230000 89712
rect 229200 86912 230000 87024
rect 229200 84224 230000 84336
rect 229200 81536 230000 81648
rect 229200 78848 230000 78960
rect 229200 76160 230000 76272
rect 229200 73472 230000 73584
rect 229200 70784 230000 70896
rect 229200 68096 230000 68208
rect 229200 65408 230000 65520
rect 229200 62720 230000 62832
rect 229200 60032 230000 60144
rect 229200 57344 230000 57456
rect 229200 54656 230000 54768
rect 229200 51968 230000 52080
rect 229200 49280 230000 49392
rect 229200 46592 230000 46704
rect 229200 43904 230000 44016
rect 229200 41216 230000 41328
rect 229200 38528 230000 38640
rect 229200 35840 230000 35952
rect 229200 33152 230000 33264
rect 229200 30464 230000 30576
rect 229200 27776 230000 27888
rect 229200 25088 230000 25200
rect 229200 22400 230000 22512
rect 229200 19712 230000 19824
rect 229200 17024 230000 17136
rect 229200 14336 230000 14448
rect 229200 11648 230000 11760
rect 229200 8960 230000 9072
rect 229200 6272 230000 6384
rect 229200 3584 230000 3696
<< obsm3 >>
rect 1698 146220 229200 148820
rect 1698 145988 229140 146220
rect 1698 143532 229200 145988
rect 1698 143300 229140 143532
rect 1698 140844 229200 143300
rect 1698 140612 229140 140844
rect 1698 138156 229200 140612
rect 1698 137924 229140 138156
rect 1698 135468 229200 137924
rect 1698 135236 229140 135468
rect 1698 132780 229200 135236
rect 1698 132548 229140 132780
rect 1698 130092 229200 132548
rect 1698 129860 229140 130092
rect 1698 127404 229200 129860
rect 1698 127172 229140 127404
rect 1698 124716 229200 127172
rect 1698 124484 229140 124716
rect 1698 122028 229200 124484
rect 1698 121796 229140 122028
rect 1698 119340 229200 121796
rect 1698 119108 229140 119340
rect 1698 116652 229200 119108
rect 1698 116420 229140 116652
rect 1698 113964 229200 116420
rect 1698 113732 229140 113964
rect 1698 111276 229200 113732
rect 1698 111044 229140 111276
rect 1698 108588 229200 111044
rect 1698 108356 229140 108588
rect 1698 105900 229200 108356
rect 1698 105668 229140 105900
rect 1698 103212 229200 105668
rect 1698 102980 229140 103212
rect 1698 100524 229200 102980
rect 1698 100292 229140 100524
rect 1698 97836 229200 100292
rect 1698 97604 229140 97836
rect 1698 95148 229200 97604
rect 1698 94916 229140 95148
rect 1698 92460 229200 94916
rect 1698 92228 229140 92460
rect 1698 89772 229200 92228
rect 1698 89540 229140 89772
rect 1698 87084 229200 89540
rect 1698 86852 229140 87084
rect 1698 84396 229200 86852
rect 1698 84164 229140 84396
rect 1698 81708 229200 84164
rect 1698 81476 229140 81708
rect 1698 79020 229200 81476
rect 1698 78788 229140 79020
rect 1698 76332 229200 78788
rect 1698 76100 229140 76332
rect 1698 73644 229200 76100
rect 1698 73412 229140 73644
rect 1698 70956 229200 73412
rect 1698 70724 229140 70956
rect 1698 68268 229200 70724
rect 1698 68036 229140 68268
rect 1698 65580 229200 68036
rect 1698 65348 229140 65580
rect 1698 62892 229200 65348
rect 1698 62660 229140 62892
rect 1698 60204 229200 62660
rect 1698 59972 229140 60204
rect 1698 57516 229200 59972
rect 1698 57284 229140 57516
rect 1698 54828 229200 57284
rect 1698 54596 229140 54828
rect 1698 52140 229200 54596
rect 1698 51908 229140 52140
rect 1698 49452 229200 51908
rect 1698 49220 229140 49452
rect 1698 46764 229200 49220
rect 1698 46532 229140 46764
rect 1698 44076 229200 46532
rect 1698 43844 229140 44076
rect 1698 41388 229200 43844
rect 1698 41156 229140 41388
rect 1698 38700 229200 41156
rect 1698 38468 229140 38700
rect 1698 36012 229200 38468
rect 1698 35780 229140 36012
rect 1698 33324 229200 35780
rect 1698 33092 229140 33324
rect 1698 30636 229200 33092
rect 1698 30404 229140 30636
rect 1698 27948 229200 30404
rect 1698 27716 229140 27948
rect 1698 25260 229200 27716
rect 1698 25028 229140 25260
rect 1698 22572 229200 25028
rect 1698 22340 229140 22572
rect 1698 19884 229200 22340
rect 1698 19652 229140 19884
rect 1698 17196 229200 19652
rect 1698 16964 229140 17196
rect 1698 14508 229200 16964
rect 1698 14276 229140 14508
rect 1698 11820 229200 14276
rect 1698 11588 229140 11820
rect 1698 9132 229200 11588
rect 1698 8900 229140 9132
rect 1698 6444 229200 8900
rect 1698 6212 229140 6444
rect 1698 3756 229200 6212
rect 1698 3524 229140 3756
rect 1698 700 229200 3524
<< metal4 >>
rect 4448 3076 4768 146668
rect 19808 3076 20128 146668
rect 35168 3076 35488 146668
rect 50528 3076 50848 146668
rect 65888 3076 66208 146668
rect 81248 3076 81568 146668
rect 96608 3076 96928 146668
rect 111968 3076 112288 146668
rect 127328 3076 127648 146668
rect 142688 3076 143008 146668
rect 158048 3076 158368 146668
rect 173408 3076 173728 146668
rect 188768 3076 189088 146668
rect 204128 3076 204448 146668
rect 219488 3076 219808 146668
<< obsm4 >>
rect 7868 146728 226100 148830
rect 7868 3016 19748 146728
rect 20188 3016 35108 146728
rect 35548 3016 50468 146728
rect 50908 3016 65828 146728
rect 66268 3016 81188 146728
rect 81628 3016 96548 146728
rect 96988 3016 111908 146728
rect 112348 3016 127268 146728
rect 127708 3016 142628 146728
rect 143068 3016 157988 146728
rect 158428 3016 173348 146728
rect 173788 3016 188708 146728
rect 189148 3016 204068 146728
rect 204508 3016 219428 146728
rect 219868 3016 226100 146728
rect 7868 690 226100 3016
<< labels >>
rlabel metal3 s 229200 3584 230000 3696 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 229200 30464 230000 30576 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 229200 33152 230000 33264 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 229200 35840 230000 35952 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 229200 38528 230000 38640 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 229200 41216 230000 41328 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 229200 43904 230000 44016 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 229200 46592 230000 46704 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 229200 49280 230000 49392 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 229200 51968 230000 52080 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 229200 54656 230000 54768 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 229200 6272 230000 6384 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 229200 57344 230000 57456 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 229200 60032 230000 60144 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 229200 62720 230000 62832 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 229200 65408 230000 65520 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 229200 68096 230000 68208 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 229200 70784 230000 70896 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 229200 73472 230000 73584 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 229200 76160 230000 76272 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 229200 78848 230000 78960 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 229200 81536 230000 81648 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 229200 8960 230000 9072 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 229200 84224 230000 84336 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 229200 86912 230000 87024 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 229200 89600 230000 89712 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 229200 11648 230000 11760 6 io_in[3]
port 27 nsew signal input
rlabel metal3 s 229200 14336 230000 14448 6 io_in[4]
port 28 nsew signal input
rlabel metal3 s 229200 17024 230000 17136 6 io_in[5]
port 29 nsew signal input
rlabel metal3 s 229200 19712 230000 19824 6 io_in[6]
port 30 nsew signal input
rlabel metal3 s 229200 22400 230000 22512 6 io_in[7]
port 31 nsew signal input
rlabel metal3 s 229200 25088 230000 25200 6 io_in[8]
port 32 nsew signal input
rlabel metal3 s 229200 27776 230000 27888 6 io_in[9]
port 33 nsew signal input
rlabel metal2 s 114912 149200 115024 150000 6 io_oeb
port 34 nsew signal output
rlabel metal3 s 229200 92288 230000 92400 6 io_out[0]
port 35 nsew signal output
rlabel metal3 s 229200 119168 230000 119280 6 io_out[10]
port 36 nsew signal output
rlabel metal3 s 229200 121856 230000 121968 6 io_out[11]
port 37 nsew signal output
rlabel metal3 s 229200 124544 230000 124656 6 io_out[12]
port 38 nsew signal output
rlabel metal3 s 229200 127232 230000 127344 6 io_out[13]
port 39 nsew signal output
rlabel metal3 s 229200 129920 230000 130032 6 io_out[14]
port 40 nsew signal output
rlabel metal3 s 229200 132608 230000 132720 6 io_out[15]
port 41 nsew signal output
rlabel metal3 s 229200 135296 230000 135408 6 io_out[16]
port 42 nsew signal output
rlabel metal3 s 229200 137984 230000 138096 6 io_out[17]
port 43 nsew signal output
rlabel metal3 s 229200 140672 230000 140784 6 io_out[18]
port 44 nsew signal output
rlabel metal3 s 229200 143360 230000 143472 6 io_out[19]
port 45 nsew signal output
rlabel metal3 s 229200 94976 230000 95088 6 io_out[1]
port 46 nsew signal output
rlabel metal3 s 229200 146048 230000 146160 6 io_out[20]
port 47 nsew signal output
rlabel metal3 s 229200 97664 230000 97776 6 io_out[2]
port 48 nsew signal output
rlabel metal3 s 229200 100352 230000 100464 6 io_out[3]
port 49 nsew signal output
rlabel metal3 s 229200 103040 230000 103152 6 io_out[4]
port 50 nsew signal output
rlabel metal3 s 229200 105728 230000 105840 6 io_out[5]
port 51 nsew signal output
rlabel metal3 s 229200 108416 230000 108528 6 io_out[6]
port 52 nsew signal output
rlabel metal3 s 229200 111104 230000 111216 6 io_out[7]
port 53 nsew signal output
rlabel metal3 s 229200 113792 230000 113904 6 io_out[8]
port 54 nsew signal output
rlabel metal3 s 229200 116480 230000 116592 6 io_out[9]
port 55 nsew signal output
rlabel metal2 s 172256 0 172368 800 6 rst_n
port 56 nsew signal input
rlabel metal4 s 4448 3076 4768 146668 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 146668 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 65888 3076 66208 146668 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 96608 3076 96928 146668 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 127328 3076 127648 146668 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 158048 3076 158368 146668 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 188768 3076 189088 146668 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 219488 3076 219808 146668 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 146668 6 vss
port 58 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 146668 6 vss
port 58 nsew ground bidirectional
rlabel metal4 s 81248 3076 81568 146668 6 vss
port 58 nsew ground bidirectional
rlabel metal4 s 111968 3076 112288 146668 6 vss
port 58 nsew ground bidirectional
rlabel metal4 s 142688 3076 143008 146668 6 vss
port 58 nsew ground bidirectional
rlabel metal4 s 173408 3076 173728 146668 6 vss
port 58 nsew ground bidirectional
rlabel metal4 s 204128 3076 204448 146668 6 vss
port 58 nsew ground bidirectional
rlabel metal2 s 57344 0 57456 800 6 wb_clk_i
port 59 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 230000 150000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 30125198
string GDS_FILE /run/media/tholin/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1_group/openlane/wrapped_sid/runs/23_10_31_02_06/results/signoff/wrapped_sid.magic.gds
string GDS_START 553200
<< end >>

