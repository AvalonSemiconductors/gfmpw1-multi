* NGSPICE file created from wrapped_qcpu.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_4 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_4 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_2 I Z VDD VNW VPW VSS
.ends

.subckt wrapped_qcpu custom_settings[0] custom_settings[10] custom_settings[11] custom_settings[12]
+ custom_settings[13] custom_settings[14] custom_settings[15] custom_settings[16]
+ custom_settings[17] custom_settings[18] custom_settings[19] custom_settings[1] custom_settings[20]
+ custom_settings[21] custom_settings[22] custom_settings[23] custom_settings[24]
+ custom_settings[25] custom_settings[26] custom_settings[27] custom_settings[28]
+ custom_settings[29] custom_settings[2] custom_settings[30] custom_settings[31] custom_settings[3]
+ custom_settings[4] custom_settings[5] custom_settings[6] custom_settings[7] custom_settings[8]
+ custom_settings[9] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15]
+ io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23]
+ io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31]
+ io_in[32] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0]
+ io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17]
+ io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[24] io_oeb[25] io_oeb[26]
+ io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[3]
+ io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10]
+ io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18]
+ io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25]
+ io_out[27] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[3] io_out[4]
+ io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] rst_n sram_addr[0] sram_addr[1]
+ sram_addr[2] sram_addr[3] sram_addr[4] sram_addr[5] sram_gwe sram_in[0] sram_in[1]
+ sram_in[2] sram_in[3] sram_in[4] sram_in[5] sram_in[6] sram_in[7] sram_out[0] sram_out[1]
+ sram_out[2] sram_out[3] sram_out[4] sram_out[5] sram_out[6] sram_out[7] vdd vss
+ wb_clk_i io_oeb[22] io_oeb[23] io_out[28] io_out[26]
X_05903_ _00764_ _00957_ _01566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07534__A1 _02480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09671_ _00985_ _04012_ _04796_ _04797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06883_ cpu.timer\[6\] _02509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_68_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05834_ _01493_ _01495_ _01497_ _01498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08622_ cpu.orig_IO_addr_buff\[2\] _03864_ _03865_ _00919_ _03872_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08553_ _02394_ _03813_ _03814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05765_ _01149_ _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_77_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08484_ cpu.timer_capture\[12\] _03764_ _03758_ _03765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07504_ _02971_ _02987_ _02988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07435_ _01636_ _02911_ _02922_ _00694_ _00191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05696_ net80 _01357_ _01359_ _01361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_77_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07366_ _02860_ _02861_ _02862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09105_ _04305_ _04306_ _04110_ _04307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07297_ _02809_ _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_17_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06317_ _01955_ _01956_ _00745_ _01974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06248_ _01905_ _00021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_79_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09036_ _04070_ _02569_ _04240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06462__I _02105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05078__I _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06179_ cpu.timer_top\[15\] _01411_ _01252_ _01838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09938_ _00197_ clknet_leaf_41_wb_clk_i cpu.spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_5_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09869_ _00128_ clknet_leaf_96_wb_clk_i cpu.regs\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output37_I net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_104_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05697__B _01190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08073__B _03430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer7 _02128_ net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07417__B _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06567__A2 _02223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_60_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_60_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10009_ _00268_ clknet_leaf_33_wb_clk_i cpu.uart.receiving vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05550_ _01212_ _01214_ _01215_ _01216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05481_ _01115_ _01103_ _01146_ _00983_ _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_116_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07220_ _02763_ _02764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_109_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07151_ _02722_ _02714_ _02723_ _00106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06102_ _01047_ _01358_ net37 _01762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06282__I _01938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07082_ cpu.uart.receive_counter\[3\] _02679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06033_ _01670_ _01694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07984_ _03371_ _03375_ _00287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06935_ _02548_ _02549_ _02550_ _02551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07507__A1 cpu.timer_top\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09723_ _00873_ _01971_ _04839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09654_ _01037_ _04780_ _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06866_ _02470_ _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07507__B2 cpu.timer_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05817_ net8 _01370_ _01481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08605_ _03850_ _03856_ _01093_ _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06797_ _02434_ _02437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09585_ _02532_ _04718_ _04721_ _00542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08536_ _03798_ _03793_ _03800_ _00414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05748_ cpu.timer_top\[9\] _01247_ _01249_ _01413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05679_ _01314_ _01344_ _01345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08467_ _03740_ _03749_ _03750_ _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07418_ _02906_ _02907_ _02909_ _00187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_107_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08398_ _02974_ _03687_ _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07349_ _01752_ _02840_ _02847_ _00180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06246__A1 _01897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10291_ _00549_ clknet_leaf_60_wb_clk_i net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09019_ cpu.PC\[4\] _04190_ _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09735__A2 _04846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08068__B _03430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05080__S1 _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09671__A1 _00985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06324__I2 _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07926__I cpu.uart.receive_div_counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08531__B _03774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04981_ _00673_ _00681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06720_ _00579_ _01921_ _01922_ _02371_ _02372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_06651_ _00575_ _02303_ _02304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_65_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05602_ _01266_ _01267_ _01268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09370_ _02914_ _04558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06582_ _02182_ _02198_ _02202_ _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05533_ _01054_ _01199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09662__A1 _00674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08321_ cpu.timer_div_counter\[6\] _03630_ _03621_ _02404_ _03632_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_24_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07610__B _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05464_ _01031_ _01129_ _01130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08252_ _03584_ _02365_ _00346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07203_ _02756_ cpu.regs\[10\]\[6\] _02745_ _02757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05395_ _00994_ cpu.IO_addr_buff\[0\] _01061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_61_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08183_ cpu.toggle_top\[2\] _03532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_70_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07134_ _01352_ _02710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07065_ _02654_ _02657_ _02661_ _02664_ _02665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_76_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09717__A2 _01906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06016_ _01677_ _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07728__A1 _02440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05356__I _00615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07967_ cpu.uart.receive_div_counter\[7\] _03333_ _03361_ _03362_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06918_ cpu.timer_top\[5\] _02534_ _02537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09706_ _02818_ cpu.regs\[9\]\[4\] _04819_ _04827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07898_ _03308_ _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09637_ _02317_ _02324_ _04765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_87_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06849_ _01450_ _02480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09568_ _03833_ _04703_ _04709_ _00537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_93_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08519_ _02540_ _03783_ _03788_ _00409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_38_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09499_ _01014_ _04663_ _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_65_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10274_ _00532_ clknet_leaf_49_wb_clk_i cpu.PORTB_DDR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_49_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06942__A2 _01006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08695__A2 _00784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_14_Left_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_29_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08526__B _03774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06458__A1 _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06458__B2 _01730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_104_Right_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_83_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07258__I0 _02753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05180_ _00833_ _00851_ _00852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_24_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Left_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06560__I cpu.PC\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08870_ cpu.Z cpu.base_address\[4\] _04079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07821_ cpu.uart.has_byte _03246_ _03247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_71_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05176__I _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06933__A2 _01932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07752_ cpu.uart.div_counter\[2\] _03184_ _03190_ _03191_ _03192_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_04964_ _00663_ _00664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08135__A1 cpu.toggle_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06703_ _02329_ _02356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07683_ cpu.uart.div_counter\[7\] _02631_ _01583_ cpu.uart.div_counter\[3\] _03131_
+ _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08686__A2 _00748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04895_ _00590_ _00597_ _00598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_32_Left_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09422_ cpu.ROM_spi_dat_out\[0\] _04583_ _04601_ _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06634_ _02284_ _02285_ _02288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09353_ _04481_ _04541_ _04542_ _03398_ _00489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_94_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06565_ _02221_ _02222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08304_ _02944_ _03621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_4_5_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06449__A1 _02105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09284_ _02370_ _03809_ _04479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05516_ _01178_ _01180_ _01181_ _01182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_82_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06496_ _02147_ _02151_ _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08235_ _03497_ _03573_ _03574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05447_ _01106_ _01112_ _01113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_117_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05378_ _01036_ _01006_ _01043_ _01044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__05672__A2 _01335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08166_ cpu.toggle_ctr\[4\] _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07949__A1 _02662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07117_ cpu.regs\[13\]\[0\] _02700_ _02701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_41_Left_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08097_ _02210_ _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07048_ cpu.uart.divisor\[12\] _02648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_11_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08999_ _00747_ _04166_ _04204_ _04205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08126__A1 cpu.toggle_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08397__I _03621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_117_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_117_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_57_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06160__I0 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08860__I cpu.PC\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10326_ net49 net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10257_ _00515_ clknet_leaf_45_wb_clk_i net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_56_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08365__A1 _02998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10188_ _00446_ clknet_leaf_72_wb_clk_i cpu.ROM_addr_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_56_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06350_ _02006_ _02004_ _02007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_72_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06281_ _00983_ _01312_ _00674_ _01937_ _01938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_05301_ _00926_ _00969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08020_ cpu.orig_IO_addr_buff\[0\] _03404_ _03303_ _03405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08840__A2 _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06851__A1 _02480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05232_ _00897_ _00902_ _00903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_112_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05163_ _00834_ _00835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_40_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09971_ _00230_ clknet_leaf_24_wb_clk_i net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_05094_ _00771_ _00786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06603__A1 _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08922_ _03057_ _04128_ _04129_ _04130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_0_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08853_ _01427_ _01273_ _04058_ _04062_ _04063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08784_ cpu.ROM_addr_buff\[10\] _03991_ _04000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05965__I0 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07804_ _03230_ _03195_ _03190_ _03232_ _03233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05996_ _01432_ _01657_ _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04947_ net71 _00647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_07735_ _03157_ _03176_ _03177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_84_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09405_ _02312_ _02313_ _04550_ _04586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_04878_ _00571_ _00580_ _00581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07666_ cpu.uart.div_counter\[12\] _03115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07597_ cpu.spi.div_counter\[5\] _03065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06617_ _02271_ _01799_ _02268_ _02272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09336_ _01916_ _04482_ _02338_ _04529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06548_ _02204_ _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_75_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05893__A2 _01107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09267_ _02204_ _01537_ _04463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08218_ _03552_ _03562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06479_ _02133_ _02135_ _02136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_105_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09198_ _04257_ _04382_ _04396_ _04260_ _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_95_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08149_ _03497_ _01512_ _03492_ cpu.toggle_ctr\[9\] _03498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_10111_ _00370_ clknet_leaf_4_wb_clk_i cpu.timer_top\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output67_I net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10042_ _00301_ clknet_leaf_52_wb_clk_i cpu.orig_IO_addr_buff\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09444__C _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04908__A1 cpu.base_address\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_10_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05008__S1 _00704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09075__A2 _00636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_85_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_85_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_109_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_14_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_14_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_53_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08590__I _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05850_ _01264_ _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__07010__A1 cpu.toggle_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07520_ _03001_ _03002_ _01893_ _03003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_89_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05572__A1 _01231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05781_ _00844_ _00840_ _01284_ _01446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_99_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07451_ cpu.timer_div\[7\] _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_92_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06402_ _01947_ _01295_ _02059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06285__I _01941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07382_ _01939_ _02873_ _02876_ _02877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_84_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09121_ _04299_ _04318_ _04322_ _04323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06333_ _00727_ _01990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_29_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06264_ _01911_ _01916_ _01920_ _01921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_09052_ _04116_ _04256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08003_ _03385_ _03388_ _03391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05215_ _00855_ _00874_ _00885_ _00886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06195_ _00880_ _01853_ _01854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_53_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08577__A1 _03801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05146_ cpu.PORTA_DDR\[6\] net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_12_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09954_ _00213_ clknet_leaf_37_wb_clk_i cpu.spi.div_counter\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05077_ _00752_ _00770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_90_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08905_ _04078_ _04113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09885_ _00144_ clknet_leaf_88_wb_clk_i cpu.regs\[7\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08836_ _01151_ _01969_ _04046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07001__A1 _00986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08767_ cpu.last_addr\[6\] _03981_ _03987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05979_ _01638_ _01639_ _01640_ _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05563__A1 cpu.timer_capture\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07718_ cpu.spi.counter\[1\] _03162_ _03164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08698_ _03932_ _00444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07649_ cpu.uart.receive_buff\[3\] _03102_ _03103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_36_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09319_ cpu.ROM_addr_buff\[6\] _04504_ _04512_ _04513_ _04514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_8_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06815__A1 cpu.uart.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08568__A1 cpu.uart.divisor\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput42 net42 io_oeb[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput64 net64 io_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput75 net75 io_out[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06043__A2 _01121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput53 net53 io_oeb[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput97 net97 sram_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput86 net86 sram_addr[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10025_ _00284_ clknet_leaf_30_wb_clk_i cpu.uart.receive_div_counter\[7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05229__S1 _00899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08740__A1 _02366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09048__A2 _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06806__A1 _02441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06833__I _02465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05000_ _00000_ _00697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_50_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06951_ _02551_ _02567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09670_ _01356_ _01274_ _02465_ _01514_ _04795_ _04796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05902_ _00765_ _00932_ _01565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08621_ _03860_ _03871_ _00428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06882_ _01693_ _02508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05545__A1 _01209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05833_ _01496_ _01398_ _01222_ _01497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_6_Left_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08552_ _03812_ _03813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05764_ _01426_ _01428_ _01092_ _01429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08483_ _03739_ _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07503_ _02970_ cpu.timer\[7\] _02973_ _02986_ _02987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_07434_ cpu.spi.data_in_buff\[4\] _02921_ _02922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05695_ _01357_ _01359_ net51 _01360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_33_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07365_ _02053_ _02079_ _02861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09104_ _02212_ _02423_ _04306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_60_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07296_ _02783_ _02811_ _02814_ _00160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06316_ _01942_ _01960_ _01966_ _01971_ _01972_ _00872_ _01973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai33_4
XFILLER_0_32_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06247_ _01894_ net69 _01904_ _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_79_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09035_ _02216_ _03446_ _04132_ _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__07470__A1 cpu.timer_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07470__B2 cpu.timer_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08014__A3 _00622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06178_ cpu.timer_top\[7\] _01500_ _01247_ _01837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05129_ cpu.regs\[4\]\[7\] cpu.regs\[5\]\[7\] cpu.regs\[6\]\[7\] cpu.regs\[7\]\[7\]
+ _00816_ _00817_ _00819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09937_ _00196_ clknet_leaf_44_wb_clk_i net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_5_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05084__I0 cpu.regs\[12\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09868_ _00127_ clknet_leaf_96_wb_clk_i cpu.regs\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08819_ _00811_ _01692_ _04029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09799_ _00062_ clknet_leaf_10_wb_clk_i cpu.timer_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07289__A1 _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer8 _00925_ net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_79_Left_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10008_ _00267_ clknet_leaf_23_wb_clk_i cpu.uart.data_buff\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06828__I _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05480_ _01116_ _01145_ _01103_ _01146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_39_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07150_ cpu.regs\[12\]\[3\] _02720_ _02723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07081_ cpu.uart.receive_counter\[2\] _02673_ _02678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06101_ _01760_ _01761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06032_ _01692_ _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07983_ cpu.uart.receive_div_counter\[10\] _03366_ _03342_ _03374_ _03375_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09722_ _03439_ _02579_ _04838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06934_ _02394_ _01906_ _02411_ _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09653_ _02314_ _04552_ _04779_ _04780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06865_ _02493_ _00050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05816_ _01477_ _01478_ _01479_ _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08604_ _03837_ _03855_ _03856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09584_ cpu.PORTA_DDR\[4\] _04719_ _04720_ _04721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_118_Right_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06796_ _02435_ _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08535_ cpu.timer_div\[4\] _03799_ _03774_ _03800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05747_ cpu.timer_top\[1\] _01237_ _01411_ _01412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_65_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09680__A2 _00918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05678_ _01339_ _01341_ _01343_ _01333_ _01344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08466_ cpu.timer_capture\[9\] _03746_ _03727_ _03750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07417_ cpu.spi.dout\[0\] _02908_ _02675_ _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07691__B2 cpu.uart.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07691__A1 _02640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08397_ _03621_ _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07348_ cpu.regs\[3\]\[5\] _02843_ _02847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05129__S0 _00816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07279_ _02788_ _02797_ _02803_ _00154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05089__I cpu.multiplier.a\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10290_ _00548_ clknet_leaf_60_wb_clk_i net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09018_ _04179_ _04213_ _04222_ _04186_ _04223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_60_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05757__A1 cpu.toggle_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09452__C _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06182__A1 cpu.toggle_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08863__I _04071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07682__B2 _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09671__A2 _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08812__B _03395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_87_Left_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05748__A1 cpu.timer_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04980_ _00679_ _00680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_4_12_0_wb_clk_i clknet_0_wb_clk_i clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_06650_ _02297_ _02298_ _02302_ _02303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_79_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06558__I cpu.PC\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05601_ _01115_ _01267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_86_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06581_ _02236_ _02237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_96_Left_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05532_ _01197_ _01198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08320_ _03622_ _03630_ _03631_ _00367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_19_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05463_ _01128_ _01129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09662__A2 _01329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06020__S1 _00969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08251_ cpu.pwm_counter\[0\] _03584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07202_ _01814_ _02756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_27_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05394_ _01057_ _01059_ _01060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08182_ _03488_ cpu.toggle_top\[7\] cpu.toggle_top\[6\] _03530_ _03531_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_15_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06228__A2 _01390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07133_ _01869_ _02700_ _02709_ _00102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07064_ _02651_ cpu.uart.receive_div_counter\[15\] _02662_ cpu.uart.divisor\[3\]
+ _02663_ _02664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_76_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05987__A1 cpu.toggle_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05451__A3 _00611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06015_ _01658_ _01676_ _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07966_ _03352_ _03360_ _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input29_I sram_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06917_ _02459_ _02536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09705_ _01615_ _04820_ _04826_ _00557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07073__B _02623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07897_ _03307_ _03308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09636_ _01915_ _04763_ _04764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_69_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08153__A2 _01723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06848_ _02479_ _00047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06779_ _01101_ _02421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09567_ cpu.PORTB_DDR\[7\] _04704_ _04705_ _04709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08683__I _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09498_ _01068_ _02432_ _04663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08518_ cpu.spi.divisor\[7\] _03784_ _03788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08449_ _03729_ _03654_ _03730_ _03735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_37_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06219__A2 cpu.spi.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output97_I net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09169__A1 _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05978__A1 cpu.timer_capture\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08916__A1 _04106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10273_ _00531_ clknet_leaf_53_wb_clk_i cpu.PORTB_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_29_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_39_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_39_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_49_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08542__B _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08768__I _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07820_ cpu.uart.clr_hb _03246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09580__A1 _02529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07751_ cpu.uart.div_counter\[2\] cpu.uart.div_counter\[1\] cpu.uart.div_counter\[0\]
+ _03191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_19_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06702_ _02323_ _02355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_04963_ _00609_ _00663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07682_ _02632_ cpu.uart.div_counter\[13\] cpu.uart.div_counter\[6\] _02633_ _03130_
+ _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_04894_ _00591_ _00596_ _00597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09421_ _04600_ _04551_ _04601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06633_ _02264_ _02274_ _02276_ _02286_ _02287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09352_ _01908_ _04535_ _04542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06564_ _02210_ _02211_ _02220_ _02221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__05920__I cpu.uart.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05515_ _01176_ _01181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_75_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06449__A2 _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08303_ _03618_ _03620_ _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09283_ _02369_ _04478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_82_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06495_ _02147_ _02151_ _02152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08008__I _02929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08234_ _03562_ _03572_ _03573_ _00339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05446_ _01109_ _01111_ _01112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05377_ _01042_ _01043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08165_ cpu.toggle_ctr\[5\] _03514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07116_ _02698_ _02700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_113_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08096_ _02856_ _03459_ _03460_ _00314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07047_ cpu.uart.receive_div_counter\[5\] _01695_ _02638_ cpu.uart.receive_div_counter\[2\]
+ _02646_ _02647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_2_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08678__I _00648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08998_ _04167_ _04178_ _04204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06385__A1 _00854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07949_ _02662_ _03340_ _03347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09619_ _02310_ _04748_ _04735_ _04749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08346__C _03648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08834__B1 _04043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06160__I1 cpu.PORTA_DDR\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09177__C _04321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05277__I _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10325_ net49 net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10256_ _00514_ clknet_leaf_46_wb_clk_i net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__08588__I _03839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09562__A1 _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10187_ _00445_ clknet_leaf_67_wb_clk_i cpu.ROM_addr_buff\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06128__A1 cpu.toggle_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_89_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07876__A1 _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06280_ _01924_ _01937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05300_ _00890_ _00968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05231_ _00900_ _00901_ _00832_ _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05162_ _00004_ _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_09970_ _00229_ clknet_leaf_36_wb_clk_i cpu.uart.dout\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05093_ _00770_ _00785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_110_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08921_ _03439_ _04072_ _04129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09553__A1 _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08852_ _01266_ _02416_ _04061_ _04062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07803_ _03230_ _03231_ _03232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08783_ cpu.last_addr\[10\] _03999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05995_ _01619_ _01155_ _01656_ _01657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04946_ _00634_ _00646_ _00010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07734_ _00599_ _01895_ _03176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_84_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07665_ net68 _03114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09404_ _04560_ _02296_ _04585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04877_ _00575_ _00579_ _00580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__04975__B _00674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06616_ _00815_ _02271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_109_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09122__I _00693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07596_ _03064_ _00210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05342__A2 _01007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09335_ _04528_ _00485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06547_ cpu.PC\[12\] _02204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_51_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09266_ _00671_ _01160_ _04460_ _04461_ _04462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_63_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06478_ _02114_ _02117_ _02134_ _02135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05429_ _00663_ _00610_ _01094_ _01095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08217_ _03553_ _03561_ _00334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09197_ _02882_ _04258_ _04396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08148_ cpu.toggle_ctr\[10\] _03497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08079_ _03446_ _03434_ _03448_ _00309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_31_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10110_ _00369_ clknet_leaf_21_wb_clk_i cpu.timer_div_counter\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09544__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10041_ _00300_ clknet_leaf_50_wb_clk_i cpu.orig_IO_addr_buff\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_59_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_6_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08092__B _03457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_54_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_54_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_21_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_60_Left_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10239_ _00497_ clknet_leaf_62_wb_clk_i cpu.spi_clkdiv vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05780_ _01440_ _01444_ _01445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_107_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07450_ cpu.timer_div_counter\[5\] _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_91_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06401_ _01940_ _02057_ _02058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07381_ _02573_ _02874_ _02875_ _02876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_09120_ _04267_ _04303_ _04320_ _04235_ _04321_ _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_45_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06332_ _01973_ _01985_ _01988_ _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_45_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09051_ _04249_ _04252_ _04253_ _04254_ _04255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_45_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08002_ cpu.uart.receive_div_counter\[14\] _03389_ _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06263_ _01918_ _01919_ _01920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06194_ _01326_ _01297_ _01853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05214_ _00882_ _00884_ _00885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05145_ cpu.PORTB_DDR\[6\] net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_13_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09953_ _00212_ clknet_leaf_47_wb_clk_i cpu.spi.div_counter\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05076_ cpu.regs\[2\]\[4\] _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08904_ _03438_ _01151_ _04111_ _04112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09884_ _00143_ clknet_leaf_87_wb_clk_i cpu.regs\[7\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_90_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08835_ _04042_ _04045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08766_ _03984_ _03985_ _03986_ _00458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_56_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input11_I io_in[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07717_ _03160_ _03013_ _03163_ _00231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05978_ cpu.timer_capture\[4\] _01401_ _01227_ _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06760__A1 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08697_ _03931_ cpu.ROM_addr_buff\[5\] _03921_ _03932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_95_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04929_ _00624_ _00625_ _00630_ _00011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09280__C _04007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07648_ _03093_ _03102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_67_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07579_ _03048_ _01884_ _03050_ _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_TAPCELL_ROW_64_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06512__B2 _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09318_ _03980_ cpu.ROM_addr_buff\[4\] _04486_ _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_94_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09249_ _02205_ _04258_ _04446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06579__A1 _00784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput43 net43 io_oeb[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput65 net65 io_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput76 net76 io_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput54 net54 io_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09517__A1 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_8_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput87 net87 sram_addr[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10024_ _00283_ clknet_leaf_30_wb_clk_i cpu.uart.receive_div_counter\[6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_101_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_101_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07303__I0 _02818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08256__A1 _03585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09365__C _02359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09508__A1 _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06950_ _01678_ _02554_ _02565_ _02566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input3_I io_in[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06881_ _02507_ _00052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05901_ _00932_ _01451_ _01563_ _01453_ _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05793__A2 _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05832_ cpu.timer_div\[2\] _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08620_ _01064_ _03861_ _03869_ _03870_ _03871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08551_ _03807_ _03809_ _03811_ _00626_ _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_68_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05763_ _01427_ _01138_ _01428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05694_ _01358_ _01359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08482_ cpu.timer\[12\] _03761_ _03762_ _03763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07502_ cpu.timer_top\[6\] _02972_ _02974_ cpu.timer_top\[5\] _02985_ _02986_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_07433_ _01901_ _02921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_77_Right_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_61_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09103_ cpu.PC\[6\] _01034_ _04304_ _04305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07364_ _02056_ _02078_ _02860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07295_ cpu.regs\[5\]\[1\] _02812_ _02814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06315_ _01964_ _01965_ _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_32_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06246_ _01897_ _01902_ _01903_ _01904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__08016__I _03400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09034_ _02570_ _04073_ _04238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_107_Left_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_79_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05481__A1 _01115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06177_ cpu.timer_capture\[15\] _01234_ _01835_ _01237_ _01836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05128_ cpu.regs\[0\]\[7\] _00815_ cpu.regs\[2\]\[7\] cpu.regs\[3\]\[7\] _00816_
+ _00817_ _00818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09936_ _00195_ clknet_leaf_57_wb_clk_i cpu.needs_timer_interrupt vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_86_Right_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_5_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05059_ _00717_ _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05084__I1 cpu.regs\[13\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06981__A1 _00798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09867_ _00126_ clknet_leaf_108_wb_clk_i cpu.regs\[10\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_116_Left_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08818_ _01334_ _01459_ _04028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09798_ _00061_ clknet_leaf_10_wb_clk_i cpu.timer_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08749_ cpu.ROM_addr_buff\[1\] _03970_ _03974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07289__A2 _02777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08486__A1 _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_95_Right_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08789__A2 _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer9 _02164_ net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05472__A1 _00655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09738__A1 _00728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06972__A1 _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10007_ _00266_ clknet_leaf_23_wb_clk_i cpu.uart.data_buff\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08529__C _03648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08477__A1 cpu.timer_capture\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07005__I _02456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07080_ _01903_ _02677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06100_ _01759_ _01760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06031_ _01691_ _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09729__A1 _01466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08401__A1 cpu.timer_capture\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07982_ _03372_ _03373_ _03374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09721_ _04835_ _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06963__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06933_ _02203_ _01932_ _02549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09652_ _04560_ _04549_ _04544_ _04779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06864_ cpu.timer_capture\[3\] _02471_ _02492_ _02484_ _02493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05815_ net23 _01199_ _01052_ _01479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06795_ _02434_ _02435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08603_ _03854_ _03844_ _03855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09583_ _02378_ _04720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08534_ _03789_ _03799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05746_ _01410_ _01411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05677_ _01342_ _01343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08465_ _02960_ _03742_ _03748_ _03749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07416_ _01890_ _02908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08396_ _03691_ _00383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07347_ _02846_ _00179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05129__S1 _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08640__A1 _02419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09017_ _04217_ _04220_ _04221_ _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07278_ cpu.regs\[6\]\[3\] _02801_ _02803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07585__I _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06229_ _01882_ _01883_ _01886_ _01887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__05057__I1 _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09919_ _00178_ clknet_leaf_94_wb_clk_i cpu.regs\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05509__A2 _01065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output42_I net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08459__A1 _02425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05445__A1 _01110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08147__B1 cpu.toggle_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06839__I _02470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05600_ cpu.C _01266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06580_ _01619_ _01043_ _01118_ _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_05531_ _01014_ _01015_ _01197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_46_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05462_ _01127_ _01128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08250_ _03494_ _03580_ _03553_ _00345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05684__A1 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08181_ cpu.toggle_ctr\[6\] _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07201_ _02725_ _02747_ _02755_ _00124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05393_ _00653_ _01058_ _01059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_9_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_9_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07132_ cpu.regs\[13\]\[7\] _02703_ _02709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05436__A1 _00618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08622__B2 _00919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07063_ cpu.uart.divisor\[11\] cpu.uart.receive_div_counter\[11\] _02663_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_76_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06014_ net30 _01527_ _01463_ _01675_ _01104_ _01676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_11_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07965_ _03359_ _03356_ _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06916_ _02532_ _02533_ _02535_ _02531_ _00059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09704_ cpu.regs\[9\]\[3\] _04824_ _04826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07896_ _03306_ net15 _03307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09635_ _02321_ _02326_ _02397_ _01911_ _04763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_87_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06847_ cpu.timer_capture\[0\] _02471_ _02477_ _02478_ _02479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06778_ _02382_ _02415_ _02420_ _00036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09566_ _02538_ _04703_ _04708_ _00536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09497_ _04660_ _04662_ _03043_ _00513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05729_ _01389_ _01391_ _01393_ _01394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09102__A2 _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08517_ _02538_ _03783_ _03787_ _00408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07113__A1 _01114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08448_ _03734_ _00392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_41_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08379_ _03653_ _03674_ _03676_ _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10272_ _00530_ clknet_leaf_53_wb_clk_i cpu.PORTB_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA_clkbuf_leaf_79_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_79_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_79_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05902__A2 _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07104__A1 _01114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08095__B _03457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05666__A1 _01329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05004__S _00002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_71_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07591__A1 _03057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07750_ _03180_ _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04962_ _00661_ _00662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06701_ cpu.ROM_addr_buff\[11\] _02335_ _02330_ _02354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07681_ _02628_ _03129_ cpu.uart.div_counter\[5\] _01695_ _03130_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_04893_ _00595_ _00596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07343__A1 _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09420_ _02295_ _04600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06632_ _02284_ _02285_ _02286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09351_ _03965_ _04483_ _04541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06563_ _02212_ _02213_ _02219_ _02220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_59_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09282_ _04457_ _04477_ _04431_ _00483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05514_ _01179_ _01180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08302_ cpu.pwm_top\[7\] _03613_ _03619_ _03620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08233_ cpu.toggle_ctr\[9\] _03571_ _03573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06494_ _02121_ _02149_ _02150_ _02151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_90_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05445_ _01110_ _01104_ _01111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09399__A2 _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05376_ _01040_ _01041_ _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08164_ cpu.toggle_ctr\[6\] _03511_ _03512_ cpu.toggle_ctr\[5\] _03513_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_7_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08095_ cpu.orig_PC\[8\] _03454_ _03457_ _03460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07115_ _02698_ _02699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08452__C _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07046_ _02639_ _02441_ _01183_ cpu.uart.receive_div_counter\[0\] _02645_ _02646_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_30_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_113_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06909__A1 cpu.timer_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08997_ _04176_ _04178_ _04201_ _04202_ _04203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07948_ _03335_ _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07879_ _03291_ _03293_ _03294_ _00263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09618_ _04746_ _04747_ _04742_ _04748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09549_ _04674_ _04698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07531__C _02404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05896__A1 _00763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05648__A1 _00910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08834__A1 _01116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08834__B2 _01151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10255_ _00513_ clknet_leaf_59_wb_clk_i net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10186_ _00444_ clknet_leaf_66_wb_clk_i cpu.ROM_addr_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_109_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05293__I _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07441__C _00694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08825__A1 _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05639__A1 _01303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07013__I _02610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06852__I _00626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05230_ cpu.regs\[8\]\[2\] cpu.regs\[9\]\[2\] cpu.regs\[10\]\[2\] cpu.regs\[11\]\[2\]
+ _00898_ _00899_ _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_05161_ _00832_ _00833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06064__A1 _01694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05092_ cpu.regs\[2\]\[5\] _00784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_40_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08779__I _03966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08920_ _00644_ _00689_ _02428_ _04127_ _04128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09002__A1 _02389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05811__A1 net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08851_ _01356_ _01514_ _01274_ _01761_ _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07802_ _03115_ _03227_ _03231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08782_ _03984_ _03997_ _03998_ _00462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05994_ _00958_ _01521_ _01653_ _01654_ _01655_ _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_07733_ _03160_ _03174_ _03175_ _00235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_04945_ _00629_ _00641_ _00644_ _00645_ _00646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_46_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07664_ _03111_ _03095_ _03112_ _03113_ _00229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_04876_ net129 _00578_ _00579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09403_ _02345_ _04584_ _04431_ _00497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_84_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08447__C _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06615_ _02130_ _01691_ _02269_ _02270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07595_ cpu.spi.div_counter\[4\] _03058_ _03063_ _02506_ _03064_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_62_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09334_ _01912_ _04481_ _04526_ _04527_ _04528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08019__I _03403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06546_ _01938_ _02203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_23_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09265_ _02254_ _04189_ _04084_ _04461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06477_ _01968_ _02116_ _02134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05428_ _00678_ _00672_ _01094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09196_ _04254_ _04393_ _04394_ _04395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_62_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08216_ _03515_ _03559_ _03561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05359_ _01024_ _01025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08147_ _03494_ cpu.toggle_top\[15\] cpu.toggle_top\[14\] _03495_ _03496_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_113_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08078_ cpu.orig_PC\[3\] _03443_ _03447_ _03448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07029_ cpu.uart.receive_div_counter\[9\] _02629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_10040_ _00299_ clknet_leaf_51_wb_clk_i cpu.orig_IO_addr_buff\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_59_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_104_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08373__B _03615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06046__A1 cpu.uart.dout\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05288__I _00955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08599__I _03850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10307_ _00565_ clknet_leaf_84_wb_clk_i cpu.multiplier.a\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_94_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_94_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10238_ _00496_ clknet_leaf_60_wb_clk_i cpu.startup_cycle\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_23_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_23_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10169_ _00427_ clknet_leaf_15_wb_clk_i cpu.IO_addr_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06400_ _00946_ _01993_ _01995_ _01731_ _02057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_57_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07380_ _02104_ _02126_ _02875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06331_ _01986_ _01959_ _01972_ _01987_ _01988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_17_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06262_ cpu.mem_cycle\[2\] _01919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09050_ _04147_ _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08001_ _03333_ _03388_ _03389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05213_ _00883_ _00884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06193_ net33 _01852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_13_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06037__A1 net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05144_ cpu.PORTA_DDR\[5\] net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_09952_ _00211_ clknet_leaf_46_wb_clk_i cpu.spi.div_counter\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05075_ _00767_ _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_110_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08903_ cpu.PC\[0\] cpu.br_rel_dest\[0\] _04111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_90_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09883_ _00142_ clknet_leaf_111_wb_clk_i cpu.regs\[8\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_90_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08834_ _01116_ _04042_ _04043_ _01151_ _04044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08765_ cpu.ROM_addr_buff\[5\] _03976_ _03986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_56_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07716_ _03009_ _03162_ _03163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05977_ cpu.timer_div\[4\] _01397_ _01221_ _01639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_95_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08696_ _02214_ _03917_ _03930_ _03931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04928_ _00628_ cpu.instr_cycle\[3\] _00629_ _00630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_0_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07647_ _03093_ _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_67_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07578_ _01902_ _03050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_64_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09317_ _04505_ _04506_ _04508_ _04511_ _04512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_06529_ _02009_ _02186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_63_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06276__A1 _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09248_ _04249_ _04443_ _04444_ _04366_ _04445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09179_ _04355_ _04378_ _04324_ _00479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_114_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06579__A2 _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput66 net66 io_out[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput55 net55 io_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07537__B _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput44 net44 io_oeb[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput77 net77 io_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput88 net88 sram_addr[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10023_ _00282_ clknet_leaf_32_wb_clk_i cpu.uart.receive_div_counter\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__06200__A1 _00826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04915__I net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05746__I _01410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06880_ cpu.timer_capture\[5\] _02494_ _02505_ _02506_ _02507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05900_ _00764_ _00931_ _01563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05831_ _01494_ _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05625__S0 _01285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08550_ _03810_ _03811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05762_ cpu.Z _01427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05693_ _01191_ _01358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07501_ _01716_ cpu.timer\[5\] _02498_ _01620_ _02984_ _02985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08481_ _02495_ _03751_ _03762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07432_ _02919_ _02920_ _02915_ _00190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_85_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09102_ _03452_ _01058_ _04279_ _04304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_57_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07363_ _01939_ _02858_ _02859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07294_ _02776_ _02811_ _02813_ _00159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06314_ _01969_ _01970_ _01971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06245_ _00626_ _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09033_ _04211_ _04237_ _04210_ _00474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_115_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06176_ _01832_ _01833_ _01834_ _01835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05127_ _00786_ _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09935_ _00194_ clknet_leaf_37_wb_clk_i cpu.spi.dout\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08032__I _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05058_ _00730_ _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__05084__I2 cpu.regs\[14\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09866_ _00125_ clknet_leaf_111_wb_clk_i cpu.regs\[10\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08817_ _01747_ _01811_ _01865_ _04026_ _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06733__A2 _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09797_ _00060_ clknet_leaf_10_wb_clk_i cpu.timer_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08748_ cpu.last_addr\[1\] _03967_ _03973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08679_ _03916_ _03917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_101_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06972__A2 _02569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10006_ _00265_ clknet_leaf_23_wb_clk_i cpu.uart.data_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08098__B _03457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08826__B _04035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09501__I _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08117__I _03473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06860__I _00933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06030_ _01685_ _01690_ _01691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_10_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07981_ _03365_ _03367_ cpu.uart.receive_div_counter\[10\] _03373_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09720_ _04836_ _00562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06932_ _02547_ _02548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09651_ _02351_ _04777_ _04778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06715__A2 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06863_ _02489_ _02473_ _02474_ _02491_ _02492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05814_ net61 _01195_ _01188_ _01478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_89_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08602_ _03839_ _03854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06794_ _01184_ _02433_ _02434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09582_ _04710_ _04719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05745_ _01213_ _01080_ _01410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08533_ _02453_ _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06100__I _01759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05676_ _01336_ _01157_ _01328_ _01342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_46_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08464_ _02480_ _03743_ _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07415_ _01890_ _02907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_92_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08395_ cpu.timer_capture\[5\] _03678_ _03689_ _03690_ _03691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_18_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07346_ _02818_ cpu.regs\[3\]\[4\] _02838_ _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_116_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09016_ _04217_ _04220_ _04110_ _04221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07277_ _02785_ _02797_ _02802_ _00153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06228_ cpu.spi.div_counter\[1\] _01390_ cpu.spi.divisor\[4\] _01875_ _01885_ _01886_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__06770__I _02413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06159_ cpu.uart.divisor\[7\] _01818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05057__I2 _00748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09918_ _00177_ clknet_leaf_93_wb_clk_i cpu.regs\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_69_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07815__B _03242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09849_ _00108_ clknet_leaf_106_wb_clk_i cpu.regs\[12\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output35_I net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_14_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08395__A1 cpu.timer_capture\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07016__I _02456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07370__A2 _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05530_ cpu.PORTB_DDR\[0\] _01021_ _01195_ _01196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05461_ _00605_ _01002_ _01117_ _01127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_74_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05392_ _00602_ _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07200_ cpu.regs\[10\]\[5\] _02750_ _02755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08180_ _03526_ cpu.toggle_top\[1\] cpu.toggle_top\[0\] _03528_ _03529_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_82_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07131_ _02708_ _00101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08622__A2 _03864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07062_ cpu.uart.receive_div_counter\[3\] _02662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_76_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05436__A2 _00583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06013_ _01454_ _01659_ _01674_ _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_clkbuf_leaf_103_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08925__A3 cpu.PC\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07964_ cpu.uart.receive_div_counter\[7\] _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08138__A1 _02467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07895_ cpu.uart.receiving _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06915_ cpu.timer_top\[4\] _02534_ _02535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09703_ _01551_ _04820_ _04825_ _00556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09634_ _02302_ _04761_ _04551_ _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06846_ _01903_ _02478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_69_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_87_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06777_ _02419_ _02414_ _00685_ _02420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09565_ cpu.PORTB_DDR\[6\] _04704_ _04705_ _04708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09496_ net89 _04661_ _00649_ _04662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05728_ _01392_ _01393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_65_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08516_ cpu.spi.divisor\[6\] _03784_ _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07113__A2 _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05659_ _01324_ _01325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08447_ cpu.timer_capture\[14\] _03714_ _03733_ _03722_ _03734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_80_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08378_ cpu.timer_capture\[3\] _03660_ _03675_ _03676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07329_ _02821_ cpu.regs\[4\]\[6\] _02825_ _02835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_33_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06624__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10271_ _00529_ clknet_leaf_42_wb_clk_i net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_14_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05038__S1 _00731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07104__A2 _02684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08852__A2 _02416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06863__A1 _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_71_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04961_ _00659_ _00660_ _00661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06700_ _02334_ _02353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07680_ cpu.uart.div_counter\[9\] _03129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_04892_ _00594_ _00595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08540__A1 _03801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06631_ _02130_ _02069_ _02070_ _01761_ _02285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_09350_ _04540_ _00488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_87_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09096__A2 _04273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06562_ _02214_ _02216_ _02218_ _02219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09281_ _04206_ _04473_ _04476_ _04477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05513_ _01009_ _00998_ _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08301_ _02466_ _03602_ _03619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08843__A2 _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06854__A1 cpu.timer_capture\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05657__A2 _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08232_ cpu.toggle_ctr\[9\] _03571_ _03572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06493_ _02148_ _02118_ _02150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_117_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05444_ _00652_ _01110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_62_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05375_ _00652_ cpu.br_rel_dest\[6\] _01041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_08163_ cpu.toggle_top\[5\] _03512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08094_ _03403_ _03459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_70_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07114_ _02697_ _02698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_113_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07045_ _02640_ _02641_ cpu.uart.receive_div_counter\[8\] _02642_ _02644_ _02645_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__06082__A2 _00980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08996_ _04161_ _04202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07947_ _03308_ _03345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05593__A1 _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07878_ cpu.uart.data_buff\[6\] _03288_ _03289_ _03294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09617_ cpu.ROM_addr_buff\[5\] _02355_ _02356_ cpu.ROM_addr_buff\[9\] cpu.ROM_addr_buff\[13\]
+ _02340_ _04747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_06829_ _02462_ _02463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09548_ _04695_ _04697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09087__A2 _03854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08834__A2 _04042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09479_ cpu.pwm_top\[7\] cpu.pwm_counter\[7\] _04646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06845__A1 _02425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08598__A1 _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06073__A2 _01733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09011__A2 _01107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10254_ _00512_ clknet_leaf_102_wb_clk_i net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10185_ _00443_ clknet_leaf_72_wb_clk_i cpu.ROM_addr_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07022__A1 _02467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09078__A2 _02421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06836__A1 _02467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05195__S0 _00858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05160_ _00831_ _00832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_110_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05091_ _00782_ _00783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05811__A2 _01190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08850_ _01278_ _04012_ _04058_ _04059_ _04060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07801_ cpu.uart.div_counter\[13\] _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05484__I _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08781_ cpu.ROM_addr_buff\[9\] _03988_ _03998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05993_ _01044_ _01304_ _01655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_46_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07732_ _03007_ _01898_ _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04944_ _00627_ _00645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08513__A1 _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07663_ _03055_ _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04875_ _00577_ _00578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_84_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09402_ cpu.spi_clkdiv _04583_ _04584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_84_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06614_ _01759_ _02069_ _02130_ _02269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09333_ _00627_ _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07594_ _01875_ _03038_ _02921_ _03050_ _03062_ _03063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_48_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06545_ _02178_ _02200_ _02202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_90_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06827__A1 _02460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09264_ _03849_ _04458_ _04460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06476_ _02130_ _02132_ _02133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09195_ _04249_ _04382_ _04394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05427_ _00583_ _01093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08215_ _03555_ _03559_ _03560_ _00333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08146_ cpu.toggle_ctr\[14\] _03495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09241__A2 _03863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05358_ _00605_ _01007_ _01024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08077_ _03410_ _03447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05289_ _00957_ _00958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_07028_ cpu.uart.divisor\[9\] _02628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08979_ _04181_ _04182_ _04184_ _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_59_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05110__S0 _00799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05869__A2 _00916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06046__A2 _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10306_ _00564_ clknet_leaf_85_wb_clk_i cpu.multiplier.a\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_115_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10237_ _00495_ clknet_leaf_44_wb_clk_i cpu.startup_cycle\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08743__A1 _02366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10168_ _00426_ clknet_leaf_36_wb_clk_i cpu.uart.divisor\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05101__S0 _00770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10099_ _00358_ clknet_leaf_11_wb_clk_i cpu.pwm_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_63_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_63_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_89_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06330_ _01977_ _01978_ _01982_ _01983_ _01987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__05168__S0 _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06261_ _01917_ _01918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_96_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07482__A1 cpu.timer_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08000_ cpu.uart.receive_div_counter\[14\] _03385_ _03330_ _03388_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05212_ _00853_ _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07482__B2 cpu.timer_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06192_ _01033_ _01431_ _01306_ _01851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05143_ cpu.PORTB_DDR\[5\] net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_40_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09951_ _00210_ clknet_leaf_37_wb_clk_i cpu.spi.div_counter\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05074_ cpu.multiplier.a\[4\] _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08902_ _04081_ _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05796__A1 _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08734__A1 _02254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09882_ _00141_ clknet_leaf_113_wb_clk_i cpu.regs\[8\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_90_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08833_ _01969_ _04043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08764_ cpu.last_addr\[5\] _03981_ _03985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05976_ _01633_ _01635_ _01637_ _01638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07715_ _01897_ _03161_ _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_04927_ _00622_ _00629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08695_ _03926_ _00784_ _03930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07646_ cpu.uart.dout\[3\] _03100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_0_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07577_ _03046_ _03045_ _03048_ _03049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_64_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09316_ net130 _03964_ _04509_ _04510_ _04511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_06528_ _02161_ _02183_ _02184_ _02185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09247_ _04138_ _04436_ _04444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06459_ _02065_ _02115_ _02116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_105_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09178_ _04299_ _04373_ _04377_ _04378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08129_ _03473_ _03482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput34 net34 io_oeb[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput67 net67 io_out[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput56 net56 io_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput45 net45 io_oeb[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput78 net78 io_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput89 net89 sram_gwe vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10022_ _00281_ clknet_leaf_33_wb_clk_i cpu.uart.receive_div_counter\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05539__A1 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_113_Right_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07779__I _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06267__A2 _01434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_110_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_110_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_41_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09610__C1 cpu.ROM_addr_buff\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08964__A1 _02389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_9_0_wb_clk_i clknet_0_wb_clk_i clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08716__A1 _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06990__A3 _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08559__B _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05830_ cpu.spi.dout\[2\] _01177_ _01397_ _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_27_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05625__S1 _01286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05761_ _01356_ _01283_ _01425_ _01299_ _01426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_07500_ cpu.timer_top\[3\] _02975_ _02976_ cpu.timer_top\[4\] _02983_ _02984_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_89_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05692_ _01047_ _01357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05002__I0 cpu.regs\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08480_ _03741_ _03761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07431_ cpu.spi.data_in_buff\[3\] _02908_ _02920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05702__A1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07362_ _02856_ _02857_ _02858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_61_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09101_ _04302_ _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06313_ _01952_ _00883_ _01970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07293_ cpu.regs\[5\]\[0\] _02812_ _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06244_ _01898_ _01901_ _01902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09032_ _04175_ _04231_ _04236_ _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06175_ cpu.timer_capture\[7\] _01402_ _01228_ _01834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05126_ _00785_ _00816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_40_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09934_ _00193_ clknet_leaf_47_wb_clk_i cpu.spi.dout\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05084__I3 cpu.regs\[15\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05057_ cpu.regs\[0\]\[3\] _00747_ _00748_ cpu.regs\[3\]\[3\] _00749_ _00750_ _00751_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_clkbuf_leaf_59_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08707__A1 _02597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09865_ _00124_ clknet_leaf_108_wb_clk_i cpu.regs\[10\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08816_ _01547_ _01570_ _01675_ _04025_ _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_09796_ _00059_ clknet_leaf_10_wb_clk_i cpu.timer_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05959_ net2 _01621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08747_ _03159_ _03972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05941__A1 cpu.toggle_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08678_ _00648_ _03916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08983__I _04150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07629_ _02364_ _03088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_95_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09683__A2 _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05472__A3 _01118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09199__A1 _00913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_98_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08946__A1 _04150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_2_Left_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_39_Left_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10005_ _00264_ clknet_leaf_22_wb_clk_i cpu.uart.data_buff\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05932__A1 cpu.timer_capture\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_48_Left_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_57_Left_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_10_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07980_ cpu.uart.receive_div_counter\[10\] _03365_ _03367_ _03372_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__06412__A2 _00798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06931_ _02543_ _02546_ _02547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09650_ _02398_ _04776_ _02353_ _04777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08601_ _03838_ _03846_ _03852_ _03853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_66_Left_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06176__A1 _01832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06862_ _02490_ _02475_ _02491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05223__I0 cpu.regs\[4\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05923__A1 _00615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05813_ _01474_ _01475_ _01476_ _01477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06793_ _02432_ _02433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09581_ _04710_ _04718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08532_ _03796_ _03793_ _03797_ _00413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05744_ _01404_ _01406_ _01408_ _01409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07676__A1 cpu.uart.divisor\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09665__A2 _01990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08463_ _03740_ _03745_ _03747_ _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07414_ cpu.spi.data_in_buff\[0\] _02906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05675_ _01340_ _01341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_46_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08394_ _02483_ _03690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07345_ _01615_ _02839_ _02845_ _00178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_75_Left_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07276_ cpu.regs\[6\]\[2\] _02801_ _02802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06227_ _01884_ cpu.spi.divisor\[0\] _01390_ cpu.spi.div_counter\[1\] _01885_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09015_ _04218_ _04219_ _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09139__I _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07368__B _02573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08043__I _03410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06158_ _01817_ _00019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06089_ _01307_ _01749_ _01750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__06403__A2 _01691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05109_ _00771_ _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09917_ _00176_ clknet_leaf_93_wb_clk_i cpu.regs\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06167__A1 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07203__I1 cpu.regs\[10\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09848_ _00107_ clknet_leaf_115_wb_clk_i cpu.regs\[12\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05914__A1 net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09779_ _00042_ clknet_leaf_24_wb_clk_i cpu.uart.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_96_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08662__B _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09719__I0 _04042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04956__A2 _00655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09512__I _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05460_ _01125_ _01126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_15_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08128__I _03473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05391_ _00584_ _00657_ _01057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_55_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07130_ _01816_ cpu.regs\[13\]\[6\] _02698_ _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07130__I0 _01816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07061_ _02648_ _02658_ _02659_ _02633_ _02660_ _02661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_76_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06012_ _01664_ _01666_ _01673_ _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07963_ _03357_ _03358_ _00283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07894_ _03305_ _00267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06914_ _02519_ _02534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09702_ cpu.regs\[9\]\[2\] _04824_ _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09633_ _02308_ _04758_ _02311_ _04761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06845_ _02425_ _02473_ _02474_ _02476_ _02477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_97_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09564_ _02536_ _04703_ _04707_ _00535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06776_ _02418_ _02419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08515_ _02536_ _03783_ _03786_ _00407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09495_ _00682_ _03810_ _04661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05727_ _01067_ _01128_ _01392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_93_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05658_ _00908_ _01324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06321__A1 _01941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08446_ _03681_ _03731_ _03732_ _03662_ _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_108_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_83_Left_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08377_ _03608_ _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07328_ _02791_ _02827_ _02834_ _00172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05589_ cpu.pwm_top\[0\] _01252_ _01254_ _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08074__A1 _03442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07259_ _02790_ _00147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06624__A2 _02229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10270_ _00528_ clknet_leaf_42_wb_clk_i net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_61_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09574__A1 _02518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_92_Left_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08501__I _03776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05346__B _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07888__A1 _02513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08301__A2 _03602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_88_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_88_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_24_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_17_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_17_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_51_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06615__A2 _01691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09565__A1 cpu.PORTB_DDR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04960_ cpu.uart.busy cpu.spi.busy _00640_ _00660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__07179__I0 _01816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04891_ _00592_ _00593_ _00594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06630_ _02267_ _02273_ _02272_ _02284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05770__I _01434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06866__I _02470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06561_ _02217_ cpu.PC\[2\] cpu.PC\[1\] _02218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_59_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09280_ _04374_ _04459_ _04475_ _04404_ _04007_ _04476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05512_ cpu.spi.divisor\[0\] _01178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08300_ _02379_ _03618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_47_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06492_ _02148_ _02118_ _02149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05443_ _01108_ _01092_ _01097_ _00911_ _01109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_08231_ _03555_ _03570_ _03571_ _00338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09398__B _00693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06815__B _02391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05374_ _00618_ _00571_ _01039_ _01040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_08162_ cpu.toggle_top\[6\] _03511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08093_ _02597_ _03449_ _03458_ _00313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07113_ _01114_ _02546_ _02697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07044_ cpu.uart.divisor\[10\] _02641_ _02643_ cpu.uart.divisor\[0\] _02644_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_3_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09556__A1 cpu.PORTB_DDR\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05290__A1 _00911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05010__I _00002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08995_ _04187_ _04196_ _04200_ _04201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07946_ _03327_ _03344_ _00280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input27_I sram_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05593__A2 _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07877_ cpu.uart.data_buff\[5\] _03282_ _03292_ _03293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09616_ cpu.ROM_addr_buff\[1\] _04738_ _02327_ _04746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_92_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06828_ _01693_ _02462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09547_ _04695_ _04696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06759_ _02403_ _02406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09478_ cpu.pwm_top\[4\] cpu.pwm_counter\[4\] _04645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_108_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_11_0_wb_clk_i clknet_0_wb_clk_i clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_53_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08429_ _03718_ _00389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output95_I net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10253_ _00511_ clknet_leaf_65_wb_clk_i net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10184_ _00442_ clknet_leaf_64_wb_clk_i cpu.ROM_addr_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_109_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06781__A1 _02385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06533__A1 _00815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05195__S1 _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09538__A1 net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05090_ _00781_ _00782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05765__I _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08780_ cpu.last_addr\[9\] _03996_ _03997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07800_ _03214_ _03229_ _00249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07731_ cpu.spi.counter\[4\] _03173_ _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05992_ _00980_ _01277_ _01282_ _01654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05575__A2 _01240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04943_ _00643_ _00644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07662_ cpu.uart.receive_buff\[7\] _03093_ _03112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_04874_ cpu.mem_cycle\[1\] cpu.mem_cycle\[0\] _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_46_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09401_ _02351_ _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07593_ cpu.spi.div_counter\[4\] _03058_ _03062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_84_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06613_ _01759_ _02071_ _02268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09332_ _04482_ _04525_ _04526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08277__A1 _01073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06544_ _02178_ _02200_ _02201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_51_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05005__I _00002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09263_ _04458_ _04459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06475_ _00955_ _02131_ _02040_ _00947_ _02132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09194_ _04340_ _04392_ _04393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05426_ _01012_ _01018_ _01021_ _01091_ _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_08214_ _03522_ _03556_ _03519_ _03560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05357_ _01022_ _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_55_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08145_ cpu.toggle_ctr\[15\] _03494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_95_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09529__A1 net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08076_ _03445_ _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05288_ _00955_ _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_30_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07027_ _02387_ _02627_ _02409_ _00078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08978_ _04181_ _04182_ _04183_ _04184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_59_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05566__A2 _01225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06763__A1 _02385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05110__S1 _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07929_ _03328_ _03330_ _03331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06515__A1 _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_20_Left_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08440__A1 cpu.timer_capture\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10305_ _00563_ clknet_leaf_85_wb_clk_i cpu.multiplier.a\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_115_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10236_ _00494_ clknet_leaf_43_wb_clk_i cpu.startup_cycle\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10167_ _00425_ clknet_leaf_37_wb_clk_i cpu.uart.divisor\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10098_ _00357_ clknet_leaf_104_wb_clk_i cpu.pwm_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_32_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_32_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_84_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06260_ cpu.mem_cycle\[3\] _01917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__05168__S1 _00839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07040__I cpu.uart.divisor\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05493__A1 _00910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05211_ _00881_ _00882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06191_ _01471_ _01846_ _01849_ _01850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05142_ cpu.PORTA_DDR\[4\] net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_110_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09950_ _00209_ clknet_4_9_0_wb_clk_i cpu.spi.div_counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05073_ _00743_ _00766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_clkbuf_leaf_49_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08901_ _04108_ _04099_ _04109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06993__A1 _02283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09881_ _00140_ clknet_leaf_112_wb_clk_i cpu.regs\[8\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_90_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05548__A2 _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08832_ _01952_ _04042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08763_ _02404_ _03984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05975_ _01636_ _01176_ _01396_ _01637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07714_ _01891_ _03161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04926_ _00627_ _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08694_ _03929_ _00443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07645_ _03098_ _03094_ _03099_ _03056_ _00224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_0_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07576_ cpu.spi.div_counter\[1\] _03048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_64_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09315_ _04485_ _04507_ cpu.ROM_addr_buff\[2\] _04510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06527_ net123 _02167_ _02184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08046__I _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09246_ _03469_ _00912_ _04442_ _04443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_8_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06458_ _00945_ _02017_ _02066_ _01730_ _02115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_105_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05409_ _00585_ _00595_ _01049_ _01075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__06276__A3 _01932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09177_ _04374_ _04358_ _04375_ _04376_ _04321_ _04377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_71_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_88_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06389_ _02045_ _02025_ _02046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08128_ _03473_ _03481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08422__A1 cpu.timer_capture\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08059_ cpu.PC\[0\] _03432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__06579__A4 _01932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput57 net57 io_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05787__A2 _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput46 net46 io_oeb[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput35 net35 io_oeb[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput79 net79 io_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10021_ _00280_ clknet_leaf_31_wb_clk_i cpu.uart.receive_div_counter\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput68 net68 io_out[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06036__I0 net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output58_I net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05475__A1 _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09496__B _00649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06027__I0 cpu.regs\[8\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10219_ _00477_ clknet_leaf_75_wb_clk_i cpu.PC\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05760_ _01280_ _01423_ _01424_ _01282_ _01425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05691_ _01335_ _01356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07430_ cpu.spi.dout\[3\] _02916_ _02919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07361_ _02220_ _02857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_61_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09100_ _03433_ _02857_ _04301_ _02596_ _04302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_06312_ _01968_ _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09031_ _02389_ _04214_ _04234_ _04235_ _04207_ _04236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_07292_ _02810_ _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06243_ _01899_ _01900_ cpu.spi.counter\[4\] _01889_ _01901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_60_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06174_ cpu.timer_div\[7\] _01398_ _01222_ _01833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_5_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05125_ _00814_ _00815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09933_ _00192_ clknet_leaf_37_wb_clk_i cpu.spi.dout\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05056_ _00731_ _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06018__I0 _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09864_ _00123_ clknet_leaf_111_wb_clk_i cpu.regs\[10\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08815_ _01348_ _04023_ _04024_ _04025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05953__I _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06194__A2 _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09795_ _00058_ clknet_leaf_10_wb_clk_i cpu.timer_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05174__B _00845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08746_ _03160_ _03968_ _03971_ _00453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_84_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05958_ cpu.timer_top\[4\] _01620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08677_ _03915_ _00440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_04909_ _00611_ _00612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09132__A2 _01110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07143__A1 cpu.regs\[12\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05889_ _01166_ _01553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07628_ _03081_ _03087_ _00219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_101_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07559_ _03028_ _03033_ _03034_ _00203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08643__A1 _03885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09229_ _04351_ _04410_ _04427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_51_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06957__A1 _02570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06959__I _02573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_73_Right_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10004_ _00263_ clknet_leaf_22_wb_clk_i cpu.uart.data_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07382__A1 _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_103_Left_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_67_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05696__A1 net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_82_Right_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05999__A2 _00948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_112_Left_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_10_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_91_Right_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06869__I _02470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06930_ _01147_ _02545_ _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA_input1_I io_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08600_ _01169_ _03851_ _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06861_ cpu.timer\[3\] _02490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05812_ _01197_ _01476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06792_ _02431_ _02432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09580_ _02529_ _04711_ _04717_ _00541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08531_ cpu.timer_div\[3\] _03791_ _03774_ _03797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05743_ _01407_ _01234_ _01237_ _01408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05674_ _01158_ _01328_ _01340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_18_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08462_ cpu.timer_capture\[8\] _03746_ _03727_ _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08873__A1 _01116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07413_ _02854_ _02904_ _02905_ _00186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08393_ _02974_ _03679_ _03681_ _03688_ _03684_ _03689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_9_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08625__B2 _03870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07344_ cpu.regs\[3\]\[3\] _02843_ _02845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07275_ _02795_ _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_103_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06226_ cpu.spi.div_counter\[0\] _01884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_85_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09014_ cpu.PC\[4\] _00655_ _04219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06157_ _01816_ cpu.regs\[15\]\[6\] _01167_ _01817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06088_ net31 _01310_ _01749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05108_ _00785_ _00799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__05298__S0 _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05039_ _00732_ _00733_ _00702_ _00734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09916_ _00175_ clknet_leaf_83_wb_clk_i cpu.regs\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06167__A2 _01121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09847_ _00106_ clknet_leaf_106_wb_clk_i cpu.regs\[12\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09778_ _00041_ clknet_leaf_26_wb_clk_i cpu.uart.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08729_ _03916_ cpu.regs\[3\]\[4\] _03957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06728__B _02379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05678__B2 _01333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09493__C _03079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05390_ _01053_ _01055_ _01056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08607__A1 _03836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08607__B2 _01065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07060_ cpu.uart.receive_div_counter\[7\] _02631_ cpu.uart.divisor\[1\] _02639_ _02660_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__09280__A1 _04374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07130__I1 cpu.regs\[13\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06011_ _01543_ _01663_ _01667_ _01672_ _01673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_11_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07962_ _02659_ _03353_ _03234_ _03358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09701_ _04818_ _04824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07893_ cpu.uart.data_buff\[9\] _03264_ _03276_ _03257_ _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06149__A2 _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06913_ _02519_ _02533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09632_ _02297_ _04759_ _02353_ _04760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06844_ cpu.timer\[0\] _02475_ _02476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_87_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09099__A1 _03453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09563_ cpu.PORTB_DDR\[5\] _04704_ _04705_ _04707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06775_ _00651_ _02418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08514_ cpu.spi.divisor\[5\] _03784_ _03786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09494_ net18 _00688_ _03810_ net89 _04660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_81_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05726_ _01390_ _00999_ _01126_ _01391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_65_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05657_ _01158_ _01317_ _01321_ _01323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_08445_ _03729_ _03621_ _03732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05588_ _01253_ _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08376_ _02490_ _03669_ _03673_ _03657_ _03674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_92_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07327_ cpu.regs\[4\]\[5\] _02830_ _02834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09271__A1 _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06085__A1 _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07258_ _02753_ cpu.regs\[7\]\[4\] _02779_ _02790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07189_ _02710_ _02746_ _02748_ _00119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06209_ _01867_ _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_output40_I net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_107_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08837__A1 _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06076__A1 _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_108_Right_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09014__A1 cpu.PC\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_57_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_57_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_20_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04890_ cpu.IO_addr_buff\[7\] cpu.IO_addr_buff\[6\] cpu.IO_addr_buff\[5\] _00593_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_48_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07179__I1 cpu.regs\[11\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07043__I cpu.uart.receive_div_counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06560_ cpu.PC\[3\] _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05511_ _01176_ _01177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06491_ _02112_ _02148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07978__I _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08843__A4 _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05442_ _01107_ _01108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06882__I _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07500__A1 cpu.timer_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08230_ cpu.toggle_ctr\[8\] cpu.toggle_ctr\[7\] _03568_ _03571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_117_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05373_ _00572_ _01037_ _01038_ _01039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_70_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06067__A1 _00950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08161_ _03488_ cpu.toggle_top\[7\] _03509_ _03510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_15_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08092_ cpu.orig_PC\[7\] _03454_ _03457_ _03458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05114__I0 cpu.regs\[8\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07112_ _02696_ _00094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07043_ cpu.uart.receive_div_counter\[0\] _02643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05814__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05290__A2 _00958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08602__I _03839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08994_ _04197_ _04178_ _04198_ _04199_ _04200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07945_ cpu.uart.receive_div_counter\[3\] _03309_ _03342_ _03343_ _03344_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_76_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09615_ net72 _04745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_97_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07876_ _02495_ _03278_ _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06827_ _02460_ _02442_ _02461_ _00044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09546_ _01239_ _04663_ _04695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06758_ _02376_ _02402_ _02405_ _00031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08819__A1 _00811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05709_ _01024_ _01184_ _01374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_66_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09477_ net73 _04644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06689_ _02328_ _02330_ _02341_ _02342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06792__I _02431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08428_ cpu.timer_capture\[11\] _03714_ _03717_ _03690_ _03718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_65_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08359_ _03651_ _03660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06058__A1 cpu.timer_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10252_ _00510_ clknet_leaf_45_wb_clk_i cpu.ROM_spi_cycle\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10183_ _00441_ clknet_leaf_64_wb_clk_i cpu.ROM_addr_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06032__I _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06533__A2 _00948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_104_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_104_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_56_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09235__A1 _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_39_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04950__I _00637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07038__I _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07730_ _03172_ _01891_ _03169_ _03173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08578__B _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05991_ _01280_ _01652_ _01653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_04942_ _00642_ _00643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07721__A1 _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04873_ cpu.mem_cycle\[5\] cpu.mem_cycle\[4\] cpu.mem_cycle\[3\] cpu.mem_cycle\[2\]
+ _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_07661_ cpu.uart.dout\[7\] _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09400_ _04582_ _00496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07592_ _03061_ _00209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_84_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06612_ _02265_ _02266_ _02267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09331_ _04483_ _04524_ _04525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06543_ _02199_ _02200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09474__A1 _03079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08277__A2 _02432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09262_ cpu.PC\[13\] _04433_ _04458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_7_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06474_ _02072_ _02131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09193_ _04388_ _04391_ _04392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_78_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05425_ _01045_ _01056_ _01060_ _01090_ _01091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_08213_ cpu.toggle_ctr\[3\] cpu.toggle_ctr\[2\] _03556_ _03559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_05356_ _00615_ _01022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08144_ cpu.toggle_ctr\[9\] _03492_ _02608_ cpu.toggle_ctr\[8\] _03493_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_16_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05021__I _00704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08075_ _02217_ _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05287_ _00909_ _00955_ _00956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07026_ _02384_ _02627_ _02408_ _00077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_101_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08977_ _04081_ _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_59_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_2_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_2_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07928_ _03329_ _03330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06787__I _02426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05691__I _01335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07859_ _03207_ _03278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_3_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09529_ net80 _04682_ _04683_ _04685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_109_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06736__B _02379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10304_ _00562_ clknet_leaf_84_wb_clk_i cpu.multiplier.a\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10235_ _00493_ clknet_leaf_61_wb_clk_i cpu.startup_cycle\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_115_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06203__A1 _00826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10166_ _00424_ clknet_leaf_27_wb_clk_i cpu.uart.divisor\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10097_ _00356_ clknet_leaf_11_wb_clk_i cpu.pwm_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_112_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05210_ _00880_ _00881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06190_ _01655_ _01848_ _01849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_72_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_72_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05141_ cpu.PORTB_DDR\[4\] net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_25_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05072_ _00765_ net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_08900_ _04107_ _04108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09880_ _00139_ clknet_leaf_113_wb_clk_i cpu.regs\[8\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08831_ _04037_ _04038_ _04039_ _04040_ _04041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_0_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08762_ _03972_ _03982_ _03983_ _00457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05974_ cpu.spi.dout\[4\] _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07713_ _03159_ _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08693_ _03928_ cpu.ROM_addr_buff\[4\] _03921_ _03929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_04925_ _00626_ _00627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07644_ cpu.uart.receive_buff\[2\] _03095_ _03099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07575_ _03043_ _03047_ _00206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_64_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09314_ _03963_ cpu.ROM_addr_buff\[0\] _04509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06526_ net123 _02167_ _02183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_36_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08327__I _03635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09245_ _04440_ _04441_ _04442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_8_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06457_ _01961_ _02113_ _02114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08670__A2 _00696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05408_ _01068_ _01072_ _01073_ _01074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09176_ _00715_ _04351_ _04136_ _04376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06388_ _02022_ _02045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05339_ cpu.br_rel_dest\[5\] _00609_ _00611_ _01004_ _01005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__05686__I _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08127_ _02451_ _03474_ _03480_ _00325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08058_ _02945_ _03423_ _03431_ _00305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput58 net58 io_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_101_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput47 net47 io_oeb[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_07009_ _02447_ _02615_ _02618_ _00069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput36 net36 io_oeb[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput69 net69 io_out[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10020_ _00279_ clknet_leaf_32_wb_clk_i cpu.uart.receive_div_counter\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__06036__I1 cpu.PORTA_DDR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07834__C _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05095__S1 _00786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09686__A1 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08110__A1 _03469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09610__B2 cpu.ROM_addr_buff\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10218_ _00476_ clknet_leaf_76_wb_clk_i cpu.PC\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10149_ _00408_ clknet_leaf_12_wb_clk_i cpu.spi.divisor\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05690_ _01168_ _01353_ _01355_ _00013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05002__I2 _00696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07360_ _02211_ _02856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_61_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06311_ _01967_ _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09030_ _04034_ _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09687__B _04169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07291_ _02810_ _02811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06242_ cpu.spi.counter\[2\] _01900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__05466__A2 _01126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09601__A1 net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06173_ cpu.spi.dout\[7\] _01393_ _01218_ _01831_ _01832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_53_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05124_ _00813_ _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06415__A1 cpu.multiplier.a\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09932_ _00191_ clknet_leaf_38_wb_clk_i cpu.spi.dout\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05055_ _00730_ _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_40_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09863_ _00122_ clknet_leaf_108_wb_clk_i cpu.regs\[10\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06018__I1 cpu.regs\[15\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08814_ _03903_ _01330_ _01436_ _04024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_09794_ _00057_ clknet_leaf_9_wb_clk_i cpu.timer_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08745_ cpu.ROM_addr_buff\[0\] _03970_ _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05957_ _01618_ _01619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08676_ _03914_ cpu.ROM_addr_buff\[1\] _03813_ _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_68_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04908_ cpu.base_address\[1\] cpu.base_address\[0\] _00610_ _00611_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_05888_ _01551_ _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08340__A1 cpu.timer_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07627_ cpu.spi.data_in_buff\[4\] _03083_ _03085_ cpu.spi.data_in_buff\[5\] _03087_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_101_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07558_ cpu.spi.data_out_buff\[4\] _03011_ _03026_ _03034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06509_ _02139_ _02165_ _02166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07489_ cpu.timer_top\[6\] _02972_ _02973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_91_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09228_ _04137_ _04410_ _04425_ _04162_ _04426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09159_ cpu.orig_PC\[9\] _04244_ _04359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output70_I net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10003_ _00262_ clknet_leaf_22_wb_clk_i cpu.uart.data_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07382__A2 _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07580__B _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08331__A1 cpu.timer_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08882__A2 _00984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_78_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06948__A2 _02557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09526__I _04674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06860_ _00933_ _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05811_ net41 _01190_ _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_38_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06791_ _02429_ _02430_ _02431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_54_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05223__I2 cpu.regs\[6\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08530_ _02450_ _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05742_ cpu.timer_capture\[9\] _01407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_49_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05673_ _00712_ _01333_ _01339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08461_ _03739_ _03746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07412_ _00748_ _02869_ _02905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08392_ cpu.timer\[5\] _03687_ _03688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_73_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07343_ _01551_ _02839_ _02844_ _00177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07274_ _02783_ _02797_ _02800_ _00152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06636__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06225_ cpu.spi.div_counter\[6\] cpu.spi.divisor\[6\] _01883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09013_ _02215_ _01618_ _04218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08389__A1 cpu.timer_capture\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06156_ _01815_ _01816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07061__A1 _02648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07061__B2 _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06087_ _01313_ _01747_ _01748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05298__S1 _00899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05107_ cpu.multiplier.a\[6\] _00798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09915_ _00174_ clknet_leaf_89_wb_clk_i cpu.regs\[4\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05038_ cpu.regs\[4\]\[2\] cpu.regs\[5\]\[2\] cpu.regs\[6\]\[2\] cpu.regs\[7\]\[2\]
+ _00730_ _00731_ _00733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09846_ _00105_ clknet_leaf_107_wb_clk_i cpu.regs\[12\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09777_ _00040_ clknet_leaf_36_wb_clk_i cpu.uart.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05375__A1 _00652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06989_ net119 _02079_ _02601_ _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08728_ _03956_ _00450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08659_ _02376_ _03900_ _03902_ _00435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_95_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06627__A1 cpu.regs\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09041__A2 _04244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07355__A2 _01906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05823__B _01142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08855__A2 _04008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04953__I _00652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06010_ _01670_ _01343_ _01671_ _01341_ _01434_ _01672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_112_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08791__A1 _00686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07961_ _02659_ _03345_ _03346_ _03356_ _03357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07594__A2 _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06912_ _02453_ _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09700_ _01468_ _04820_ _04823_ _00555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07892_ _03291_ _03302_ _03304_ _00266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08543__A1 _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09631_ _02311_ _04756_ _04758_ _04759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06843_ _02472_ _02475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06774_ _02376_ _02415_ _02417_ _00035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09562_ _02532_ _04703_ _04706_ _00534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05725_ cpu.spi.divisor\[1\] _01390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_08513_ _02532_ _03783_ _03785_ _00406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05225__S _00832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08846__A2 _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06157__I0 _01816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09493_ _04644_ _04657_ _04658_ _04659_ _03079_ _00512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_93_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06857__A1 _00906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05656_ _01158_ _01317_ _01321_ _01322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08444_ _03729_ _03730_ _03731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_105_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05587_ _01083_ _01085_ _01253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08375_ _02975_ _03667_ _03673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05959__I net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07326_ _02833_ _00171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07257_ _02788_ _02780_ _02789_ _00146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09023__A2 _03854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06208_ _01850_ _01851_ _01866_ _01432_ _01867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_07188_ cpu.regs\[10\]\[0\] _02747_ _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07034__B2 _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07034__A1 cpu.uart.divisor\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06139_ _01798_ _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09166__I _04147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05596__A1 cpu.toggle_top\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09829_ _00088_ clknet_leaf_99_wb_clk_i cpu.regs\[14\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07350__S _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09014__A2 _00655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_29_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08773__A1 cpu.ROM_addr_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05131__S0 _00816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_97_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_97_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_26_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_26_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_48_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08828__A2 _01990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05510_ _01009_ _01175_ _01176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_47_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06490_ _02137_ _02143_ _02146_ _02147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_05441_ cpu.br_rel_dest\[3\] _01107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_68_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08160_ _03491_ _03493_ _03503_ _03508_ _03509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_43_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05372_ _00574_ _01038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08155__I cpu.toggle_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07111_ cpu.regs\[14\]\[7\] _02283_ _02692_ _02696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08091_ _03456_ _03457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_82_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07042_ _01209_ _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_3_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08993_ _04106_ _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07944_ _02662_ _03340_ _03343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07875_ _03269_ _03291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08516__A1 cpu.spi.divisor\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09614_ _04744_ _00548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06826_ cpu.uart.divisor\[5\] _02435_ _02457_ _02461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09545_ _03833_ _04688_ _04694_ _00529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06757_ _01169_ _02401_ _02404_ _02405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08819__A2 _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09476_ _04558_ _04643_ _00511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06688_ _02333_ _02336_ _02340_ _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05708_ net7 _01204_ _01373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05639_ _01303_ _01299_ _01304_ _01305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08427_ _02953_ _03668_ _03680_ _03716_ _03677_ _03717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_108_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08358_ cpu.timer\[0\] _03657_ _03658_ _03659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07309_ _02822_ _00165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08289_ _02447_ _03604_ _03611_ _00356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_104_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10251_ _00509_ clknet_leaf_45_wb_clk_i cpu.ROM_spi_cycle\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07007__A1 _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10182_ _00440_ clknet_leaf_63_wb_clk_i cpu.ROM_addr_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_70_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08507__A1 _02527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_102_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08703__I _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08746__A1 _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05990_ _00957_ _01265_ _01651_ _01137_ _01652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_04941_ _00566_ _00642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05980__A1 cpu.timer_capture\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04872_ _00572_ _00573_ _00574_ _00575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_07660_ _03109_ _03101_ _03110_ _03104_ _00228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07591_ _03057_ _03059_ _03060_ _03061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_84_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06611_ _02246_ _02248_ _02266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09330_ _02337_ _02395_ _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06542_ _02182_ _02198_ _02199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09261_ cpu.PC\[13\] _04379_ _04457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08212_ _03553_ _03558_ _00332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06473_ _00813_ _02130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_09192_ _04362_ _04389_ _04390_ _04391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05424_ _01011_ _01082_ _01086_ _01089_ _01090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_16_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05355_ _01020_ _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_55_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08143_ cpu.toggle_top\[9\] _03492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08074_ _03442_ _03434_ _03444_ _00308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08613__I _03863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08985__A1 _04173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07025_ _02381_ _02627_ _02407_ _00076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05286_ _00954_ _00955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_30_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input32_I sram_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08976_ _04173_ _01108_ _04182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07927_ _03306_ _02666_ _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_59_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07858_ _03273_ _03275_ _03277_ _00259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07789_ _03138_ _03219_ _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06809_ _02446_ _02447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_3_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07899__I _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09528_ _03815_ _04681_ _04684_ _00522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_104_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08009__B _03395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09459_ cpu.ROM_spi_cycle\[3\] _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_93_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08976__A1 _04173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10303_ _00561_ clknet_leaf_92_wb_clk_i cpu.regs\[9\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10234_ _00492_ clknet_leaf_60_wb_clk_i cpu.startup_cycle\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_115_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10165_ _00423_ clknet_leaf_27_wb_clk_i cpu.uart.divisor\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06203__A2 _01759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07400__A1 _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10096_ _00355_ clknet_leaf_3_wb_clk_i cpu.pwm_top\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09456__A2 _04592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06218__I cpu.spi.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05122__I cpu.multiplier.a\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07219__A1 _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08416__B1 _03681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05140_ cpu.PORTA_DDR\[3\] net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_25_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05071_ _00764_ _00765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_41_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_41_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07049__I _02648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08830_ _01531_ _00728_ _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_90_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06888__I _02465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08761_ cpu.ROM_addr_buff\[4\] _03976_ _03983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05973_ _01213_ _01175_ _01634_ _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09144__A1 _00984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08692_ _02556_ _03917_ _03927_ _03928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04924_ _00619_ _00626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_07712_ _02403_ _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07643_ cpu.uart.dout\[2\] _03098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09313_ _03920_ _04485_ _04507_ _04508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09447__A2 _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07574_ _03044_ _03045_ _03046_ _03047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_64_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06525_ _02181_ _02182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09244_ cpu.PC\[11\] _00877_ _04419_ _04441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06456_ _01798_ _01993_ _01995_ _01296_ _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_105_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09175_ _04166_ _04357_ _04375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05407_ _01014_ _01029_ _01073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_44_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06387_ _02041_ _02043_ _02044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08126_ cpu.toggle_top\[3\] _03475_ _03477_ _03480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05338_ _00647_ cpu.instr_cycle\[2\] _00576_ _00577_ _01004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_113_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08057_ cpu.orig_flags\[3\] _03428_ _03430_ _03431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05236__A3 _00906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05269_ _00006_ _00937_ _00938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_113_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput48 net48 io_oeb[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_07008_ cpu.toggle_top\[10\] _02612_ _02616_ _02618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput37 net37 io_oeb[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput59 net59 io_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06197__A1 _00810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05244__I0 _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08959_ _04165_ _04166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05944__A1 _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09686__A2 _02465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09123__B _04324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08110__A2 _03404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06121__A1 cpu.timer_capture\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08949__A1 _00661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08253__I _03370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05307__S0 _00891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10217_ _00475_ clknet_leaf_73_wb_clk_i cpu.PC\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06188__A1 _01618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06027__I2 cpu.regs\[10\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10148_ _00407_ clknet_leaf_12_wb_clk_i cpu.spi.divisor\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09126__A1 _03432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10079_ _00338_ clknet_leaf_118_wb_clk_i cpu.toggle_ctr\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08856__C _04035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09677__A2 _00884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07290_ _02809_ _02810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_17_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06310_ _00714_ _01967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06241_ cpu.spi.counter\[3\] _01899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07860__A1 _02480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06172_ _01828_ _01829_ _01830_ _01831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08163__I cpu.toggle_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07612__A1 _01896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05123_ _00812_ _00813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09931_ _00190_ clknet_leaf_38_wb_clk_i cpu.spi.dout\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05054_ cpu.regs\[2\]\[3\] _00748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_110_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09208__B _04324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09862_ _00121_ clknet_leaf_108_wb_clk_i cpu.regs\[10\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08813_ _01438_ _01461_ _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09793_ _00056_ clknet_leaf_10_wb_clk_i cpu.timer_top\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08744_ _03969_ _03970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05956_ cpu.br_rel_dest\[4\] _01618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__09668__A2 _04244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04907_ cpu.base_address\[3\] cpu.base_address\[2\] _00610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08675_ _03439_ _00649_ _03913_ _03914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05887_ _01550_ _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07626_ _03081_ _03086_ _00218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08338__I _03635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07557_ cpu.spi.data_out_buff\[5\] _03021_ _03032_ _03033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06508_ _02142_ _02165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_36_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06103__A1 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07488_ cpu.timer\[6\] _02972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09227_ _04412_ _04424_ _04425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07851__A1 _02677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06439_ _02064_ _02068_ _02096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_16_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09158_ _04357_ _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08109_ cpu.orig_PC\[12\] _03464_ _03467_ _03470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09089_ _04285_ _04289_ _04291_ _04292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_112_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08159__A2 _01842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output63_I net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08022__B _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10002_ _00261_ clknet_leaf_22_wb_clk_i cpu.uart.data_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05393__A2 _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06590__A1 _02119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_17_Left_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_26_Left_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05810_ _01472_ _01473_ _01363_ _01474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06790_ _00639_ _00668_ _02430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07263__S _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08858__B1 _04036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05741_ _01228_ _01405_ _01406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05672_ _00712_ _01335_ _01337_ _01338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08460_ _03702_ _03742_ _03744_ _03745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08391_ _02490_ _02498_ _03667_ _03687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_46_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_35_Left_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07411_ _01613_ _02234_ _02903_ _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07342_ cpu.regs\[3\]\[2\] _02843_ _02844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07273_ cpu.regs\[6\]\[1\] _02798_ _02800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06636__A2 _02229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06224_ cpu.spi.div_counter\[5\] cpu.spi.divisor\[5\] _01882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09012_ _04181_ _04215_ _04216_ _04217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_14_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_1_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09586__A1 cpu.PORTA_DDR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06155_ _01814_ _01815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05106_ _00766_ _00797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_44_Left_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06086_ _01315_ net95 _01746_ _01747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09338__A1 _03588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09914_ _00173_ clknet_leaf_91_wb_clk_i cpu.regs\[4\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05037_ cpu.regs\[0\]\[2\] _00728_ _00729_ cpu.regs\[3\]\[2\] _00730_ _00731_ _00732_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09845_ _00104_ clknet_leaf_105_wb_clk_i cpu.regs\[12\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09776_ _00039_ clknet_leaf_18_wb_clk_i cpu.uart.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_06988_ net119 _02079_ _02558_ _02601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08727_ _03955_ cpu.ROM_addr_buff\[11\] _03952_ _03956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05939_ cpu.pwm_top\[3\] _01251_ _01601_ _01253_ _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09510__A1 _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08658_ _00984_ _03901_ _03830_ _03902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_53_Left_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07609_ _01873_ _03002_ _03070_ _03075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_4_8_0_wb_clk_i clknet_0_wb_clk_i clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08589_ _03840_ _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_83_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09120__C _04321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07824__A1 _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_19_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_62_Left_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09577__A1 cpu.PORTA_DDR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06760__B _02406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_71_Left_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05366__A2 _01031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_58_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09568__A1 _03833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09537__I _04674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07258__S _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07960_ _02659_ _03353_ _03356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06911_ _02529_ _02520_ _02530_ _02531_ _00058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07891_ cpu.uart.data_buff\[9\] _03266_ _03303_ _03304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09630_ _04757_ _04758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_65_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06842_ _02470_ _02474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06773_ _02416_ _02414_ _02406_ _02417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09561_ cpu.PORTB_DDR\[4\] _04704_ _04705_ _04706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_97_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05724_ _01387_ _01388_ _01134_ _01389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08512_ cpu.spi.divisor\[4\] _03784_ _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09492_ _03584_ cpu.pwm_counter\[1\] cpu.pwm_counter\[3\] _03589_ _04659_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_93_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05655_ _00711_ _01320_ _01321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_18_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08443_ _02965_ _02949_ _03719_ _03730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_73_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08616__I _03850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08374_ _03653_ _03671_ _03672_ _00380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05586_ _01251_ _01252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07325_ _02818_ cpu.regs\[4\]\[4\] _02825_ _02833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07256_ cpu.regs\[7\]\[3\] _02786_ _02789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06207_ _01852_ _01527_ _01462_ _01865_ _01866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_33_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07187_ _02745_ _02747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06138_ _01797_ _01798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06069_ _00967_ _00971_ _00976_ _00974_ _01730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_09828_ _00087_ clknet_leaf_99_wb_clk_i cpu.regs\[14\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09759_ _00022_ clknet_leaf_97_wb_clk_i cpu.regs\[2\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08298__A1 cpu.pwm_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06784__A1 _02388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05587__A2 _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05131__S1 _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06536__A1 _01941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09722__A1 _03439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_66_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_66_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_86_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05125__I _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08289__A1 _02447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04964__I _00663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05440_ _01100_ _01105_ _01106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05371_ _00573_ _01037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07110_ _02695_ _00093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08090_ _02455_ _03456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__05114__I2 cpu.regs\[10\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07041_ cpu.uart.receive_div_counter\[10\] _02641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_11_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08992_ cpu.orig_PC\[3\] _03841_ _04198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07943_ _03335_ _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07874_ _03273_ _03287_ _03290_ _00262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09713__A1 _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09613_ net65 _04735_ _04737_ _04743_ _02439_ _04744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_06825_ _02459_ _02460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09544_ net58 _04689_ _04690_ _04694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06756_ _02403_ _02404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__05035__I _00716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09475_ net74 _03551_ _04643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06687_ _02337_ _02339_ _02340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_05707_ _01366_ _01368_ _01371_ _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05638_ _01012_ _01018_ _01021_ _01091_ _01304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_08426_ _02953_ _03715_ _03716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_19_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05569_ _01026_ _01031_ _01235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_46_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08357_ cpu.timer\[0\] _03654_ _03658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07308_ _02821_ cpu.regs\[5\]\[6\] _02810_ _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08288_ cpu.pwm_top\[2\] _03605_ _03609_ _03611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07239_ _02742_ _02766_ _02775_ _00142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10250_ _00508_ clknet_leaf_45_wb_clk_i cpu.ROM_spi_cycle\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10181_ _00439_ clknet_leaf_72_wb_clk_i cpu.ROM_addr_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05569__A2 _01031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07191__A1 _02717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_53_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07246__A2 _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_113_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_113_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_40_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06757__A1 _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04940_ _00635_ _00640_ _00641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07335__I _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04871_ cpu.startup_cycle\[3\] cpu.startup_cycle\[2\] _00574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_79_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07182__A1 cpu.regs\[11\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07590_ _01879_ _03052_ _01872_ _03060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_9_Left_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06610_ _02186_ _02247_ _02265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06541_ _02185_ _02189_ _02197_ _02198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09260_ _04432_ _04456_ _04431_ _00482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06472_ _02119_ _00917_ _02129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05496__A1 _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05423_ _01083_ _01088_ _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08211_ _03523_ _03556_ _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09191_ cpu.PC\[9\] _00881_ _04390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05354_ _01016_ _01019_ _01020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08142_ _03489_ _02620_ cpu.toggle_top\[11\] _03490_ _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__08434__A1 cpu.timer_capture\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08073_ cpu.orig_PC\[2\] _03443_ _03430_ _03444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05285_ _00953_ _00954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07024_ _02375_ _02627_ _02405_ _00075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08975_ _04141_ _04142_ _04180_ _04181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07926_ cpu.uart.receive_div_counter\[0\] _03328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_59_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07245__I _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input25_I rst_n vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07857_ cpu.uart.data_buff\[2\] _03276_ _03041_ _03277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07788_ _03129_ _03218_ _03220_ _03113_ _00246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06808_ _00905_ _02446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_3_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09527_ net79 _04682_ _04683_ _04684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06739_ _02387_ _02388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_104_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09458_ _00568_ _04630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05487__A1 _00650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09389_ _04568_ _04571_ _02914_ _04574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05487__B2 _00882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08409_ cpu.timer\[8\] _03702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08976__A2 _01108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output93_I net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10302_ _00560_ clknet_leaf_92_wb_clk_i cpu.regs\[9\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06987__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10233_ _00491_ clknet_leaf_60_wb_clk_i cpu.startup_cycle\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10164_ _00422_ clknet_leaf_27_wb_clk_i cpu.uart.divisor\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10095_ _00354_ clknet_leaf_3_wb_clk_i cpu.pwm_top\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06911__A1 _02529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05270__S0 _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08664__A1 _00913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05022__S0 _00716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07219__A2 _02729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05070_ _00763_ _00764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_4_6_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_10_0_wb_clk_i clknet_0_wb_clk_i clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_57_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08760_ _03980_ _03981_ _03982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05972_ cpu.spi.divisor\[4\] _01180_ _01634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_81_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_81_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_04923_ cpu.TIE cpu.needs_timer_interrupt _00625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08691_ _03926_ _00769_ _03927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07711_ _03114_ _03152_ _03153_ _00236_ _00230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_73_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07155__A1 cpu.regs\[12\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_10_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_10_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07642_ _01385_ _03094_ _03097_ _03056_ _00223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_79_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09312_ cpu.last_addr\[1\] _03963_ cpu.last_addr\[2\] _04507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07573_ _03044_ _01902_ _03046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_87_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05313__I _00980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06524_ _02160_ _02179_ _02180_ _02181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09243_ _02206_ _01099_ _04440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06455_ _02111_ _02106_ _02112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09174_ _00679_ _04374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05406_ _01064_ _01071_ _01072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_63_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06386_ _00783_ _02042_ _02043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08407__A1 cpu.timer_capture\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05337_ _01002_ _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08125_ _02447_ _03474_ _03479_ _00324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08056_ _03410_ _03430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05268_ cpu.regs\[4\]\[4\] cpu.regs\[5\]\[4\] cpu.regs\[6\]\[4\] cpu.regs\[7\]\[4\]
+ _00890_ _00892_ _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_101_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput49 net49 io_oeb[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_05199_ net127 _00871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07007_ _02614_ _02615_ _02617_ _00068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput38 net38 io_oeb[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07394__A1 _02573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08958_ _04091_ _04165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07909_ cpu.uart.receive_buff\[2\] _03313_ _03316_ cpu.uart.receive_buff\[1\] _03318_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_98_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08889_ _04074_ _04097_ _03395_ _00470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_85_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05880__A1 _00904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09071__A1 _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05307__S1 _00893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10216_ _00474_ clknet_leaf_76_wb_clk_i cpu.PC\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06027__I3 cpu.regs\[11\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07385__A1 _01466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10147_ _00406_ clknet_leaf_12_wb_clk_i cpu.spi.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10078_ _00337_ clknet_leaf_118_wb_clk_i cpu.toggle_ctr\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_99_Left_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_72_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06240_ _01888_ _01898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05871__A1 _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06171_ cpu.spi.divisor\[7\] _01180_ _01181_ _01830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_80_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05122_ cpu.multiplier.a\[7\] _00812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09930_ _00189_ clknet_leaf_37_wb_clk_i cpu.spi.dout\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_92_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05053_ _00746_ _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_5_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09861_ _00120_ clknet_leaf_111_wb_clk_i cpu.regs\[10\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07376__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08812_ _04020_ _04022_ _03395_ _00468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09792_ _00055_ clknet_leaf_9_wb_clk_i cpu.timer_top\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08743_ _02366_ _03965_ _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_05955_ _01168_ _01616_ _01617_ _00016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_108_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_04906_ _00607_ cpu.instr_buff\[14\] _00608_ cpu.base_address\[4\] _00609_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_08674_ _03909_ _00715_ _03913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08876__A1 _03432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05886_ _01549_ _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07625_ cpu.spi.data_in_buff\[3\] _03083_ _03085_ cpu.spi.data_in_buff\[4\] _03086_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_101_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07556_ _02503_ _03022_ _03032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08628__A1 _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06507_ _02163_ _02164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_91_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09226_ _04346_ _04423_ _04424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07487_ _02970_ _02514_ _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06438_ _02064_ _02068_ _02095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_90_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09157_ _02222_ _04212_ _04356_ _03461_ _04357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__05862__A1 _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06369_ _02022_ _02025_ _02026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_44_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07064__B1 _02662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08108_ cpu.PC\[12\] _03469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09088_ _04010_ _04276_ _04290_ _04158_ _04291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_31_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08039_ _03407_ _03418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_112_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10001_ _00260_ clknet_leaf_21_wb_clk_i cpu.uart.data_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output56_I net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10225__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05888__I _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05853__B2 _00884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_87_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04967__I _00654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05740_ cpu.timer_capture\[1\] _01223_ _01405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08439__I _03608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05671_ _01327_ _01098_ _01336_ _00856_ _01337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_58_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08390_ _03686_ _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_46_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07410_ _02259_ _02902_ _02903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_73_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07341_ _02837_ _02843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07272_ _02776_ _02797_ _02799_ _00151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06223_ cpu.spi.div_counter\[0\] _01178_ cpu.spi.divisor\[2\] _01879_ _01880_ _01881_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_09011_ _02217_ _01107_ _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07046__B1 _01183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06154_ _01796_ _01813_ _01814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XPHY_EDGE_ROW_103_Right_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05105_ _00796_ net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_41_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06085_ _01316_ _01739_ _01742_ _01745_ _01746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_41_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09913_ _00172_ clknet_leaf_89_wb_clk_i cpu.regs\[4\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05036_ _00717_ _00731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07349__A1 _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07962__B _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09844_ _00103_ clknet_leaf_105_wb_clk_i cpu.regs\[12\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06572__A2 _01040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09775_ _00038_ clknet_leaf_14_wb_clk_i cpu.br_rel_dest\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06987_ net20 _02559_ _02600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08726_ _03466_ _03949_ _03954_ _03955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05938_ _01597_ _01599_ _01600_ _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_96_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08657_ _03899_ _03901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05869_ _00909_ _00916_ _01532_ _01533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07521__A1 cpu.spi.data_out_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07608_ cpu.spi.div_counter\[7\] _03071_ _03074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07372__I1 _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08588_ _03839_ _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07539_ _02446_ _03008_ _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06088__A1 net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07824__A2 _01895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09209_ _02207_ _04379_ _04407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05835__A1 cpu.timer_capture\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_73_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_4_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07512__A1 _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04877__A2 _00579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09265__A1 _02254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05826__A1 cpu.spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08722__I _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06910_ _02523_ _02531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07890_ _03025_ _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_65_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06841_ _02472_ _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06772_ _01267_ _02416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09560_ _02378_ _04705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08169__I cpu.toggle_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05723_ cpu.uart.has_byte _01136_ _01388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08511_ _03776_ _03784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09491_ cpu.pwm_counter\[5\] _03594_ cpu.pwm_counter\[7\] cpu.pwm_counter\[6\] _04658_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_08442_ cpu.timer\[14\] _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05654_ _01319_ _00879_ _01320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05585_ _01083_ _01073_ _01251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_46_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08373_ cpu.timer_capture\[2\] _03660_ _03615_ _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07324_ _02788_ _02826_ _02832_ _00170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05817__A1 net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05321__I _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07255_ _01614_ _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06206_ _01315_ net97 _01864_ _01865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07186_ _02745_ _02746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06137_ _01682_ _01684_ _01689_ _01687_ _01797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_06068_ _01140_ _01170_ _01728_ _01729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__07248__I _01467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05045__A2 _00737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05019_ cpu.regs\[2\]\[1\] _00715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09827_ _00086_ clknet_leaf_80_wb_clk_i _00003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_09758_ _00021_ clknet_leaf_40_wb_clk_i net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_69_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08709_ _03941_ _00446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_68_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09689_ _04035_ _04799_ _04814_ _04815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_107_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09247__A1 _04138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06233__A1 _01888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07733__A1 _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05339__A3 _00611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06946__B _02203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09238__A1 _03469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05370_ _00655_ _01036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_35_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_35_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_15_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09548__I _04695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05114__I3 cpu.regs\[11\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07040_ cpu.uart.divisor\[10\] _02640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__05275__A2 _00006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06472__A1 _02119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08991_ _04009_ _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07942_ _02630_ _03339_ _03341_ _03310_ _00279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07873_ cpu.uart.data_buff\[5\] _03288_ _03289_ _03290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07724__A1 _02440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09612_ _04740_ _04741_ _04742_ _04743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06824_ _00981_ _02459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07017__B _02623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09543_ _03804_ _04688_ _04693_ _00528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_92_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06755_ _00620_ _02403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06686_ _01918_ _02338_ _02321_ _02339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09474_ _03079_ _04639_ _04642_ _00510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05706_ _01369_ _01189_ _01370_ _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05637_ _01302_ _01303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08425_ _02989_ _03710_ _03715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_108_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08356_ _03656_ _03657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05568_ _01233_ _01234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07307_ _01814_ _02821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08287_ _02614_ _03604_ _03610_ _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_33_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05499_ _01148_ _01154_ _01164_ _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_07238_ cpu.regs\[8\]\[7\] _02769_ _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06463__A1 _02119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07169_ _02717_ _02732_ _02735_ _00112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10180_ _00438_ clknet_leaf_78_wb_clk_i cpu.base_address\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_70_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07715__A1 _01897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05226__I _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08691__A2 _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04870_ cpu.startup_cycle\[6\] cpu.startup_cycle\[5\] cpu.startup_cycle\[4\] _00573_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_99_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06540_ _02190_ _02196_ _02197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06471_ _02104_ _02126_ _02127_ _02128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__08131__A1 _02454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06693__A1 _00622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05422_ _01030_ _01087_ _01088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08210_ _03555_ _03556_ _03557_ _00331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09190_ cpu.PC\[9\] _00881_ _04389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05353_ _00996_ _01013_ _01019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08141_ cpu.toggle_ctr\[11\] _03490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08072_ _03407_ _03443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05284_ _00952_ _00953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_31_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07023_ _02401_ _02627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08974_ _04143_ _04180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07925_ _03213_ _03327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_89_Right_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05420__A2 _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09698__A1 _01352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07856_ _03269_ _03276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input18_I io_in[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08785__C _03993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06807_ _02440_ _02445_ _00040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07787_ cpu.uart.div_counter\[9\] _03184_ _03181_ _03219_ _03220_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_04999_ cpu.regs\[2\]\[0\] _00696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_94_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04931__A1 cpu.IE vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09526_ _04674_ _04683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06738_ net20 _02374_ _02387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09457_ _04628_ _04629_ _00506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08122__A1 _01417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06669_ _01913_ _02316_ _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_98_Right_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_22_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08408_ _03663_ _03700_ _03701_ _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09388_ _04568_ _04556_ _04569_ _04572_ _04573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_93_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08339_ _03635_ _03644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09622__B2 cpu.ROM_addr_buff\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10301_ _00559_ clknet_leaf_109_wb_clk_i cpu.regs\[9\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10232_ _00490_ clknet_leaf_43_wb_clk_i cpu.startup_cycle\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10163_ _00421_ clknet_leaf_27_wb_clk_i cpu.uart.divisor\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09137__B _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09689__A1 _04035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10094_ _00353_ clknet_leaf_103_wb_clk_i cpu.pwm_counter\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_83_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05270__S1 _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08113__A1 _02440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05022__S1 _00717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09613__B2 _04743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09098__I _04101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06427__B2 _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04989__A1 _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05971_ _01630_ _01631_ _01632_ _01633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07710_ _03158_ _00236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08690_ _03908_ _03926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04922_ _00617_ _00621_ _00623_ _00624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_07641_ cpu.uart.receive_buff\[1\] _03095_ _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_73_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07572_ _01897_ _02910_ _03045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_0_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09311_ cpu.last_addr\[1\] cpu.ROM_addr_buff\[1\] _03963_ _04506_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xclkbuf_leaf_50_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_50_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_48_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06523_ _02168_ _02172_ _02180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_36_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09242_ _04197_ _04437_ _04438_ _04199_ _04439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_8_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06454_ _02110_ _02108_ _02111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_90_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09173_ _04300_ _04358_ _04372_ _04317_ _04373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05405_ _01070_ _01071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06385_ _00854_ _02018_ _02002_ _00915_ _02042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05336_ _01001_ _01002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08124_ cpu.toggle_top\[2\] _03475_ _03477_ _03479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08055_ _03427_ _03423_ _03429_ _00304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05267_ _00935_ _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07006_ cpu.toggle_top\[9\] _02612_ _02616_ _02617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05198_ _00869_ _00864_ _00870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
Xoutput39 net39 io_oeb[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08957_ _04136_ _04163_ _04164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07908_ _03243_ _03317_ _00269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08888_ _00644_ _00689_ _02428_ _04096_ _04097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07839_ _03152_ _03259_ _03261_ _03252_ _03262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08087__I _03400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08894__A2 _04101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_38_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09509_ net62 _04666_ _04667_ _04671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_117_Right_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_93_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09071__A2 _04273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10215_ _00473_ clknet_leaf_76_wb_clk_i cpu.PC\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08582__A1 _03833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06070__I _01730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10146_ _00405_ clknet_leaf_15_wb_clk_i cpu.spi.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10077_ _00336_ clknet_leaf_118_wb_clk_i cpu.toggle_ctr\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05320__A1 _00984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06245__I _00626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06170_ cpu.uart.dout\[7\] _01023_ _01589_ _01829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_80_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05121_ _00811_ net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_13_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05052_ _00745_ _00746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09860_ _00119_ clknet_leaf_111_wb_clk_i cpu.regs\[10\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08573__A1 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08811_ cpu.orig_flags\[2\] _04017_ _04014_ _04021_ _04022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_84_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09791_ _00054_ clknet_leaf_7_wb_clk_i cpu.timer_capture\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08742_ _03963_ _03967_ _03968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05954_ cpu.regs\[15\]\[3\] _01553_ _01617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08673_ _03912_ _00439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_04905_ cpu.base_address\[5\] _00608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_07624_ _03077_ _03085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05885_ _01524_ _01526_ _01548_ _01307_ _01549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_88_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07555_ _03028_ _03030_ _03031_ _00202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06506_ _00813_ _02162_ _02163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06639__A1 cpu.regs\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07486_ cpu.timer_top\[7\] _02970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09225_ _04254_ _04416_ _04422_ _04423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06437_ _02093_ _02089_ _02094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09156_ _04325_ _04327_ _04356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06368_ _01980_ _02023_ _02024_ _02025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06155__I _01814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07064__B2 cpu.uart.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08107_ _03466_ _03459_ _03468_ _00317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09087_ cpu.orig_PC\[6\] _03854_ _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06299_ _00714_ _00727_ _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05319_ _00985_ _00986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06811__A1 _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08038_ cpu.IO_addr_buff\[6\] _03417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_111_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08564__A1 _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10000_ _00259_ clknet_leaf_21_wb_clk_i cpu.uart.data_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09989_ _00248_ clknet_leaf_25_wb_clk_i cpu.uart.div_counter\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_67_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06878__A1 _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05234__I _00904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08280__I _03602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10129_ _00388_ clknet_leaf_1_wb_clk_i cpu.timer\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08858__A2 _03870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05670_ _01156_ _01336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_54_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05144__I cpu.PORTA_DDR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07340_ _01468_ _02839_ _02842_ _00176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08455__I _03739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09010_ cpu.PC\[3\] cpu.br_rel_dest\[3\] _04215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07271_ cpu.regs\[6\]\[0\] _02798_ _02799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_rebuffer8_I _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06222_ _01878_ cpu.spi.divisor\[2\] cpu.spi.divisor\[3\] _01871_ _01880_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__09035__A2 _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07046__B2 cpu.uart.receive_div_counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06153_ net32 _01527_ _01311_ _01812_ _01813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_5_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08794__A1 _00686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05104_ _00766_ _00789_ _00795_ _00796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_111_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06084_ _01457_ _01743_ _01744_ _01332_ _01745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_13_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08546__A1 _00648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09912_ _00171_ clknet_leaf_91_wb_clk_i cpu.regs\[4\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05035_ _00716_ _00730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05319__I _00985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09843_ _00102_ clknet_leaf_96_wb_clk_i cpu.regs\[13\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09774_ _00037_ clknet_leaf_14_wb_clk_i cpu.br_rel_dest\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_06986_ _02597_ _02598_ _02599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05255__S _00830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05937_ cpu.timer_top\[11\] _01242_ _01248_ _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08725_ _03942_ cpu.regs\[3\]\[3\] _03954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_95_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08656_ _03899_ _03900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05868_ _00909_ _01531_ _01532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07607_ _03043_ _03073_ _00212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08587_ _00603_ _00656_ _03839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_49_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07538_ _03013_ _03015_ _03017_ _00199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05799_ _01438_ _01461_ _01463_ _01464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09274__A2 _03863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07469_ cpu.timer\[11\] _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_91_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09208_ _04380_ _04406_ _04324_ _00480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_51_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07037__B2 _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09139_ _04110_ _04340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05599__A1 _01057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07444__I _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_107_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_107_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07276__A1 cpu.regs\[6\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08776__A1 cpu.last_addr\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05139__I cpu.PORTB_DDR\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08528__A1 _00919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06840_ _01220_ _02472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06771_ _02414_ _02415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05722_ _00993_ _01213_ _01384_ _01386_ _01387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_08510_ _03776_ _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09490_ _04650_ _04653_ _04656_ _04657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_81_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05653_ _00908_ _00870_ _01318_ _01319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08441_ _03663_ _03726_ _03728_ _00391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_105_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08372_ _03669_ _03670_ _03671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05584_ cpu.timer_top\[8\] _01247_ _01249_ _01250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_85_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07267__A1 _02684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07323_ cpu.regs\[4\]\[3\] _02830_ _02832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07254_ _02785_ _02780_ _02787_ _00145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06205_ _01316_ _01858_ _01860_ _01863_ _01864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07019__A1 cpu.toggle_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07185_ _02744_ _02745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_30_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06136_ _01306_ _01795_ _01796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06067_ _00950_ _01283_ _01655_ _01727_ _01728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__08519__A1 _02540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05018_ cpu.multiplier.a\[1\] _00714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09826_ _00085_ clknet_leaf_82_wb_clk_i _00002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_100_Left_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09757_ _00020_ clknet_leaf_102_wb_clk_i cpu.regs\[15\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_5_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_5_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06969_ _02552_ _02582_ _02583_ _00064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08708_ _03940_ cpu.ROM_addr_buff\[7\] _03937_ _03941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_69_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09688_ _04800_ _04801_ _04813_ _04814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_107_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08639_ cpu.orig_IO_addr_buff\[5\] _03842_ _03845_ _01733_ _03886_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05512__I cpu.spi.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05116__S0 _00799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07430__A1 cpu.spi.dout\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05992__A1 _00980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_75_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_75_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_113_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07421__A1 cpu.spi.dout\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06224__A2 cpu.spi.divisor\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08889__B _03395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08990_ _00662_ _04195_ _04196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05283__I0 _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07941_ cpu.uart.receive_div_counter\[2\] _03333_ _03335_ _03340_ _03341_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07872_ _03025_ _03289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09611_ _04729_ _04742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08921__A1 _03439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06823_ _02454_ _02436_ _02458_ _00043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09542_ net57 _04689_ _04690_ _04693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06754_ _02401_ _02402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_92_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05705_ _01203_ _01370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06685_ _01919_ _02338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09473_ _00567_ _04627_ _04641_ _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__09232__C _03836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05636_ cpu.C _01302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08424_ _03677_ _03714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05567_ _01232_ _01233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08355_ _03655_ _03656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07306_ _02791_ _02812_ _02820_ _00164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_34_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05498_ _01155_ _01163_ _01164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_46_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08286_ cpu.pwm_top\[1\] _03605_ _03609_ _03610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07237_ _02774_ _00141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07168_ cpu.regs\[11\]\[1\] _02733_ _02735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06119_ cpu.spi.dout\[6\] _01393_ _01218_ _01778_ _01779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__07412__A1 _00748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05274__I0 cpu.regs\[12\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07099_ _01469_ _02686_ _02689_ _00088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_70_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05726__A1 _01390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09809_ _00072_ clknet_leaf_116_wb_clk_i cpu.toggle_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05041__I3 cpu.regs\[11\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06206__A2 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06801__I _02439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08903__A1 cpu.PC\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06142__A1 _00810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06470_ _02122_ _02125_ _02127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05152__I cpu.PORTB_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05421_ _00992_ _01050_ _01087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09559__I _04695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08140_ cpu.toggle_ctr\[12\] _03489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_16_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05352_ _01017_ _01018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07642__A1 _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08071_ _03441_ _03442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05283_ _00925_ _00929_ _00848_ _00952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_3_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07022_ _02467_ _02611_ _02626_ _00074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_24_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06711__I _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08973_ _04138_ _04179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07924_ _03326_ _00276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05708__A1 net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07855_ cpu.uart.data_buff\[1\] _03264_ _03274_ _03275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07786_ cpu.uart.div_counter\[9\] _03215_ _03208_ _03219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06806_ _02441_ _02442_ _02444_ _02445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08638__I _03370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04998_ _00695_ cpu.ROM_spi_mode net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_clkbuf_leaf_28_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09525_ _04680_ _04682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06737_ _02373_ _02385_ _02386_ _00029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_39_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09456_ _00569_ _04592_ _03234_ _04629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06668_ cpu.mem_cycle\[5\] _01909_ _02321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_78_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05619_ _00968_ _01285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_08407_ cpu.timer_capture\[7\] _03652_ _03675_ _03701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_108_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09387_ _04568_ _04571_ _04572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_74_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06599_ _02254_ _02225_ _02255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_22_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05997__I _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08338_ _03635_ _03643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07633__A1 _03088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08269_ cpu.pwm_counter\[5\] _03594_ _03593_ _03597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_116_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10300_ _00558_ clknet_leaf_92_wb_clk_i cpu.regs\[9\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10231_ _00489_ clknet_leaf_62_wb_clk_i cpu.mem_cycle\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__04998__A2 cpu.ROM_spi_mode vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08189__A2 _01723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09418__B _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07236__I1 cpu.regs\[8\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output79_I net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10162_ _00420_ clknet_leaf_27_wb_clk_i cpu.uart.divisor\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05947__A1 _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_67_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10093_ _00352_ clknet_leaf_102_wb_clk_i cpu.pwm_counter\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06777__B _00685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04922__A2 _00621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08113__A2 _03396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06124__A1 cpu.timer_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05970_ cpu.uart.dout\[4\] _01022_ _01589_ _01632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_57_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08727__I1 cpu.ROM_addr_buff\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04921_ net18 _00622_ _00623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07640_ _03091_ _03094_ _03096_ _03056_ _00222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__04986__I _00685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06363__A1 _00783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07571_ cpu.spi.div_counter\[0\] _03044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_0_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09310_ cpu.last_addr\[3\] cpu.ROM_addr_buff\[3\] _04485_ _04505_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06522_ _02168_ _02172_ _02179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_36_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09241_ cpu.orig_PC\[12\] _03863_ _04438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06453_ _02109_ _00812_ _02110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_113_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09172_ _04360_ _04371_ _04372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05404_ _01069_ _01048_ _01070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06384_ _00871_ _02040_ _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_8_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_90_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_90_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_7_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05335_ _00691_ _01000_ _00575_ _01001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_71_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08123_ _02614_ _03474_ _03478_ _00323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08054_ cpu.orig_flags\[2\] _03428_ _03421_ _03429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05266_ cpu.base_address\[4\] _00935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07005_ _02456_ _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_101_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05197_ _00866_ _00868_ _00869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08591__A2 _01618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input30_I sram_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08956_ _04137_ _04135_ _04160_ _04162_ _04163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07907_ cpu.uart.receive_buff\[1\] _03313_ _03316_ cpu.uart.receive_buff\[0\] _03317_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08887_ _00643_ _04095_ _04096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09540__A1 net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07838_ _03250_ _03260_ _03261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09508_ _03823_ _04665_ _04670_ _00516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07769_ _03145_ _03195_ _03190_ _03204_ _03205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09439_ cpu.ROM_spi_dat_out\[3\] _04579_ _04606_ _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07854__A1 _02426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06616__I _00815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10214_ _00472_ clknet_4_13_0_wb_clk_i cpu.PC\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07891__B _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10145_ _00404_ clknet_leaf_15_wb_clk_i cpu.spi.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10076_ _00335_ clknet_leaf_118_wb_clk_i cpu.toggle_ctr\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_4_10_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09531__A1 net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08278__I _03602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05320__A2 _00986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05120_ _00810_ _00811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08741__I _03966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08270__A1 _03588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05051_ _00744_ _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_21_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08810_ _00905_ _04017_ _04021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_5_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09790_ _00053_ clknet_leaf_7_wb_clk_i cpu.timer_capture\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08741_ _03966_ _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05953_ _01615_ _01616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09522__A1 _03833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08672_ _03911_ cpu.ROM_addr_buff\[0\] _03813_ _03912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_04904_ cpu.instr_buff\[15\] _00607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_05884_ net28 _01527_ _01463_ _01547_ _01548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_07623_ _03081_ _03084_ _00217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08089__A1 _03453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07554_ cpu.spi.data_out_buff\[3\] _03016_ _03026_ _03031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07485_ _02951_ _02967_ _02968_ _02969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06505_ _00947_ _02131_ _02039_ _01732_ _02162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_91_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09224_ _04183_ _04409_ _04421_ _04366_ _04422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_8_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06436_ _02090_ _02092_ _02093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_63_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09589__A1 _02538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09155_ _02209_ _04273_ _04355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06367_ _01947_ _01944_ _01731_ _02024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_44_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08106_ cpu.orig_PC\[11\] _03464_ _03467_ _03468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09086_ _00662_ _04288_ _04289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05318_ _00873_ _00985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06298_ _01954_ _01955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08261__A1 _03588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08037_ _03415_ _03413_ _03416_ _00299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05249_ _00918_ _00919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__05614__A3 _01007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_112_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09988_ _00247_ clknet_leaf_25_wb_clk_i cpu.uart.div_counter\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05378__A2 _01006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06575__A1 _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08939_ _04108_ _04134_ _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_67_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08561__I _02443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05369__A2 _01034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10128_ _00387_ clknet_leaf_1_wb_clk_i cpu.timer\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09504__A1 _03815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10059_ _00318_ clknet_leaf_70_wb_clk_i cpu.orig_PC\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_29_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_29_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_89_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07270_ _02796_ _02798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08672__S _03813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06221_ _01878_ _01879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07046__A2 _02441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06152_ _01313_ _01811_ _01812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06083_ _01740_ _00979_ _01744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05103_ _00790_ _00792_ _00794_ _00766_ _00795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_09911_ _00170_ clknet_leaf_87_wb_clk_i cpu.regs\[4\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05034_ cpu.regs\[2\]\[2\] _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_41_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08546__A2 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Left_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09842_ _00101_ clknet_leaf_105_wb_clk_i cpu.regs\[13\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09773_ _00036_ clknet_leaf_52_wb_clk_i cpu.br_rel_dest\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08724_ _03953_ _00449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06985_ _02585_ _02569_ _02598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08849__A3 _00985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05936_ cpu.timer_top\[3\] _01236_ _01598_ _01599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08655_ _02394_ _02850_ _03898_ _02371_ _03899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_05867_ cpu.br_rel_dest\[2\] _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_07606_ cpu.spi.div_counter\[6\] _03071_ _03072_ _03073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_95_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08586_ _03837_ _03838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07537_ cpu.spi.data_out_buff\[0\] _03016_ _02675_ _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05798_ _01462_ _01463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_91_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Left_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05070__I _00763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07468_ cpu.timer\[12\] _02952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09207_ _04299_ _04401_ _04405_ _04406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06419_ _02041_ _02043_ _02076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07399_ _01549_ _02234_ _02892_ _02893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09138_ _04334_ _04337_ _04338_ _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09477__I net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08785__A2 _03970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09069_ _04238_ _04272_ _04210_ _00475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_31_Left_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09734__A1 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output61_I net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06720__A1 _00579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09670__B1 _02465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08473__A1 _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06804__I _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09725__A1 _04043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06770_ _02413_ _02414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05721_ _01385_ _01142_ _01386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08700__A2 cpu.regs\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05652_ _00908_ _01116_ _01318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08440_ cpu.timer_capture\[13\] _03652_ _03727_ _03728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08371_ _02977_ _03658_ _02980_ _03670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05583_ _01248_ _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07267__A2 _02777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07322_ _02785_ _02826_ _02831_ _00169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08464__A1 _02480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06475__B1 _02040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07253_ cpu.regs\[7\]\[2\] _02786_ _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06204_ _01457_ _01861_ _01862_ _01332_ _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07184_ _02684_ _02729_ _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06227__B1 _01390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06135_ _01058_ _01155_ _01794_ _01795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06778__A1 _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06066_ _01277_ _01693_ _01726_ _01521_ _01727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_111_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09716__A1 _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05017_ _00003_ _00713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09825_ _00084_ clknet_leaf_100_wb_clk_i _00001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09756_ _00019_ clknet_leaf_106_wb_clk_i cpu.regs\[15\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06968_ _02186_ _02567_ _02583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06950__A1 _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08707_ _02597_ _03933_ _03939_ _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05919_ _01186_ _01580_ _01581_ _01582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09687_ _04024_ _04812_ _04169_ _01937_ _04813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08638_ _03370_ _03885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06899_ _02403_ _02523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_107_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08569_ _03796_ _03817_ _03825_ _00422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_36_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05269__A1 _00006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09000__I _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05116__S1 _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06941__A1 _02556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07249__A2 _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08446__A1 _03681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08749__A2 _03970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_7_0_wb_clk_i clknet_0_wb_clk_i clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07940_ cpu.uart.receive_div_counter\[2\] cpu.uart.receive_div_counter\[1\] cpu.uart.receive_div_counter\[0\]
+ _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
Xclkbuf_leaf_44_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_44_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07871_ _03269_ _03288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09610_ cpu.ROM_addr_buff\[4\] _02355_ _02356_ cpu.ROM_addr_buff\[8\] cpu.ROM_addr_buff\[12\]
+ _02340_ _04741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_06822_ cpu.uart.divisor\[4\] _02437_ _02457_ _02458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09541_ _03801_ _04688_ _04692_ _00527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06753_ _02400_ _02401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05704_ net22 _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06684_ _01912_ _01915_ _02337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09472_ _04630_ _00570_ _04640_ _04641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05043__S0 _00716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05635_ _01279_ _01283_ _01300_ _01301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08423_ _03713_ _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05566_ _01026_ _01225_ _01232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08354_ _03654_ _02997_ _03655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07305_ cpu.regs\[5\]\[5\] _02815_ _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05497_ _01139_ _01159_ _01162_ _01096_ _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_61_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08285_ _03608_ _03609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07236_ _02756_ cpu.regs\[8\]\[6\] _02764_ _02774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07167_ _02710_ _02732_ _02734_ _00111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06118_ _01775_ _01776_ _01777_ _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05274__I1 cpu.regs\[13\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07098_ cpu.regs\[14\]\[1\] _02687_ _02689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06049_ cpu.spi.dout\[5\] _01393_ _01218_ _01709_ _01710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_10_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09808_ _00071_ clknet_leaf_116_wb_clk_i cpu.toggle_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05726__A2 _00999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09739_ _04837_ _04852_ _04853_ _00564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_4_15_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08428__A1 cpu.timer_capture\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_96_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08600__A1 _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07913__I _03213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08667__A1 _02388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06529__I _02009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05025__S0 _00697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08744__I _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05420_ _01083_ _01085_ _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07788__C _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05351_ _01014_ _01016_ _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09092__A1 _00798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07642__A2 _03094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05282_ _00936_ _00950_ _00951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08070_ cpu.PC\[2\] _03441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05653__A1 _00908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07021_ _01842_ _02621_ _02623_ _02626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08972_ _04177_ _04178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07923_ cpu.uart.receive_buff\[7\] _03313_ _03314_ net15 _02439_ _03326_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_07854_ _02426_ _03260_ _03274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06805_ _02443_ _02434_ _02444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07785_ _03215_ _03208_ _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04997_ net75 _00695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06381__A2 cpu.multiplier.a\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09524_ _04680_ _04681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06736_ _00673_ _02377_ _02379_ _02386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08658__A1 _00984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06667_ _02317_ _02318_ _02319_ _02320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_09455_ _04627_ _04628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_94_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05618_ _00965_ _01284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_19_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08406_ _02514_ _03692_ _03657_ _03699_ _03700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06133__A2 _01761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09386_ _04570_ _04571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06598_ cpu.PC\[13\] _02254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XTAP_TAPCELL_ROW_50_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05892__A1 _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05549_ cpu.uart.busy _01135_ _01134_ _01215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_74_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09083__A1 _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08337_ _02450_ _03636_ _03642_ _03641_ _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08268_ _03594_ _03593_ cpu.pwm_counter\[5\] _03596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08830__A1 _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07219_ _02711_ _02729_ _02763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10230_ _00488_ clknet_leaf_56_wb_clk_i cpu.mem_cycle\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08199_ _03531_ _03547_ _03548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_115_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06902__I _02443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Left_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07397__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10161_ _00419_ clknet_leaf_27_wb_clk_i cpu.uart.divisor\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10092_ _00351_ clknet_leaf_103_wb_clk_i cpu.pwm_counter\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08897__A1 _04103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08649__B2 _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07321__A1 cpu.regs\[4\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09074__A1 cpu.PC\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09328__C _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09129__A2 _04244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04920_ _00581_ _00622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07560__A1 _02508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07570_ _02914_ _03043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_69_Left_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05163__I _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06521_ _02154_ _02175_ _02177_ _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_87_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09240_ _04436_ _04437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07312__A1 _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06452_ _00915_ _02072_ _02039_ _00954_ _02109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09171_ _04248_ _04367_ _04370_ _04371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05403_ cpu.IO_addr_buff\[3\] _01069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_56_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06383_ _02039_ _02040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05334_ cpu.ROM_spi_cycle\[4\] cpu.ROM_spi_cycle\[1\] cpu.ROM_spi_cycle\[0\] _00570_
+ _01000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_0_44_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08122_ _01417_ _03475_ _03477_ _03478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08053_ _03407_ _03428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_78_Left_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05265_ _00934_ net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07004_ _02610_ _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06722__I _00579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05196_ _00833_ _00867_ _00849_ _00868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_08955_ _04161_ _04162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06051__A1 cpu.timer_capture\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07906_ _03315_ _03316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input23_I io_in[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08886_ _00671_ _04094_ _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_79_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07837_ _03176_ _03260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07768_ _03145_ _03201_ _03204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09507_ net61 _04666_ _04667_ _04670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06719_ _02369_ _02370_ _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_07699_ _02648_ _03144_ _03145_ _02633_ _03147_ _03148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_66_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09438_ _04615_ _00501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_109_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09369_ _04554_ _04557_ _02524_ _00490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08803__A1 _03403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09429__B _04603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output91_I net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10213_ _00471_ clknet_leaf_55_wb_clk_i cpu.PC\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06042__A1 _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10144_ _00403_ clknet_leaf_12_wb_clk_i cpu.spi.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09164__B _04108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10075_ _00334_ clknet_leaf_119_wb_clk_i cpu.toggle_ctr\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07542__A1 _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06079__I _00796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_qcpu_110 io_out[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_58_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05608__A1 _00636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05050_ cpu.multiplier.a\[3\] _00744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08022__A2 _03404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05158__I _00006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08740_ _02366_ _03965_ _03966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__04997__I net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05952_ _01614_ _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08671_ _03433_ _00649_ _03910_ _03911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04903_ _00605_ _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05883_ _01436_ _00742_ _01546_ _01547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07622_ cpu.spi.data_in_buff\[2\] _03083_ _03078_ cpu.spi.data_in_buff\[3\] _03084_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_88_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07553_ cpu.spi.data_out_buff\[4\] _03021_ _03029_ _03030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_101_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07484_ _02946_ cpu.timer\[15\] cpu.timer\[14\] _02948_ _02968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06504_ _02105_ _00955_ _02161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09223_ _04417_ _04419_ _04420_ _04421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06435_ _00812_ _02091_ _02092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_33_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_86_Left_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09154_ _04326_ _04354_ _04324_ _00478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06880__C _02506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06366_ _00946_ _01731_ _01946_ _02023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08105_ _03456_ _03467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09085_ _02421_ _04188_ _04287_ _04194_ _04288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05317_ _00983_ _00984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06297_ cpu.multiplier.a\[1\] _00727_ _01954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08036_ cpu.orig_IO_addr_buff\[5\] _03408_ _03411_ _03416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05248_ _00917_ _00918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_112_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05179_ cpu.regs\[8\]\[1\] cpu.regs\[9\]\[1\] cpu.regs\[10\]\[1\] cpu.regs\[11\]\[1\]
+ _00836_ _00839_ _00851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XPHY_EDGE_ROW_95_Left_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09987_ _00246_ clknet_leaf_29_wb_clk_i cpu.uart.div_counter\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08938_ _04141_ _04144_ _04145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08869_ _00607_ _00673_ _01160_ _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__07524__A1 _00694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09277__B2 _04162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09029__A1 _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08252__A2 _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05369__A3 _01007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10127_ _00386_ clknet_leaf_1_wb_clk_i cpu.timer\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10058_ _00317_ clknet_leaf_70_wb_clk_i cpu.orig_PC\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07515__A1 _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05621__S0 _01285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_69_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_69_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06220_ cpu.spi.div_counter\[2\] _01878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_70_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08752__I _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06151_ _01810_ _01804_ _01811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_5_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06082_ _01740_ _00980_ _01743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05102_ _00790_ _00793_ _00794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09910_ _00169_ clknet_leaf_89_wb_clk_i cpu.regs\[4\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05033_ _00727_ _00728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09841_ _00100_ clknet_leaf_96_wb_clk_i cpu.regs\[13\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06984_ _02596_ _02597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_09772_ _00035_ clknet_leaf_98_wb_clk_i cpu.br_rel_dest\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08723_ _03951_ cpu.ROM_addr_buff\[10\] _03952_ _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05935_ _01410_ _01598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05080__I2 cpu.regs\[6\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08849__A4 _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08654_ _02398_ _02850_ _03898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05866_ _01529_ _01440_ _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07605_ cpu.spi.div_counter\[6\] _03050_ _03066_ _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08585_ _00658_ _03837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05797_ _01312_ _01309_ _01462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07109__I1 _01815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07536_ _03010_ _03016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09206_ _04374_ _04383_ _04403_ _04404_ _04321_ _04405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_64_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07467_ _02948_ cpu.timer\[14\] _02950_ _02951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06418_ _02064_ _02068_ _02074_ _02075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_07398_ _02259_ _02891_ _02892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09137_ _04334_ _04337_ _04183_ _04338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06349_ _01979_ _01984_ _02006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09068_ _04175_ _04266_ _04271_ _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08019_ _03403_ _03404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_20_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06910__I _02523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08330__C _02542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05287__A2 _00955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06092__I _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_116_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_116_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06820__I _02455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08747__I _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05720_ cpu.uart.dout\[1\] _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05651_ _01302_ cpu.base_address\[0\] _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08370_ _02996_ _03667_ _03668_ _03669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05582_ _01027_ _01073_ _01248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07321_ cpu.regs\[4\]\[2\] _02830_ _02831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07600__B _00645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07252_ _02778_ _02786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06475__A1 _00955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06203_ _00826_ _01759_ _01862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_07183_ _02742_ _02733_ _02743_ _00118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06134_ _01733_ _01521_ _01655_ _01793_ _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_6_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06065_ _01471_ _01725_ _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_47_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05016_ _00712_ net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_10_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09824_ _00083_ clknet_leaf_99_wb_clk_i _00000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05202__A2 _00873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09755_ _00018_ clknet_leaf_101_wb_clk_i cpu.regs\[15\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06967_ _01751_ _02581_ _02553_ _02582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05918_ net9 _01204_ _01581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08706_ _03926_ cpu.regs\[2\]\[7\] _03939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08657__I _03899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09686_ net97 _02465_ _04802_ _04810_ _04811_ _04812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_06898_ cpu.timer_top\[0\] _02521_ _02522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08637_ _03860_ _03884_ _00431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05849_ _01512_ _01258_ _01126_ _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08568_ cpu.uart.divisor\[11\] _03818_ _03821_ _03825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07519_ _01898_ _01901_ _03002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_77_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08499_ _02430_ _01040_ _01004_ _00999_ _03776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XTAP_TAPCELL_ROW_40_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_86_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_48_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07471__I cpu.timer_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07709__A1 _00621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07870_ cpu.uart.data_buff\[4\] _03282_ _03286_ _03287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05166__I _00837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06821_ _02456_ _02457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09540_ net56 _04689_ _04690_ _04692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06752_ _02394_ _02397_ _02399_ _02371_ _02400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XPHY_EDGE_ROW_50_Left_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_84_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_84_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09471_ _04631_ _04632_ _00568_ _04640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_92_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05703_ _01055_ _01367_ _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_13_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_13_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08134__A1 _02460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06683_ _02334_ _02335_ _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08422_ cpu.timer_capture\[10\] _03678_ _03712_ _03690_ _03713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05634_ _01283_ _01297_ _01299_ _01300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05043__S1 _00717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05565_ cpu.timer_capture\[8\] _01231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08353_ _02944_ _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__06725__I _02372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07304_ _02819_ _00163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08284_ _03607_ _03608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05496_ _01160_ _00935_ _01161_ _01162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_46_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07235_ _02725_ _02766_ _02773_ _00140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_81_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07166_ cpu.regs\[11\]\[0\] _02733_ _02734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_3_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06117_ cpu.spi.divisor\[6\] _01179_ _01176_ _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07097_ _01353_ _02686_ _02688_ _00087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06048_ _01706_ _01707_ _01708_ _01709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05274__I2 cpu.regs\[14\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08373__A1 cpu.timer_capture\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07999_ _03371_ _03387_ _00290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_70_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09807_ _00070_ clknet_leaf_115_wb_clk_i cpu.toggle_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__04934__A1 cpu.uart.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05726__A3 _01126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09738_ _00728_ _04837_ _04853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08125__A1 _02447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05804__I _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09669_ _01266_ _01263_ _03843_ _01041_ _04050_ _04795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__09625__A1 _03618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05695__B net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05178__A1 _00843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08116__A1 _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05025__S1 _00698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05350_ _01015_ _01016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_112_Right_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05281_ _00949_ _00950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05653__A2 _00870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07020_ _02463_ _02611_ _02625_ _00073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_101_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06602__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08971_ _04173_ _04132_ _04177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07922_ _03320_ _03325_ _00275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07853_ _03266_ _03273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06804_ _01450_ _02443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04996_ _00624_ _00688_ _00632_ _00690_ _00694_ _00009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_07784_ _03214_ _03217_ _00245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09523_ _01028_ _04663_ _04680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06735_ _02384_ _02385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_104_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06666_ _01917_ _01919_ _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_09454_ _00569_ _04592_ _04627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09385_ _04548_ _04543_ _02307_ _04570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05617_ _01282_ _01283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08405_ _03697_ _03698_ _03699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_52_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08336_ cpu.timer_top\[11\] _03637_ _03642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06597_ net116 _02252_ _02253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05548_ cpu.uart.dout\[0\] _01023_ _00993_ _01213_ _01214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_62_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05479_ _00654_ _01119_ _01124_ _01144_ _01145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_61_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08267_ _03585_ _03595_ _00350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08830__A2 _00728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08198_ _03513_ _03546_ _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07218_ _01869_ _02762_ _00134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07149_ _01615_ _02722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_115_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07286__I _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10160_ _00012_ clknet_leaf_17_wb_clk_i cpu.uart.clr_hb vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08594__B2 _00986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10091_ _00350_ clknet_leaf_11_wb_clk_i cpu.pwm_counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_76_Right_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_58_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_106_Left_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_83_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09074__A2 _00636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07085__A1 _02677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_85_Right_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_94_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_115_Left_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10289_ _00547_ clknet_leaf_62_wb_clk_i net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XPHY_EDGE_ROW_94_Right_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05444__I _00652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06520_ _02157_ _02176_ _02177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_88_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07312__A2 _02777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06451_ _02083_ _02087_ _02107_ _02108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05402_ _00596_ _01068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09170_ _03903_ _04256_ _04369_ _04262_ _04370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06382_ _02038_ _02039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05333_ _00998_ _00999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_44_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08121_ _03456_ _03477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08052_ cpu.IE _03427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06823__A1 _02454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05264_ _00911_ _00922_ _00933_ _00934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__05626__A2 _01291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07003_ _02443_ _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05195_ cpu.regs\[8\]\[0\] cpu.regs\[9\]\[0\] cpu.regs\[10\]\[0\] cpu.regs\[11\]\[0\]
+ _00858_ _00859_ _00867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_08954_ _00678_ _00669_ _04161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07905_ _03307_ _03314_ _03315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08885_ _00666_ _04090_ _04093_ _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07836_ _03252_ _03154_ _03259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input16_I io_in[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07767_ _03133_ _03197_ _03203_ _03113_ _00242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_04979_ _00678_ _00679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09506_ _03820_ _04665_ _04669_ _00515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06718_ _02332_ _02367_ _02370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07698_ _03146_ _02631_ _02441_ _03136_ _03147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_09437_ cpu.ROM_spi_dat_out\[3\] _04609_ _04614_ _04527_ _04615_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_109_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06649_ cpu.startup_cycle\[6\] _02299_ _02301_ _02302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_63_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09368_ _04544_ _04556_ _04557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05303__B _00845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09299_ cpu.last_addr\[11\] _04490_ _04494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08319_ cpu.timer_div_counter\[5\] _03628_ _03631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08567__A1 _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10212_ _00470_ clknet_leaf_54_wb_clk_i cpu.PC\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10143_ _00402_ clknet_leaf_15_wb_clk_i cpu.spi.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10074_ _00333_ clknet_leaf_119_wb_clk_i cpu.toggle_ctr\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08575__I _03829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_qcpu_100 io_oeb[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_69_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_qcpu_111 io_oeb[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_84_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06805__A1 _02443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05608__A2 _01273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input8_I io_in[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05951_ _01613_ _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08670_ _03909_ _00696_ _03910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04902_ _00604_ _00605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05882_ _01536_ _01539_ _01545_ _01546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07621_ _01893_ _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08730__A1 _03469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07552_ _02495_ _03022_ _03029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06503_ _02158_ _02159_ _02160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07483_ _02954_ _02964_ _02966_ _02967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09222_ _04417_ _04419_ _04107_ _04420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_60_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06434_ _00854_ _02072_ _02039_ _00915_ _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09153_ _04299_ _04349_ _04353_ _04354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06365_ _00746_ _02021_ _02022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08104_ cpu.PC\[11\] _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_05316_ _00856_ _00983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09084_ _04189_ _04275_ _04286_ _04260_ _04287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_71_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06296_ _01952_ _01945_ _00916_ _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08035_ cpu.IO_addr_buff\[5\] _03415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05247_ _00916_ _00917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05178_ _00843_ _00847_ _00849_ _00850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_40_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09986_ _00245_ clknet_leaf_29_wb_clk_i cpu.uart.div_counter\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_4_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08937_ _04142_ _04143_ _04144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08868_ cpu.orig_PC\[0\] _04075_ _04076_ _04077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07819_ _03243_ _03245_ _00252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_67_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08799_ _01041_ _03843_ _04011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07288__A1 _02807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06129__B _01137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08788__A1 _00686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06015__A2 _01676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07474__I cpu.timer_top\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05774__A1 _00711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10126_ _00385_ clknet_leaf_5_wb_clk_i cpu.timer\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10057_ _00316_ clknet_leaf_70_wb_clk_i cpu.orig_PC\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08712__A1 _02856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07515__A2 _02998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09268__A2 _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05621__S1 _01286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_38_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_38_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_81_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06150_ _01537_ _01807_ _01809_ _00811_ _01810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_110_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06081_ _00980_ _01451_ _01741_ _01453_ _01454_ _01742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05101_ cpu.regs\[12\]\[5\] cpu.regs\[13\]\[5\] cpu.regs\[14\]\[5\] cpu.regs\[15\]\[5\]
+ _00770_ _00771_ _00793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_clkbuf_leaf_37_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05032_ cpu.multiplier.a\[2\] _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09840_ _00099_ clknet_leaf_104_wb_clk_i cpu.regs\[13\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06983_ _02212_ _02596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09771_ _00034_ clknet_leaf_81_wb_clk_i cpu.br_rel_dest\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08722_ _03812_ _03952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05934_ cpu.timer_capture\[11\] _01227_ _01596_ _01032_ _01597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_89_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08653_ _03885_ _03897_ _00434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05865_ _01444_ _01529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07604_ _03038_ _02910_ _01902_ _03070_ _03071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_88_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08584_ _03835_ _03836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05796_ _01316_ _01445_ _01455_ _01460_ _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_07535_ cpu.spi.data_out_buff\[1\] _03007_ _03014_ _03015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07466_ cpu.timer_top\[13\] _02949_ _02950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09205_ _04034_ _04404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_63_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06417_ _00812_ _02073_ _02074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_17_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_76_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07397_ net19 _02855_ _02890_ _02891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_71_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09136_ _04335_ _04336_ _04337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06348_ _01986_ _02004_ _02005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_17_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05128__S0 _00816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09067_ _04267_ _04242_ _04270_ _04235_ _04207_ _04271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06279_ _01935_ _01936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08018_ _03400_ _03403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09969_ _00228_ clknet_leaf_38_wb_clk_i cpu.uart.dout\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09498__A2 _02432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output47_I net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07681__B2 _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08933__A1 cpu.PC\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10109_ _00368_ clknet_leaf_8_wb_clk_i cpu.timer_div_counter\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05880__C _01434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05650_ _00877_ _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08161__A2 cpu.toggle_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_110_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05581_ _01242_ _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09110__A1 _02423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07320_ _02824_ _02830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08763__I _02404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07251_ _01550_ _02785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06202_ _00827_ _01760_ _01861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07182_ cpu.regs\[11\]\[7\] _02736_ _02743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06227__A2 cpu.spi.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06133_ _01277_ _01761_ _01792_ _01518_ _01793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_14_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08712__B _03943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06064_ _01694_ _01516_ _01722_ _01724_ _01725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__09177__A1 _04374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05015_ _00711_ _00712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09823_ _00082_ clknet_leaf_32_wb_clk_i cpu.uart.receive_counter\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05038__I0 cpu.regs\[4\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09754_ _00017_ clknet_leaf_105_wb_clk_i cpu.regs\[15\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06966_ _02575_ _02580_ _02581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08705_ _03938_ _00445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05917_ _01122_ _01578_ _01579_ _01053_ _01580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06886__C _02506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09685_ _00811_ _01808_ _01862_ _04811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06897_ _02519_ _02521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_96_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06163__A1 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08636_ cpu.IO_addr_buff\[4\] _03861_ _03882_ _03883_ _03884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_55_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08152__A2 _01512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05848_ cpu.toggle_top\[10\] _01512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_77_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08567_ _03823_ _03817_ _03824_ _00421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05779_ net91 _01443_ _01444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_37_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07518_ _00692_ _03001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08498_ _03760_ _03773_ _03775_ _00401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_40_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07449_ cpu.timer_div_counter\[1\] _02933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_52_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09119_ _02429_ _04321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_75_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09437__C _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09168__A1 _03848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05901__A1 _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08906__A1 _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06820_ _02455_ _02456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05196__A2 _00867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06751_ _02398_ _02397_ _02399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09706__I0 _02818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06682_ _02331_ _02322_ _02335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09470_ _04631_ _04637_ _00567_ _04639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05702_ net60 _01195_ _01367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06145__A1 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08421_ _02989_ _03679_ _03680_ _03711_ _03684_ _03712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_106_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05633_ _01298_ _01299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_53_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_53_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_74_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05564_ _01219_ _01223_ _01228_ _01229_ _01230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05910__I _01108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08352_ _03652_ _03653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05495_ _00607_ _00672_ _01161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08283_ _00619_ _03607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07303_ _02818_ cpu.regs\[5\]\[4\] _02810_ _02819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07234_ cpu.regs\[8\]\[5\] _02769_ _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07165_ _02731_ _02733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06116_ cpu.uart.dout\[6\] _01022_ _01588_ _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07096_ cpu.regs\[14\]\[0\] _02687_ _02688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06047_ cpu.spi.divisor\[5\] _01180_ _01181_ _01708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05274__I3 cpu.regs\[15\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_109_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07998_ cpu.uart.receive_div_counter\[13\] _03345_ _03384_ _03386_ _03387_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08668__I _00648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09806_ _00069_ clknet_leaf_116_wb_clk_i cpu.toggle_top\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06949_ _02555_ _02564_ _02565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09737_ _01549_ _02555_ _04851_ _04852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__04934__A2 cpu.spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09668_ cpu.orig_flags\[0\] _04244_ _04789_ _04793_ _04794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09599_ _02325_ _01911_ _02322_ _04730_ _04731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_96_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07884__A1 _02508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08619_ _03835_ _03870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09448__B _04603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05178__A2 _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08116__A2 _02433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06098__I _01757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07175__I0 _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06127__A1 cpu.pwm_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05280_ _00948_ _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_3_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06602__A2 _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08970_ _04101_ _04176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_100_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_100_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07921_ cpu.uart.receive_buff\[7\] _03321_ _03315_ cpu.uart.receive_buff\[6\] _03325_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09552__A1 cpu.PORTB_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07852_ _03272_ _00258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput1 io_in[0] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_06803_ _02434_ _02442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09522_ _03833_ _04672_ _04679_ _00521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09304__A1 cpu.last_addr\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04995_ _00693_ _00694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07783_ _03215_ _03209_ _03216_ _03208_ _03217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06734_ net19 _02374_ _02384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09453_ _04626_ _00505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06665_ _01908_ _01909_ _02318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_93_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09384_ _04556_ _04553_ _04569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05616_ _01281_ _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08404_ cpu.timer\[7\] cpu.timer\[6\] _03693_ _03698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_93_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05341__A2 _01006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08335_ _02527_ _03636_ _03640_ _03641_ _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06596_ _02242_ _02251_ _02252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_117_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05547_ _01010_ _01213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05478_ _01132_ _01134_ _01136_ _01143_ _01144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__08291__A1 _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08266_ _03594_ _03593_ _03595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08197_ _03516_ _03545_ _03546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07217_ _01796_ _01813_ _02762_ _00133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07148_ _02719_ _02714_ _02721_ _00105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_115_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07079_ _02673_ _02674_ _02676_ _00081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10090_ _00349_ clknet_leaf_102_wb_clk_i cpu.pwm_counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09543__A1 _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06109__A1 net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07157__I0 _01816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08282__A1 _02427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_94_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10288_ _00546_ clknet_leaf_63_wb_clk_i cpu.ROM_spi_mode vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09534__A1 _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08101__I _03400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06450_ _01951_ _01757_ _02085_ _02033_ _02107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_118_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05401_ _00590_ _00597_ _01066_ _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_7_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06381_ _00781_ cpu.multiplier.a\[6\] _02038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05332_ _00989_ _00997_ _00998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08120_ _02427_ _03474_ _03476_ _00322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08273__A1 _02478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08051_ _03425_ _03423_ _03426_ _00303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05263_ _00932_ _00933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_43_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07002_ _02608_ _02611_ _02613_ _02542_ _00067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_12_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05194_ _00857_ _00865_ _00866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__06587__A1 _00815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08953_ _04156_ _04159_ _04160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07904_ _02666_ _03311_ _03306_ _03314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08884_ _04042_ _04091_ _04092_ _00665_ _04093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07835_ _03258_ _00255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07766_ cpu.uart.div_counter\[5\] _03184_ _03202_ _03203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_04978_ cpu.instr_buff\[15\] _00678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09505_ net60 _04666_ _04667_ _04669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06717_ _02366_ _02368_ _02369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_79_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07071__B _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09436_ _04594_ _04613_ _04614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07697_ cpu.uart.div_counter\[7\] _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_94_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06648_ _02300_ _02301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_63_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05370__I _00655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09367_ _04555_ _04556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_81_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06579_ _00784_ _01927_ _02234_ _01932_ _02235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_09298_ cpu.ROM_addr_buff\[13\] _04492_ _04493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_74_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08318_ cpu.timer_div_counter\[5\] _03628_ _03630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_34_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08264__A1 _03588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08249_ _03583_ _00344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10211_ _00469_ clknet_leaf_79_wb_clk_i cpu.Z vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10142_ _00401_ clknet_leaf_4_wb_clk_i cpu.timer_capture\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09516__A1 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10073_ _00332_ clknet_leaf_119_wb_clk_i cpu.toggle_ctr\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_qcpu_101 io_oeb[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_97_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_qcpu_112 io_oeb[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__05280__I _00948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06502__A1 _02119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08524__C _03648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06281__A3 _00674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07000__I _02610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06569__A1 _02203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09507__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05950_ _01571_ _01572_ _01612_ _01613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_108_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04901_ cpu.br_rel_dest\[4\] _00603_ _00604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05881_ _01337_ _01540_ _01542_ _01543_ _01544_ _01545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_07620_ _03081_ _03082_ _00216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_108_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07551_ _03010_ _03028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06502_ _02119_ _00917_ _02136_ _02159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07482_ cpu.timer_top\[12\] _02965_ _02949_ cpu.timer_top\[13\] _02966_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_33_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_66_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09221_ _04386_ _04418_ _04419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_60_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06433_ _02061_ _02058_ _02090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09152_ _04267_ _04329_ _04350_ _04352_ _04321_ _04353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06364_ _00914_ _01993_ _01995_ _00953_ _02021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08103_ _03463_ _03459_ _03465_ _00316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05315_ _00982_ net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08434__C _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09083_ _02585_ _04190_ _04286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06295_ _01951_ _01952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08034_ _00592_ _03413_ _03414_ _00298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05246_ _00915_ _00916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05480__A1 _01116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05177_ _00848_ _00849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_112_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09985_ _00244_ clknet_leaf_28_wb_clk_i cpu.uart.div_counter\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08936_ cpu.PC\[2\] cpu.br_rel_dest\[2\] _04143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06980__A1 _01815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08867_ _04069_ _04075_ _04076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07818_ cpu.uart.div_counter\[15\] _03239_ _03244_ _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08182__B1 cpu.toggle_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08798_ _04009_ _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06732__A1 _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_8_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_8_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07749_ cpu.uart.div_counter\[1\] _03137_ _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09419_ _04595_ _04597_ _04599_ _00498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_66_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06799__A1 _02427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09456__B _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08360__B _03615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10125_ _00384_ clknet_leaf_6_wb_clk_i cpu.timer\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10056_ _00315_ clknet_leaf_70_wb_clk_i cpu.orig_PC\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_89_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06723__A1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05082__S0 _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_100_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08535__B _03774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06080_ _01740_ _00979_ _01741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05100_ _00791_ _00792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_111_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_78_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_78_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05031_ _00726_ net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07665__I net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05214__A1 _00882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_107_Right_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09770_ _00033_ clknet_leaf_81_wb_clk_i cpu.br_rel_dest\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06982_ _02552_ _02594_ _02595_ _00065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08721_ _03463_ _03949_ _03950_ _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05933_ _01593_ _01594_ _01595_ _01596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08652_ cpu.IO_addr_buff\[7\] _03858_ _03896_ _03883_ _03897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08496__I _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07603_ _03069_ _03070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_89_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05864_ net91 _01443_ _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_95_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08583_ _01093_ _03835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05795_ _01457_ _01458_ _01459_ _01332_ _01460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07534_ _02480_ _03008_ _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07465_ cpu.timer\[13\] _02949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09204_ _00729_ _04167_ _04402_ _04403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06416_ net127 _02072_ _02038_ _00854_ _02073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_17_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07396_ _02884_ _02889_ _02851_ _02890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_72_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09135_ _04325_ _00856_ _04336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06347_ _01997_ _02000_ _02003_ _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__05128__S1 _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09066_ _02186_ _04232_ _04269_ _04270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06278_ _01930_ _01935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08017_ _03401_ _03402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05229_ cpu.regs\[12\]\[2\] cpu.regs\[13\]\[2\] cpu.regs\[14\]\[2\] cpu.regs\[15\]\[2\]
+ _00898_ _00899_ _00900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_09968_ _00227_ clknet_leaf_34_wb_clk_i cpu.uart.dout\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08919_ _00643_ _04126_ _04127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09899_ _00158_ clknet_leaf_90_wb_clk_i cpu.regs\[6\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09030__I _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08630__B2 _03870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08933__A2 _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10108_ _00367_ clknet_leaf_20_wb_clk_i cpu.timer_div_counter\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09205__I _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10039_ _00298_ clknet_leaf_51_wb_clk_i cpu.orig_IO_addr_buff\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05580_ _01230_ _01238_ _01245_ _01246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_105_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07250_ _02783_ _02780_ _02784_ _00144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06201_ _01760_ _01343_ _01859_ _01453_ _01435_ _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_07181_ _01868_ _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06132_ _01790_ _01791_ _01270_ _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06063_ _01723_ _01173_ _01137_ _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05014_ _00003_ _00701_ _00710_ _00711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_09822_ _00081_ clknet_leaf_34_wb_clk_i cpu.uart.receive_counter\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09753_ _00016_ clknet_leaf_106_wb_clk_i cpu.regs\[15\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08704_ _03935_ _03936_ _03937_ _03938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06965_ _02237_ _02577_ _02578_ _02579_ _02580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05916_ net24 _01199_ _01579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09684_ _01740_ _01733_ _04031_ _04808_ _04809_ _04810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_06896_ _02519_ _02520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_68_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08635_ _03835_ _03883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05847_ _01508_ _01509_ _01510_ _01511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08566_ _02640_ _03818_ _03821_ _03824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06163__A2 _01018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07517_ net70 _03000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05778_ _01325_ _00855_ _01441_ _01442_ _01443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_71_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08497_ cpu.timer_capture\[15\] _03764_ _03774_ _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_40_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07448_ cpu.timer_div\[3\] cpu.timer_div_counter\[3\] _02932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06474__I _02072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07379_ _02104_ _02126_ _02874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_45_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09118_ _02271_ _04232_ _04319_ _04320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_75_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05426__A1 _01012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09049_ _04138_ _04241_ _04253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06926__A1 _02540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06154__A2 _01813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08851__B2 _01761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05665__A1 _00882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_97_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08603__A1 _03854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07406__A2 _02223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09159__A2 _04244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06750_ _02333_ _02398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_92_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06681_ _01039_ _02334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05701_ _01362_ _01365_ _01018_ _01366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05632_ _01044_ _01298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08420_ _02959_ _03710_ _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07342__A1 cpu.regs\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08774__I _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05563_ cpu.timer_capture\[0\] _01223_ _01229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08351_ _03651_ _03652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07645__A2 _03094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05494_ cpu.base_address\[5\] _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_58_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08842__A1 _02070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06294__I _01950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08282_ _02427_ _03604_ _03606_ _00354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_34_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07302_ _01677_ _02818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07233_ _02772_ _00139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_93_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_93_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_104_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_22_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_22_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07164_ _02731_ _02732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06115_ _01770_ _01772_ _01774_ _01775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07095_ _02685_ _02687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06046_ cpu.uart.dout\[5\] _01023_ _01589_ _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06081__A1 _00980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07997_ _03352_ _03385_ _03386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_70_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06384__A2 _02040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09805_ _00068_ clknet_leaf_115_wb_clk_i cpu.toggle_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06948_ _02257_ _02557_ _02563_ _02564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09736_ _02584_ _04850_ _04851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09667_ _02070_ _04048_ _04051_ _04792_ _04793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_96_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08618_ _03862_ _03866_ _03868_ _03869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06879_ _02483_ _02506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07333__A1 _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09598_ _04729_ _02398_ _04730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08549_ _02333_ _02369_ _03810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09389__A2 _04571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09010__A1 cpu.PC\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07572__A1 _01897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05258__S0 _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08808__B _03395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07175__I1 cpu.regs\[11\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09077__A1 _03453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05638__A1 _01012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07003__I _02443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06842__I _02470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06063__B _01137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06063__A1 _01723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07920_ _03320_ _03324_ _00274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07851_ _02677_ _03271_ _03272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xinput2 io_in[10] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06802_ cpu.uart.divisor\[1\] _02441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07782_ _03215_ _03210_ _03216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09521_ net67 _04673_ _04675_ _04679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04994_ _00692_ _00693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06733_ _02373_ _02382_ _02383_ _00028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_36_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09452_ cpu.ROM_spi_dat_out\[7\] _04609_ _04625_ _00628_ _04626_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06664_ _02316_ _02317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09383_ _02301_ _04568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05615_ _01036_ _01280_ _01281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06595_ _02244_ _02250_ _02251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08403_ _02509_ _03693_ _02514_ _03697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05546_ _01206_ _01208_ _01211_ _00616_ _01212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_47_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08334_ _02523_ _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_62_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05477_ _01137_ _01138_ _01142_ _01143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08265_ cpu.pwm_counter\[4\] _03594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08196_ _03542_ _03544_ _03520_ _03545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07216_ _01753_ _02762_ _00132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_70_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07147_ cpu.regs\[12\]\[2\] _02720_ _02721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05101__I0 cpu.regs\[12\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07078_ _02673_ _02674_ _02675_ _02676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06029_ _01687_ _01689_ _01690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_58_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09719_ _04042_ _04833_ _04835_ _04836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_2_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07157__I1 cpu.regs\[12\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05168__I0 cpu.regs\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_6_0_wb_clk_i clknet_0_wb_clk_i clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_96_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09059__A1 _02419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08806__A1 _00933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09231__A1 _00680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_17_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10287_ _00545_ clknet_leaf_99_wb_clk_i cpu.PORTA_DDR\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_29_Left_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07545__A1 _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05859__A1 cpu.IE vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_1_Left_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_56_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05400_ _01064_ _01065_ _01066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XPHY_EDGE_ROW_38_Left_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06380_ _02032_ net120 _02037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_7_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09369__B _02524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05331_ _00996_ _00997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08050_ cpu.orig_flags\[1\] _03418_ _03421_ _03426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05262_ _00931_ _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_31_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07001_ _00986_ _02612_ _02613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05193_ cpu.regs\[12\]\[0\] cpu.regs\[13\]\[0\] cpu.regs\[14\]\[0\] cpu.regs\[15\]\[0\]
+ _00858_ _00859_ _00865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XPHY_EDGE_ROW_47_Left_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06587__A2 _00948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08952_ _04009_ _04135_ _04157_ _04158_ _04159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07903_ _03312_ _03313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08883_ _04070_ _04091_ _04092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07834_ cpu.uart.counter\[1\] _03254_ _03256_ _03257_ _03258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_47_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04977_ cpu.instr_cycle\[3\] cpu.instr_cycle\[1\] _00677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07765_ _03200_ _03201_ _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_79_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_95_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06716_ _00579_ _00633_ _02367_ _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09504_ _03815_ _04665_ _04668_ _00514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07696_ cpu.uart.div_counter\[6\] _03145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09435_ cpu.ROM_spi_dat_out\[2\] _04562_ _04612_ _04613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06647_ cpu.startup_cycle\[4\] _02300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_56_Left_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05314__A3 _00981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09366_ _01000_ _02334_ _04555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06578_ _01935_ _02234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09297_ cpu.last_addr\[13\] _04491_ _04492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05529_ _01017_ _01195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08317_ _03622_ _03628_ _03629_ _00366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_35_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08248_ _02478_ _03551_ _03580_ _03582_ _03583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10210_ _00468_ clknet_leaf_53_wb_clk_i cpu.IE vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_65_Left_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08179_ cpu.toggle_ctr\[0\] _03528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10141_ _00400_ clknet_leaf_4_wb_clk_i cpu.timer_capture\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05250__A2 _00918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10072_ _00331_ clknet_leaf_0_wb_clk_i cpu.toggle_ctr\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09742__B _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_74_Left_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_qcpu_113 io_oeb[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xwrapped_qcpu_102 io_oeb[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_108_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06266__A1 _01906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09204__A1 _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04900_ cpu.br_rel_dest\[7\] _00602_ _00603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05880_ _00904_ _01343_ _01541_ _01341_ _01434_ _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_108_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07550_ _03013_ _03024_ _03027_ _00201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06501_ _02133_ _02135_ _02158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09220_ _04386_ _04387_ _04391_ _04418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07481_ _02952_ _02965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08494__A2 _02513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06432_ _00814_ _00871_ _02089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09151_ _00696_ _04351_ _04136_ _04352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06363_ _00783_ _02019_ _02020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_17_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08102_ cpu.orig_PC\[10\] _03464_ _03457_ _03465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09082_ _04179_ _04275_ _04282_ _04284_ _04186_ _04285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05314_ _00608_ _00964_ _00981_ _00982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_08033_ cpu.orig_IO_addr_buff\[4\] _03408_ _03411_ _03414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06294_ _01950_ _01951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05245_ _00914_ _00915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_31_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05480__A2 _01145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05176_ _00007_ _00848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_40_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09984_ _00243_ clknet_leaf_27_wb_clk_i cpu.uart.div_counter\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05646__I _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05232__A2 _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08935_ _03441_ _01531_ _04142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input21_I io_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08866_ _00637_ _01115_ _04049_ _04075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_98_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08797_ _03839_ _04009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07817_ cpu.uart.div_counter\[15\] _03210_ _03237_ _03244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07748_ _03188_ _00238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_67_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07679_ _03127_ cpu.uart.div_counter\[9\] cpu.uart.div_counter\[2\] _02638_ _03128_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_67_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09418_ cpu.ROM_spi_dat_out\[0\] _04598_ _03904_ _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_109_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07693__B1 _01183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09434__A1 _02359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09349_ _03057_ _04539_ _04540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_75_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10124_ _00383_ clknet_leaf_6_wb_clk_i cpu.timer\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06420__A1 _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10055_ _00314_ clknet_leaf_72_wb_clk_i cpu.orig_PC\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__04982__A1 _00680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_82_Left_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_89_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05082__S1 _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05782__I0 _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_46_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_91_Left_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05030_ _00713_ _00720_ _00725_ _00726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__05214__A2 _00884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06981_ _00798_ _02567_ _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_47_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_47_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05932_ cpu.timer_capture\[3\] _01221_ _01232_ _01595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08720_ _03942_ cpu.regs\[3\]\[2\] _03950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08651_ _03838_ _03894_ _03895_ _03896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05863_ _01309_ _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_07602_ cpu.spi.div_counter\[6\] _03065_ _03062_ _03069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08582_ _03833_ _03826_ _03834_ _00426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_88_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05794_ _00726_ _01449_ _01459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07533_ _03010_ _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08726__B _03954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07464_ cpu.timer_top\[14\] _02948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_91_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09203_ _04268_ _04383_ _04402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06415_ cpu.multiplier.a\[7\] _02069_ _02071_ _02072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__06246__B _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09134_ _02211_ _01157_ _04335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07395_ _02127_ _02874_ _02886_ _02888_ _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_44_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08017__I _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06346_ _00871_ _02002_ _02003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09065_ _04268_ _04242_ _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06277_ _01933_ _01934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08016_ _03400_ _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05453__A2 _01118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05228_ _00892_ _00899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_69_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05159_ _00830_ _00831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_110_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09967_ _00226_ clknet_leaf_36_wb_clk_i cpu.uart.dout\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08918_ _04099_ _04102_ _04125_ _00680_ _04126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_99_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09898_ _00157_ clknet_leaf_110_wb_clk_i cpu.regs\[6\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08849_ _02418_ _00667_ _00985_ _01297_ _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_95_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06603__C _02258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08597__I _03848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10107_ _00366_ clknet_leaf_7_wb_clk_i cpu.timer_div_counter\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10038_ _00297_ clknet_leaf_14_wb_clk_i cpu.orig_IO_addr_buff\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06200_ _00826_ _01760_ _01859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_116_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06880__A1 cpu.timer_capture\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07180_ _02741_ _00117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06131_ _00979_ _01515_ _01791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_41_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06062_ cpu.toggle_top\[13\] _01723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_69_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05013_ _00702_ _00706_ _00709_ _00003_ _00710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_41_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09821_ _00080_ clknet_leaf_34_wb_clk_i cpu.uart.receive_counter\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05038__I2 cpu.regs\[6\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09752_ _00015_ clknet_leaf_106_wb_clk_i cpu.regs\[15\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08703_ _03812_ _03937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08137__A1 cpu.toggle_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06964_ _01926_ _02579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05915_ _01476_ _01576_ _01577_ _01578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08300__I _02379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06895_ _01031_ _02433_ _02519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09683_ _01659_ _00949_ _01744_ _04809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_96_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08634_ _03862_ _03880_ _03881_ _03882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05846_ cpu.toggle_top\[2\] _01171_ _01173_ _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08565_ _02446_ _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05777_ _00879_ _01150_ _01324_ _01442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07516_ _00631_ _02999_ _00195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_91_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08496_ _03757_ _03774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07447_ cpu.timer_div\[4\] cpu.timer_div_counter\[4\] _02931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_40_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08970__I _04101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07378_ _02209_ _02872_ _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09117_ _04268_ _04303_ _04319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06329_ _01977_ _01978_ _01982_ _01983_ _01986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_45_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09048_ _02214_ _01140_ _04251_ _04252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__05426__A2 _01018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06623__A1 _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output52_I net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05037__S1 _00731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06614__A1 _01759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07406__A3 _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04913__I _00615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05268__I2 cpu.regs\[6\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_10_Left_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__04928__A1 _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08119__A1 cpu.toggle_top\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_2_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06680_ _02332_ _02333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05700_ cpu.PORTB_DDR\[1\] _01364_ _01365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05631_ _01296_ _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_106_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08350_ _03650_ _03651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05562_ _01227_ _01228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07301_ _02788_ _02811_ _02817_ _00162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05493_ _00910_ _00876_ _01158_ _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_46_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08281_ cpu.pwm_top\[0\] _03605_ _03484_ _03606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05656__A2 _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07232_ _02753_ cpu.regs\[8\]\[4\] _02764_ _02772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_54_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07163_ _02730_ _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06114_ _00615_ _01773_ _01774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07094_ _02685_ _02686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_62_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_62_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_100_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06045_ cpu.uart.divisor\[13\] _01382_ _01705_ _00012_ _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_2_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09804_ _00067_ clknet_leaf_116_wb_clk_i cpu.toggle_top\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07996_ _03383_ _03379_ _03385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_70_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06947_ _02559_ _02560_ _02561_ _02562_ _02563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_09735_ _02579_ _04846_ _04849_ _04850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09666_ _04039_ _04790_ _04791_ _04792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08617_ _01430_ _03867_ _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06878_ _02503_ _02496_ _02497_ _02504_ _02505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09597_ _00575_ _04729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_96_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05829_ _01491_ _01492_ _01177_ _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08548_ _00674_ _00612_ _01041_ _03808_ _03809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_77_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_53_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08479_ _03739_ _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_37_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09464__C _03398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07021__A1 _01842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05258__S1 _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05335__A1 _00691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_46_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09077__A2 _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05638__A2 _01018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05110__I1 _00798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07850_ _03268_ _03266_ _03270_ _03271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06801_ _02439_ _02440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_04993_ _00691_ _00692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07781_ cpu.uart.div_counter\[8\] _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_85_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput3 io_in[11] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09520_ _03804_ _04672_ _04678_ _00520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_108_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06732_ _01160_ _02377_ _02379_ _02383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08512__A1 cpu.spi.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09451_ _04593_ _04624_ _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06663_ cpu.mem_cycle\[0\] _02316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_94_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09382_ _04558_ _04567_ _00493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05614_ _01033_ _01101_ _01007_ _01280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_47_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05877__A2 _00904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06594_ _02239_ _02249_ _02250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08402_ _03653_ _03695_ _03696_ _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05545_ _01209_ _01010_ _01210_ _01211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_74_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08333_ cpu.timer_top\[10\] _03637_ _03640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08264_ _03588_ _03592_ _03593_ _00349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_116_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05476_ _01139_ _00599_ _01141_ _01142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_61_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08195_ _03522_ _03532_ _03543_ _03529_ _03544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07215_ _01658_ _01676_ _02762_ _00131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08579__A1 _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08025__I _03407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07146_ _02712_ _02720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07077_ _02456_ _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06028_ _00965_ _01688_ _00849_ _01689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07979_ _03370_ _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09718_ _02548_ _02549_ _04834_ _04835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_69_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08503__A1 _02518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07306__A2 _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09649_ _02331_ _04521_ _04524_ _04776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_97_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05868__A2 _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06943__I _02558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07242__A1 _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10286_ _00544_ clknet_leaf_99_wb_clk_i cpu.PORTA_DDR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_2_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05308__A1 _00843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05330_ _00995_ _00586_ _00996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05261_ _00897_ net122 _00930_ _00931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_114_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_72_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05192_ _00861_ _00863_ _00864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07000_ _02610_ _02612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05095__I0 cpu.regs\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_102_Left_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08951_ _00659_ _04158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07902_ cpu.uart.receiving _02666_ _03311_ _03312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_08882_ _01336_ _00984_ _01454_ _04091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_07833_ _02483_ _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_81_Right_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07764_ _03133_ _03197_ _03201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_79_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04976_ _00614_ _00662_ _00670_ _00675_ _00676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_78_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06715_ _00647_ net18 _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09503_ net59 _04666_ _04667_ _04668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07695_ cpu.uart.div_counter\[12\] _03144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09434_ _02359_ _04611_ _04612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06646_ cpu.startup_cycle\[5\] _02299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_94_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_111_Left_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_63_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09365_ _04545_ _04553_ _02353_ _02359_ _04554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_06577_ _01934_ _02232_ _02233_ _00022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09296_ cpu.last_addr\[12\] cpu.last_addr\[11\] _04490_ _04491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_05528_ _01190_ _01193_ _01194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08316_ cpu.timer_div_counter\[3\] _03625_ cpu.timer_div_counter\[4\] _03629_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_90_Right_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05459_ _00606_ _01003_ _01117_ _01125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_62_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08247_ _03495_ _03581_ _03582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09213__A2 _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08178_ _03526_ _01417_ _03527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_30_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07129_ _01753_ _02700_ _02707_ _00100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10140_ _00399_ clknet_leaf_4_wb_clk_i cpu.timer_capture\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10071_ _00330_ clknet_leaf_0_wb_clk_i cpu.toggle_ctr\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_qcpu_114 io_oeb[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xwrapped_qcpu_103 io_oeb[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_58_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05289__I _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08963__A1 _00728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_119_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_119_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10269_ _00527_ clknet_leaf_44_wb_clk_i net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_108_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07480_ _02957_ _02961_ _02963_ _02964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06500_ _02146_ _02155_ _02156_ _02157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_60_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06431_ _02083_ _02087_ _02088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_32_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09150_ _04103_ _04351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_84_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05701__B _01018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06362_ net127 _02018_ _02002_ _00883_ _02019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_16_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08101_ _03400_ _03464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09081_ _04249_ _04283_ _04284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05313_ _00980_ _00981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06293_ cpu.multiplier.a\[0\] _01950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08032_ _03401_ _03413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05244_ _00902_ _00896_ _00887_ _00914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07206__A1 _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05175_ cpu.regs\[12\]\[1\] cpu.regs\[13\]\[1\] cpu.regs\[14\]\[1\] cpu.regs\[15\]\[1\]
+ _00836_ _00839_ _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_40_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06009__A2 _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09983_ _00242_ clknet_leaf_27_wb_clk_i cpu.uart.div_counter\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05768__A1 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08934_ _04139_ _04111_ _04140_ _04141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_4_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08865_ _04070_ _04073_ _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07816_ _03213_ _03243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08796_ _00658_ _04008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08182__A2 cpu.toggle_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input14_I io_in[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07747_ _02677_ _03187_ _03188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_79_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04959_ _00651_ _00638_ _00658_ _00659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_67_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05940__A1 cpu.toggle_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07678_ _02628_ _03127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08973__I _04138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09417_ _04593_ _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06629_ _01867_ _02283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09348_ _04478_ _04479_ _04521_ _04538_ _04539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_118_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09279_ _00784_ _04452_ _04474_ _04475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output82_I net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10123_ _00382_ clknet_leaf_6_wb_clk_i cpu.timer\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10054_ _00313_ clknet_leaf_72_wb_clk_i cpu.orig_PC\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06184__A1 _00650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09044__I _00661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06184__B2 _01842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05782__I1 _00851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_7_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09673__A2 _04008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04916__I net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05298__I0 cpu.regs\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08551__C _00626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06980_ _01815_ _02554_ _02593_ _02594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input6_I io_in[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05931_ cpu.timer_div\[3\] _01400_ _01402_ _01594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08650_ _02423_ _03851_ _03895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06175__A1 cpu.timer_capture\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05862_ _01525_ _01431_ _01432_ _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07601_ _03067_ _03068_ _00211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_89_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08581_ cpu.uart.divisor\[15\] _03827_ _03830_ _03834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05922__A1 cpu.uart.divisor\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09113__A1 _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05793_ _01437_ _01449_ _01458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_87_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_87_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07532_ _02427_ _03007_ _03012_ _00198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_16_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_16_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_44_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06022__S1 _00969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07463_ _02946_ cpu.timer\[15\] _02947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09202_ _04300_ _04383_ _04400_ _04317_ _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06414_ cpu.multiplier.a\[7\] _02070_ _02071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07427__A1 cpu.spi.dout\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09133_ _04305_ _04332_ _04333_ _04334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__07202__I _01814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07394_ _02573_ _02887_ _02888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_72_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06345_ _02001_ _02002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09064_ _04165_ _04268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06276_ _01927_ _01931_ _01932_ _01933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08015_ _03399_ _03400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05227_ _00835_ _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_69_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05158_ _00006_ _00830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_40_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09966_ _00225_ clknet_leaf_38_wb_clk_i cpu.uart.dout\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06402__A2 _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05089_ cpu.multiplier.a\[5\] _00781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08917_ _00666_ _04105_ _04124_ _00670_ _04125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09897_ _00156_ clknet_leaf_91_wb_clk_i cpu.regs\[6\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08848_ _01278_ _00919_ _04057_ _04058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__06166__A1 _01824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08779_ _03966_ _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05913__A1 cpu.PORTB_DDR\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08918__B2 _00680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09591__A1 _02540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10106_ _00365_ clknet_leaf_22_wb_clk_i cpu.timer_div_counter\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10037_ _00296_ clknet_leaf_14_wb_clk_i cpu.orig_IO_addr_buff\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09502__I _03829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08118__I _03473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07409__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08082__A1 _02556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06130_ _01787_ _01788_ _01789_ _01790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06061_ cpu.toggle_top\[5\] _01254_ _01260_ _01721_ _01722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_10_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05012_ _00707_ _00708_ _00709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09820_ _00079_ clknet_leaf_33_wb_clk_i cpu.uart.receive_counter\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09751_ _00014_ clknet_leaf_101_wb_clk_i cpu.regs\[15\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06935__A3 _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06963_ net12 _02559_ _02578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08702_ cpu.ROM_addr_buff\[6\] _03936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05914_ net62 _01198_ _01577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06894_ _02426_ _02518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09682_ _01566_ _04806_ _04807_ _04808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_96_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08633_ _02416_ _03867_ _03881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05845_ cpu.pwm_top\[2\] _01252_ _01254_ _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08564_ _03820_ _03817_ _03822_ _00420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_89_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05776_ _00829_ _01149_ _01441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07515_ _00628_ _02998_ cpu.needs_timer_interrupt _02999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08495_ cpu.timer\[15\] _03761_ _03772_ _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07446_ _02927_ _02928_ _02930_ _00194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_91_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08028__I _02455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07377_ _02211_ _02857_ _02872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09116_ _04300_ _04303_ _04316_ _04317_ _04318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06328_ _01979_ _01984_ _01960_ _01985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_103_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09047_ _04219_ _04250_ _04251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05426__A3 _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06259_ _01913_ _01915_ _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_75_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09573__A1 cpu.PORTA_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09949_ _00208_ clknet_leaf_37_wb_clk_i cpu.spi.div_counter\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_48_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_36_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08366__C _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09564__A1 _02536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06378__A1 _01950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_75_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05630_ _01295_ _01296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_116_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09619__A2 _04748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05561_ _01226_ _01227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07300_ cpu.regs\[5\]\[3\] _02815_ _02817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05492_ _01156_ _01157_ _01158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08280_ _03602_ _03605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07231_ _02722_ _02765_ _02771_ _00138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07162_ _01165_ _02729_ _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06113_ cpu.uart.divisor\[14\] _01380_ _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07093_ _01113_ _02684_ _02685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06044_ _01695_ _01375_ _01696_ _01704_ _01484_ _01705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_2_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09555__A1 _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05935__I _01410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09803_ _00066_ clknet_leaf_84_wb_clk_i cpu.multiplier.a\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07995_ _03383_ _03379_ _03384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_70_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_31_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_31_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06946_ net1 _02236_ _02203_ _02562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09734_ _02236_ _04848_ _02590_ _02256_ _04849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07869__A1 _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09665_ _00988_ _01990_ _04037_ _04791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06877_ cpu.timer\[5\] _02499_ _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05828_ cpu.spi.divisor\[2\] _01134_ _01492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08616_ _03850_ _03867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09596_ _02297_ _02298_ _04728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08547_ _00650_ _01115_ _00647_ _00566_ _03808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_77_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05759_ _01271_ _01275_ _00904_ _01424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_25_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08478_ _03740_ _03756_ _03759_ _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08294__A1 _02454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07429_ _02917_ _02918_ _02915_ _00189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_81_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06780__A1 _02421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06532__A1 _02186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05638__A3 _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06599__A1 _02254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05110__I2 cpu.regs\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07780_ _03213_ _03214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04992_ net25 _00691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_06800_ _02390_ _02439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput4 io_in[12] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_108_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06731_ _02381_ _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09450_ cpu.ROM_spi_dat_out\[6\] _02360_ _04612_ _04624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06662_ _02300_ _02311_ _02314_ _02315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_78_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08401_ cpu.timer_capture\[6\] _03660_ _03675_ _03696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09381_ _04566_ _04561_ _04567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05613_ _01269_ _01271_ _01277_ _01278_ _01279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06593_ _02246_ _02248_ _02249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05544_ _00587_ _01207_ _01210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_47_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08332_ _02525_ _03636_ _03639_ _02542_ _00371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08276__A1 _03585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08263_ cpu.pwm_counter\[3\] _03591_ _03593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05475_ _01140_ _00638_ _00613_ _01141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_61_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07214_ _02760_ _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08194_ _03526_ _01417_ _03543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07145_ _01551_ _02719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07076_ cpu.uart.receive_counter\[2\] _02669_ _02674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09528__A1 _03815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06027_ cpu.regs\[8\]\[6\] cpu.regs\[9\]\[6\] cpu.regs\[10\]\[6\] cpu.regs\[11\]\[6\]
+ _00968_ _00969_ _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_2_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05014__A1 _00003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07978_ _02363_ _03370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09717_ _02393_ _01906_ _02397_ _04834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_58_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06762__A1 _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06929_ _01153_ _02544_ _02545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09700__A1 _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09648_ _04754_ _04772_ _04775_ _03398_ _00551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_97_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09579_ cpu.PORTA_DDR\[3\] _04712_ _04713_ _04717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_38_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08267__A1 _03585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07242__A2 _02777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09519__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10285_ _00543_ clknet_leaf_99_wb_clk_i cpu.PORTA_DDR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_103_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05260_ _00888_ _00929_ _00930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_52_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05191_ _00833_ _00862_ _00845_ _00863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05095__I1 _00783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08950_ cpu.orig_PC\[2\] _03840_ _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05485__I _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07901_ cpu.uart.receive_counter\[0\] cpu.uart.receive_counter\[1\] cpu.uart.receive_counter\[3\]
+ cpu.uart.receive_counter\[2\] _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_08881_ _00641_ _02430_ _04089_ _04090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08733__A2 cpu.regs\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07832_ _03255_ cpu.uart.counter\[1\] _03250_ _03256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09502_ _03829_ _04667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07763_ _03124_ _03149_ _03156_ _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_04975_ _00671_ _00673_ _00674_ _00675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06714_ _02294_ _02334_ _02366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07694_ _03128_ _03132_ _03135_ _03142_ _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_69_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09433_ _04610_ _04596_ _04611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06645_ _01038_ _02298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_94_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09364_ _04546_ _04547_ _02301_ _04552_ _04553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_93_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08315_ cpu.timer_div_counter\[3\] cpu.timer_div_counter\[4\] _03625_ _03628_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06576_ _00769_ _01934_ _02233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09295_ _03999_ _04489_ _04490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05527_ net79 cpu.PORTA_DDR\[0\] _01192_ _01193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_62_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05458_ _01121_ _01122_ _01123_ _01124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_62_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08246_ cpu.toggle_ctr\[13\] _03578_ _03581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06275__A3 _01118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08177_ cpu.toggle_ctr\[1\] _03526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05389_ _01054_ _01055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_70_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07128_ cpu.regs\[13\]\[5\] _02703_ _02707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07059_ cpu.uart.receive_div_counter\[6\] _02659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10070_ _00329_ clknet_leaf_117_wb_clk_i cpu.toggle_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XPHY_EDGE_ROW_102_Right_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08488__A1 cpu.timer_capture\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_qcpu_104 io_oeb[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_69_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07215__A2 _01676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05777__A2 _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10268_ _00526_ clknet_leaf_42_wb_clk_i net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10199_ _00457_ clknet_leaf_66_wb_clk_i cpu.last_addr\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06430_ _02086_ _02085_ _02087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_75_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06361_ _02017_ _02018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08100_ _02208_ _03463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09080_ _04280_ _04281_ _04279_ _04283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05312_ _00979_ _00980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06292_ _01945_ _01948_ _01949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_71_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05465__A1 _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05243_ _00912_ _00913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08031_ _01069_ _03402_ _03412_ _00297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_25_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05174_ _00843_ _00844_ _00845_ _00846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_09982_ _00241_ clknet_leaf_26_wb_clk_i cpu.uart.div_counter\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08933_ cpu.PC\[1\] _01149_ _04140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08706__A2 cpu.regs\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08167__B1 cpu.toggle_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06717__A1 _02366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08864_ _04072_ _04073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04987__C _00686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08795_ _02429_ _04007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07815_ _03240_ _03241_ _03242_ _00251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07390__A1 _02203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07746_ _03136_ _03185_ _03186_ _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04958_ _00657_ _00658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09131__A2 _00652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09416_ _04587_ _04596_ _04583_ _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07677_ cpu.uart.div_counter\[4\] _01628_ _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_04889_ cpu.IO_addr_buff\[4\] _00592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07693__A2 _02441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09150__I _04103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06628_ _01934_ _02281_ _02282_ _00024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09347_ _04535_ _04537_ _04538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06559_ _02215_ _02216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09278_ _04452_ _04459_ _04474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08229_ cpu.toggle_ctr\[7\] _03568_ cpu.toggle_ctr\[8\] _03570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_78_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output75_I net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06956__A1 _02556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10122_ _00381_ clknet_leaf_6_wb_clk_i cpu.timer\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10053_ _00312_ clknet_leaf_64_wb_clk_i cpu.orig_PC\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_89_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06184__A2 _01057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07381__A1 _02573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08633__A1 _02416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05298__I1 cpu.multiplier.a\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05930_ cpu.spi.dout\[3\] _01181_ _01392_ _01592_ _01396_ _01593_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_28_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05861_ _00988_ _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07600_ _03065_ _03062_ _00645_ _03068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08580_ _02466_ _03833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_88_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07531_ cpu.spi.data_out_buff\[0\] _03008_ _03011_ _02404_ _03012_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_66_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05792_ _01456_ _01457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_88_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07462_ cpu.timer_top\[15\] _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_45_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09201_ _04385_ _04399_ _04400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05230__S0 _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07393_ _02885_ net121 _02152_ _02887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_06413_ _00781_ cpu.multiplier.a\[6\] _02070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xclkbuf_leaf_56_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_56_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_72_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09132_ _02212_ _01110_ _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06344_ cpu.multiplier.a\[3\] _00767_ _02001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09063_ _00680_ _04267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06275_ _01619_ _01043_ _01118_ _01932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_08014_ _00617_ _00642_ _00622_ _00677_ _03399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_05226_ _00007_ _00897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05157_ cpu.base_address\[1\] _00829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08388__B1 _03681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07060__B1 cpu.uart.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09965_ _00224_ clknet_leaf_36_wb_clk_i cpu.uart.dout\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05088_ _00780_ net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_08916_ _04106_ _00660_ _04121_ _04123_ _04124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_09896_ _00155_ clknet_leaf_110_wb_clk_i cpu.regs\[6\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09145__I _00661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08847_ _00932_ _01694_ _00981_ _01693_ _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__07363__A1 _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08778_ _03984_ _03994_ _03995_ _00461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_clkbuf_leaf_26_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09104__A2 _02423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07729_ _01899_ _03172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_95_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05429__A1 _00663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_65_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10105_ _00364_ clknet_leaf_21_wb_clk_i cpu.timer_div_counter\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10036_ _00295_ clknet_leaf_50_wb_clk_i cpu.orig_IO_addr_buff\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04927__I _00622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05380__A3 _01001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05668__A1 _00711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06060_ _01718_ _01719_ _01720_ _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05011_ cpu.regs\[12\]\[0\] cpu.regs\[13\]\[0\] cpu.regs\[14\]\[0\] cpu.regs\[15\]\[0\]
+ _00703_ _00704_ _00708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__09031__A1 _02389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_103_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_103_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06962_ _02027_ _02576_ _02008_ _02577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09750_ _00013_ clknet_leaf_102_wb_clk_i cpu.regs\[15\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08701_ _03453_ _03933_ _03934_ _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05913_ cpu.PORTB_DDR\[3\] _01202_ _01239_ _01363_ _01574_ _01575_ _01576_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
X_09681_ _00765_ _00958_ _04807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08632_ cpu.orig_IO_addr_buff\[4\] _03864_ _03865_ _00950_ _03880_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06893_ _02517_ _00054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07345__A1 _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07896__A2 net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05844_ _01502_ _01504_ _01507_ _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08563_ _02628_ _03818_ _03821_ _03822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05775_ _01439_ _01323_ _01440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_76_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08494_ _03743_ _02513_ _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07514_ _02944_ _02997_ _02998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_07445_ _02929_ _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07376_ net12 _02855_ _02871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09115_ _04161_ _04317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06327_ _01982_ _01983_ _01984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06258_ _01914_ _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09046_ _04217_ _04218_ _04250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05131__I0 cpu.regs\[8\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05209_ _00879_ _00880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06189_ _01335_ _01271_ _01847_ _01692_ _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09948_ _00207_ clknet_leaf_47_wb_clk_i cpu.spi.div_counter\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09879_ _00138_ clknet_leaf_105_wb_clk_i cpu.regs\[8\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_86_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05898__A1 _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output38_I net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08836__A1 _01151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06075__A1 _00796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07111__I1 _02283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05822__A1 cpu.uart.divisor\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_1_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_1_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09494__B net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07575__A1 _03043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06378__A2 _00978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10019_ _00278_ clknet_leaf_32_wb_clk_i cpu.uart.receive_div_counter\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07742__B _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09513__I _03607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05560_ _01025_ _01225_ _01226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_106_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08827__A1 _01107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08129__I _03473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05491_ cpu.base_address\[0\] _01157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_58_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07230_ cpu.regs\[8\]\[3\] _02769_ _02771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07161_ _01109_ _01111_ _01106_ _02729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_14_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06112_ _01771_ _01374_ _01381_ _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07092_ _01929_ _02684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_06043_ net11 _01121_ _01701_ _01703_ _01704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_100_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07566__A1 cpu.spi.data_out_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09802_ _00065_ clknet_leaf_84_wb_clk_i cpu.multiplier.a\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09307__A2 cpu.ROM_addr_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07994_ cpu.uart.receive_div_counter\[13\] _03383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06945_ _01989_ _02005_ _02561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09733_ _01942_ _04847_ _04839_ _04848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06876_ _00981_ _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09664_ _04044_ _04046_ _04041_ _04790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09595_ _04600_ _02304_ _02336_ _04727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09423__I _03829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05827_ _01011_ _00999_ _01489_ _01490_ _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_08615_ cpu.orig_IO_addr_buff\[1\] _03864_ _03865_ _01278_ _03866_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_96_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08546_ _00648_ net18 _03807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08039__I _03407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05758_ _01335_ _01265_ _01421_ _01422_ _01423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_25_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_53_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05689_ cpu.regs\[15\]\[0\] _01354_ _01355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08477_ cpu.timer_capture\[11\] _03746_ _03758_ _03759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08294__A2 _03613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07428_ cpu.spi.data_in_buff\[2\] _02907_ _02918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_81_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06782__I _01110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07359_ _02851_ _02855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_103_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09029_ _00768_ _04232_ _04233_ _04234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08658__B _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06780__A2 _02413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08809__A1 cpu.IE vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09482__A1 cpu.pwm_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06296__A1 _01952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_116_Right_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07028__I cpu.uart.divisor\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04991_ _00689_ _00629_ _00690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput5 io_in[13] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_108_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06730_ net12 _02374_ _02381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06867__I _01694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06661_ _02312_ _02313_ _02296_ _02314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_05612_ _00884_ _01278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08400_ _02509_ _03692_ _03657_ _03694_ _03695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09380_ _02312_ _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06592_ _02009_ _02247_ _02248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_05543_ cpu.uart.divisor\[8\] _01209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08331_ cpu.timer_top\[9\] _03637_ _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05474_ _00601_ _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_50_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08262_ cpu.pwm_counter\[3\] _03591_ _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07213_ _01616_ _02761_ _00130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06039__A1 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08193_ _03519_ _03518_ _03532_ cpu.toggle_ctr\[2\] _03542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_07144_ _02717_ _02714_ _02718_ _00104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_30_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07075_ cpu.uart.receive_counter\[0\] cpu.uart.receive_counter\[1\] _02667_ _02673_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_112_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06026_ _01686_ _00843_ _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07977_ _03327_ _03369_ _00286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_58_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06762__A2 _02400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09716_ _01351_ _02555_ _04832_ _04833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07382__B _02876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06928_ _01164_ _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09647_ _04600_ _04774_ _04772_ _02347_ _04775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_83_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06859_ _02488_ _00049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_2_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09578_ _02527_ _04711_ _04716_ _00540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08529_ _01496_ _03790_ _03795_ _03648_ _00412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_38_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06017__I _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07778__A1 _03088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10284_ _00542_ clknet_leaf_99_wb_clk_i cpu.PORTA_DDR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09063__I _00680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05190_ cpu.regs\[0\]\[0\] cpu.multiplier.a\[0\] cpu.regs\[2\]\[0\] cpu.regs\[3\]\[0\]
+ _00858_ _00859_ _00862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_24_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05766__I _01304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05095__I2 _00784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07900_ _02679_ _02678_ _03309_ _03310_ _00268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_08880_ _00658_ _04077_ _04088_ _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07831_ cpu.uart.counter\[0\] _03255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05627__S0 _01285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06744__A2 _02388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_16_Left_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08298__B _03615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09501_ _04664_ _04666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07762_ _03198_ _03199_ _00241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_04974_ _00663_ _00674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_2_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06713_ _02350_ _02362_ _02365_ _00026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07693_ _03136_ _02441_ _01183_ _03137_ _03141_ _03142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_79_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05434__C _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09432_ _04566_ _04585_ _04571_ _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06644_ _02296_ _02297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09363_ _02298_ _04551_ _04552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06575_ _01678_ _01936_ _02231_ _02232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05526_ _01046_ _01191_ _01192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_63_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08314_ _03623_ _03627_ _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09294_ cpu.last_addr\[9\] cpu.last_addr\[8\] _04488_ _04489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__05307__I0 cpu.regs\[12\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_25_Left_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05457_ _00995_ _01071_ _01120_ _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_62_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08245_ cpu.toggle_ctr\[14\] cpu.toggle_ctr\[13\] _03578_ _03580_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_117_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05388_ _00588_ _01047_ _01050_ _01054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08176_ _03513_ _03516_ _03520_ _03524_ _03525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_113_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07127_ _02706_ _00099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06432__A1 _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07058_ cpu.uart.receive_div_counter\[12\] _02658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08052__I cpu.IE vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06009_ _01659_ _01670_ _01671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_7_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07232__I0 _02753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_34_Left_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09685__A1 _00811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_qcpu_105 io_oeb[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_85_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_43_Left_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_52_Left_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10267_ _00525_ clknet_leaf_46_wb_clk_i net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10198_ _00456_ clknet_leaf_66_wb_clk_i cpu.last_addr\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07923__B2 net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06210__I _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_61_Left_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06360_ _00781_ _02014_ _02016_ _02017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_33_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06291_ _01447_ _01446_ _00902_ _00896_ _00888_ _01947_ _01948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_05311_ _00978_ _00979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput30 sram_out[4] net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08581__B _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05242_ _00877_ _00912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08030_ cpu.orig_IO_addr_buff\[3\] _03408_ _03411_ _03412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_5_0_wb_clk_i clknet_0_wb_clk_i clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_05173_ _00007_ _00845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09981_ _00240_ clknet_leaf_30_wb_clk_i cpu.uart.div_counter\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06414__A1 cpu.multiplier.a\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08932_ cpu.PC\[1\] cpu.br_rel_dest\[1\] _04139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06965__A2 _02577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08863_ _04071_ _04072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08794_ _00686_ _04005_ _04006_ _00466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07814_ _02929_ _03242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07745_ _03136_ _03137_ _03181_ _03186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_79_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04957_ _00654_ _00656_ _00613_ _00657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_clkbuf_leaf_16_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09667__A1 _02070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07390__A2 _02883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06025__S0 _00891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09415_ _04589_ _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07676_ cpu.uart.divisor\[11\] cpu.uart.div_counter\[11\] _03125_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_04888_ cpu.IO_addr_buff\[3\] _00591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_48_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06627_ cpu.regs\[2\]\[6\] _01933_ _02282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09346_ _01910_ _04536_ _04537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06558_ cpu.PC\[4\] _02215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_90_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09277_ _04137_ _04459_ _04472_ _04162_ _04473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05509_ _01064_ _01065_ _00989_ _01175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_62_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06489_ _02106_ _02111_ _02145_ _02146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_118_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08228_ _03563_ _03569_ _00337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08159_ _03494_ _01842_ _03506_ _03507_ _03508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_31_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_55_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10121_ _00380_ clknet_leaf_8_wb_clk_i cpu.timer\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output68_I net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10052_ _00311_ clknet_leaf_73_wb_clk_i cpu.orig_PC\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08510__I _03776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06184__A3 _01273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08666__B _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08330__A1 _02518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06186__B _01273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06892__A1 cpu.timer_capture\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09497__B _03043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_94_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06247__I1 net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06947__A2 _02560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05860_ _01304_ _01523_ _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_89_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05791_ _00881_ _01330_ _01329_ _01456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__08576__B _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07530_ _03010_ _03011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_66_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08872__A2 _04080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07461_ _00687_ _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_17_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09200_ _04248_ _04395_ _04398_ _04399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_8_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05230__S1 _00899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07392_ _02885_ _02152_ _02886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06412_ _00782_ _00798_ _02069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09131_ cpu.PC\[7\] _00652_ _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06343_ _01980_ _01998_ _01999_ _02000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09062_ _04176_ _04242_ _04265_ _04202_ _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_71_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06635__A1 _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_96_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_96_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06274_ _01930_ _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08013_ _00617_ _00623_ _03397_ _03398_ _00293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xclkbuf_leaf_25_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_25_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_71_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05225_ _00894_ _00895_ _00832_ _00896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05156_ _00828_ net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09964_ _00223_ clknet_leaf_36_wb_clk_i cpu.uart.dout\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05087_ _00766_ _00774_ _00779_ _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_85_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08915_ cpu.orig_PC\[1\] _04075_ _04122_ _04106_ _04123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09895_ _00154_ clknet_leaf_88_wb_clk_i cpu.regs\[6\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08846_ cpu.orig_flags\[1\] _03841_ _04053_ _04055_ _04056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__05374__A1 _00618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08560__A1 _03815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08777_ cpu.ROM_addr_buff\[8\] _03988_ _03995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05989_ _01648_ _01649_ _01650_ _01651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07728_ _02440_ _03171_ _00234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07659_ cpu.uart.receive_buff\[6\] _03102_ _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06874__A1 cpu.timer_capture\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09329_ _04523_ _00484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_11_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08615__A2 _03864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06626__A1 _01815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10104_ _00363_ clknet_leaf_20_wb_clk_i cpu.timer_div_counter\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10035_ _00294_ clknet_leaf_50_wb_clk_i cpu.orig_IO_addr_buff\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08303__A1 _03618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05668__A2 _01333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06617__A1 _02271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05010_ _00002_ _00707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08790__A1 cpu.ROM_addr_buff\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06961_ _02010_ _02013_ _02576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08700_ _03926_ cpu.regs\[2\]\[6\] _03934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05912_ net82 _00596_ _01358_ _01127_ _01575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_72_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09680_ _00742_ _00918_ _04805_ _04806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08631_ _03860_ _03879_ _00430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06892_ cpu.timer_capture\[7\] _02494_ _02516_ _02506_ _02517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_55_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05843_ _01506_ _01507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_89_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08562_ _03757_ _03821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05774_ _00711_ _01320_ _01439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08493_ _03760_ _03770_ _03771_ _00400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07513_ _02996_ _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_07444_ _02363_ _02929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08845__A2 _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07375_ _02854_ _02868_ _02870_ _00183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09114_ _04309_ _04313_ _04315_ _04316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06326_ _01951_ _01980_ _00954_ _01983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_44_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06257_ cpu.mem_cycle\[0\] _01914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09045_ _04108_ _04249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05208_ cpu.base_address\[1\] _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06188_ _01618_ _01270_ _01847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05139_ cpu.PORTB_DDR\[3\] net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XPHY_EDGE_ROW_8_Left_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09947_ _00206_ clknet_leaf_45_wb_clk_i cpu.spi.div_counter\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08060__I _03432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09878_ _00137_ clknet_leaf_105_wb_clk_i cpu.regs\[8\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08829_ _01108_ _01942_ _04039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_86_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09105__B _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06847__A1 cpu.timer_capture\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08836__A2 _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09013__A2 _01618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05808__B cpu.PORTA_DDR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10018_ _00277_ clknet_leaf_31_wb_clk_i cpu.uart.receive_div_counter\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_47_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08827__A2 _01942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05490_ _00829_ _01156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07160_ _01869_ _02715_ _02728_ _00110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06111_ cpu.uart.divisor\[6\] _01771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07091_ _02387_ _02683_ _02424_ _00086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_54_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06066__A2 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06042_ _01702_ _01189_ _01370_ _01703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07015__A1 _02454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09801_ _00064_ clknet_leaf_84_wb_clk_i cpu.multiplier.a\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07993_ _03371_ _03382_ _00289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09732_ _01960_ _01966_ _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08515__A1 _02536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06944_ _01989_ _02005_ _02560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09663_ _02419_ _04050_ _04789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06875_ _02502_ _00051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09594_ _03618_ _04726_ _00546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05826_ cpu.spi.busy _01136_ _01490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08614_ _03844_ _03865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08545_ _02467_ _03790_ _03806_ _00417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05757_ cpu.toggle_top\[9\] _01260_ _01261_ _01422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_25_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05188__S0 _00858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05688_ _01167_ _01354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08476_ _03757_ _03758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07427_ cpu.spi.dout\[2\] _02916_ _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_40_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_40_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07358_ _02853_ _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09243__A2 _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06309_ _01962_ _01964_ _01965_ _01966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_07289_ _02546_ _02777_ _02809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09028_ _04167_ _04214_ _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08349__A4 _02431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07006__A1 cpu.toggle_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08004__B _03242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08506__A1 cpu.spi.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output50_I net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07134__I _01352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05740__A1 cpu.timer_capture\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05179__S0 _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04990_ cpu.instr_cycle\[1\] _00689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09524__I _04680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput6 io_in[14] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_108_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06660_ cpu.startup_cycle\[2\] _02313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__09170__A1 _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05611_ _01276_ _01277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07979__I _03370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06591_ _00814_ _01732_ _02247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05542_ _01065_ _01207_ _01129_ _01208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_52_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08330_ _02518_ _03636_ _03638_ _02542_ _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05473_ _00584_ _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_74_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08261_ _03588_ _03590_ _03591_ _00348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_15_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07212_ _01552_ _02761_ _00129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_116_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_89_Left_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08192_ _03496_ _03540_ _03541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_6_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07143_ cpu.regs\[12\]\[1\] _02715_ _02718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_30_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07074_ _02668_ _02671_ _02672_ _00080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06025_ cpu.regs\[12\]\[6\] cpu.regs\[13\]\[6\] cpu.regs\[14\]\[6\] cpu.regs\[15\]\[6\]
+ _00891_ _00893_ _01686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_10_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07976_ _03365_ _03366_ _03342_ _03368_ _03369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_98_Left_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_58_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06927_ _01106_ _01112_ _02543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09715_ _04070_ _02257_ _02553_ _04831_ _04832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09646_ _04760_ _04773_ _04774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_97_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06858_ cpu.timer_capture\[2\] _02471_ _02487_ _02484_ _02488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_2_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05022__I0 cpu.regs\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06789_ _00566_ _02428_ _02429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05809_ net81 _01357_ _01359_ _01473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09577_ cpu.PORTA_DDR\[2\] _04712_ _04713_ _04716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_38_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05911__B net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08528_ _00919_ _03791_ _03795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06793__I _02432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08459_ _02425_ _03743_ _03744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08941__C _04147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06450__A2 _01757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10283_ _00541_ clknet_leaf_13_wb_clk_i cpu.PORTA_DDR\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06033__I _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05961__A1 net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05713__A1 cpu.uart.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07466__A1 cpu.timer_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04951__I _00650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08966__A1 _03885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05095__I3 cpu.regs\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07830_ _03248_ _03250_ _03249_ _03253_ _03254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05627__S1 _01286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08194__A2 _01417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07761_ cpu.uart.div_counter\[4\] _03196_ _00645_ _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06712_ _02364_ _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_09500_ _04664_ _04665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04973_ _00672_ _00673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09143__A1 _02856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07692_ _02640_ _03138_ cpu.uart.div_counter\[8\] _02642_ _03140_ _03141_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_69_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09431_ _04593_ _04609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06643_ _00572_ _02296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09362_ _04550_ _04551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_87_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06574_ _02228_ _02230_ _01931_ _02231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09446__A2 _04571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05525_ _01061_ _01070_ _01191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_63_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08313_ cpu.timer_div_counter\[3\] _03625_ _03627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__05180__A2 _00851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09293_ _03990_ _04487_ _04488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_05456_ _01084_ _01120_ _01122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08244_ _03563_ _03579_ _00343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05387_ _01052_ _01053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08175_ _03521_ cpu.toggle_top\[3\] cpu.toggle_top\[2\] _03523_ _03524_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_15_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07126_ _01679_ cpu.regs\[13\]\[4\] _02698_ _02706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05957__I _01618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_45_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07057_ _02655_ _02652_ cpu.uart.receive_div_counter\[13\] _02632_ _02656_ _02657_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_2_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06008_ _01668_ _01669_ _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09382__A1 _04558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06196__A1 _00810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07232__I1 cpu.regs\[8\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07959_ _03351_ _03348_ _03355_ _03310_ _00282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__05943__A1 _00918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09685__A2 _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09629_ _04546_ _02299_ _02300_ _04757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xwrapped_qcpu_106 io_oeb[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_84_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_84_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08948__A1 _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10266_ _00524_ clknet_leaf_46_wb_clk_i net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10197_ _00455_ clknet_leaf_66_wb_clk_i cpu.last_addr\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05934__A1 cpu.timer_capture\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05107__I cpu.multiplier.a\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08723__I1 cpu.ROM_addr_buff\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09428__A2 _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06290_ _01946_ _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05310_ _00972_ _00977_ _00978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput20 io_in[3] net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_116_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput31 sram_out[5] net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05241_ _00910_ _00911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08939__A1 _04108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05172_ cpu.regs\[4\]\[1\] cpu.regs\[5\]\[1\] cpu.regs\[6\]\[1\] cpu.regs\[7\]\[1\]
+ _00836_ _00839_ _00844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_4_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09980_ _00239_ clknet_leaf_29_wb_clk_i cpu.uart.div_counter\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06414__A2 _02070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08931_ _04107_ _04138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08862_ _00642_ cpu.instr_cycle\[3\] _00689_ _02428_ _04071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__08167__A2 cpu.toggle_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08102__B _03457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07813_ _03232_ _03238_ _03241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08793_ cpu.ROM_addr_buff\[13\] _03991_ _04006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07744_ _03139_ _03181_ _03184_ _03185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_04956_ _00600_ _00655_ _00656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_74_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09667__A2 _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07675_ _03116_ _03118_ _03121_ _03123_ _03124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_67_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06025__S1 _00893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05017__I _00003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09414_ _04594_ _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04887_ cpu.IO_addr_buff\[2\] _00590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_66_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06626_ _01815_ _01936_ _02280_ _02281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_109_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08328__I _03635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09345_ _04531_ _04530_ _04536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06557_ cpu.PC\[5\] _02214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_74_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09276_ _04469_ _04471_ _04472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05508_ cpu.timer_div\[0\] _01174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06488_ _02108_ _02144_ _02145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05439_ _01101_ _01104_ _01105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08227_ _03488_ _03568_ _03569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_1_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05687__I _01352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08158_ cpu.toggle_ctr\[8\] _02608_ _03507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08089_ _03453_ _03449_ _03455_ _00312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_91_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07109_ cpu.regs\[14\]\[6\] _01815_ _02692_ _02695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10120_ _00379_ clknet_leaf_6_wb_clk_i cpu.timer\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10051_ _00310_ clknet_leaf_73_wb_clk_i cpu.orig_PC\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05916__A1 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07669__B2 cpu.uart.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06186__C _01057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07142__I _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05298__I3 cpu.regs\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09594__A1 _03618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06947__A3 _02561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08149__A2 _01512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10249_ _00507_ clknet_leaf_58_wb_clk_i cpu.ROM_spi_cycle\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07761__B _00645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05790_ _01450_ _01451_ _01452_ _01453_ _01454_ _01455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_44_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07460_ _02931_ _02932_ _02940_ _02943_ _02944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XTAP_TAPCELL_ROW_17_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06411_ _02067_ _02065_ _02068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_07391_ _02147_ _02151_ _02885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09130_ _04243_ _04329_ _04330_ _04246_ _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06342_ _01947_ _01944_ _00947_ _01999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09061_ _04247_ _04264_ _04265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08012_ _03001_ _03398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06273_ _01106_ _01112_ _01929_ _01930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_77_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05224_ cpu.regs\[0\]\[2\] cpu.multiplier.a\[2\] cpu.regs\[2\]\[2\] cpu.regs\[3\]\[2\]
+ _00891_ _00893_ _00895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_25_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09585__A1 _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05155_ net75 cpu.ROM_spi_mode _00828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09963_ _00222_ clknet_leaf_37_wb_clk_i cpu.uart.dout\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05086_ _00756_ _00776_ _00778_ _00743_ _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
Xclkbuf_leaf_65_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_65_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08914_ _04075_ _04099_ _04122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09894_ _00153_ clknet_leaf_89_wb_clk_i cpu.regs\[6\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08845_ _01267_ _04049_ _04011_ _04054_ _04055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_08776_ cpu.last_addr\[8\] _03981_ _03994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input12_I io_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07727_ _01899_ _03162_ _03170_ _03161_ _03171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05988_ cpu.toggle_top\[12\] _01258_ _01126_ _01650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__06571__A1 _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_04939_ _00637_ _00638_ _00639_ _00640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07658_ cpu.uart.dout\[6\] _03109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05191__B _00845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07589_ _01872_ _03038_ _02921_ _03050_ _03058_ _03059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_48_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06609_ _02244_ _02250_ _02263_ _02264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09328_ _02317_ _04481_ _04522_ _03722_ _04523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_90_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_80_Left_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09259_ _04206_ _04451_ _04455_ _04456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07846__B _03242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09576__A1 _02525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output80_I net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10103_ _00362_ clknet_leaf_21_wb_clk_i cpu.timer_div_counter\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10034_ _00293_ clknet_leaf_58_wb_clk_i cpu.needs_interrupt vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06562__A1 _02214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06314__A1 _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06617__A2 _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05120__I _00810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06960_ _02569_ _02572_ _02574_ _02575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input4_I io_in[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05911_ _01357_ _01359_ net53 _01574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_72_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06891_ _02496_ _02513_ _02497_ _02515_ _02516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08630_ _00591_ _03861_ _03878_ _03870_ _03879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05842_ cpu.timer_top\[10\] _01242_ _01505_ _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08561_ _02443_ _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05773_ _01436_ _01437_ _01438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08492_ cpu.timer_capture\[14\] _03764_ _03758_ _03771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07512_ _02945_ _02995_ _02996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07443_ cpu.spi.data_in_buff\[7\] _02908_ _02928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_112_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_112_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08058__A1 _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09113_ _04010_ _04303_ _04314_ _04158_ _04315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05231__S _00832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07374_ _00696_ _02869_ _02870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07105__I0 cpu.regs\[14\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06325_ _01980_ _01981_ _01982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_5_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06256_ _01912_ _01913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_88_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09044_ _00661_ _04248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05207_ _00877_ _00878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06187_ _01516_ _01808_ _01844_ _01845_ _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_13_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05138_ _00827_ net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_110_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09946_ _00205_ clknet_leaf_16_wb_clk_i cpu.spi.data_out_buff\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05069_ _00743_ _00755_ _00762_ _00763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09877_ _00136_ clknet_leaf_112_wb_clk_i cpu.regs\[8\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09730__A1 _01963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08497__B _03774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_79_Right_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08828_ _00988_ _01990_ _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08759_ _03966_ _03981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_86_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08297__A1 _02460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_109_Left_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_88_Right_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_118_Left_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06783__A1 _02423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10017_ _00276_ clknet_leaf_33_wb_clk_i cpu.uart.receive_buff\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_97_Right_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_47_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06535__A1 _02105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06110_ _01186_ _01768_ _01769_ _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_81_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07090_ _02384_ _02683_ _02422_ _00085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06041_ net3 _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05785__I _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07992_ cpu.uart.receive_div_counter\[12\] _03366_ _03379_ _03381_ _03382_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06223__B1 cpu.spi.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09800_ _00063_ clknet_leaf_83_wb_clk_i cpu.multiplier.a\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09731_ _04131_ _03436_ _04846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_66_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06774__A1 _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06943_ _02558_ _02559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09662_ _00674_ _01329_ _03835_ _04788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06874_ cpu.timer_capture\[4\] _02494_ _02501_ _02484_ _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09593_ cpu.ROM_spi_mode _04725_ _04726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08613_ _03863_ _03864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05825_ _01487_ _01488_ _01136_ _01489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_89_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08544_ cpu.timer_div\[7\] _03799_ _03802_ _03806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05756_ _01414_ _01416_ _01420_ _01421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05188__S1 _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05687_ _01352_ _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_37_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08475_ _03607_ _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_107_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07426_ _02910_ _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_92_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07240__I _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07357_ _01939_ _01935_ _01932_ _02852_ _02853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_06308_ _01952_ _01963_ _00916_ _01965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__08451__A1 _02998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09027_ _04165_ _04232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_80_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_80_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07288_ _02807_ _02798_ _02808_ _00158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06239_ _01896_ _01897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_103_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07396__B _02851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08203__A1 _00621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06765__A1 _02388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09929_ _00188_ clknet_leaf_44_wb_clk_i cpu.spi.dout\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09703__A1 _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08020__B _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output43_I net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05179__S1 _00839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06296__A3 _00916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08745__A2 _03970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07753__C _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput7 io_in[15] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__04949__I _00648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05610_ _01271_ _01275_ _01276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06590_ _02119_ _02245_ _02246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05541_ _01075_ _01207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08681__A1 _03442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05472_ _00655_ _01042_ _01118_ _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_74_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08260_ cpu.pwm_counter\[0\] cpu.pwm_counter\[1\] cpu.pwm_counter\[2\] _03591_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_80_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08191_ _03506_ _03539_ _03540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07211_ _01469_ _02761_ _00128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07142_ _01468_ _02717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07073_ _02668_ _02671_ _02623_ _02672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_112_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_35_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06024_ _01682_ _01684_ _01685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07975_ _03365_ _03367_ _03368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_58_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09714_ _04045_ _02425_ _02559_ _02562_ _04831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__05270__I1 cpu.multiplier.a\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06926_ _02540_ _02533_ _02541_ _02542_ _00062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09645_ _04729_ _04764_ _04773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06857_ _00906_ _02473_ _02474_ _02486_ _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05808_ _01202_ _01028_ cpu.PORTA_DDR\[2\] _01472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_2_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06788_ _00582_ _02428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_38_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09576_ _02525_ _04711_ _04715_ _00539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_92_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05739_ _01394_ _01399_ _01403_ _01404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08527_ _02614_ _03793_ _03794_ _00411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08458_ _03741_ _03743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_74_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05486__A1 _01151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07409_ net20 _02855_ _02901_ _02902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_107_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08389_ cpu.timer_capture\[4\] _03678_ _03685_ _03257_ _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_46_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05639__B _01304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06986__A1 _02597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10282_ _00540_ clknet_leaf_103_wb_clk_i cpu.PORTA_DDR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06738__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07346__S _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07145__I _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08663__A1 _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05477__A1 _01137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_114_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09535__I _04680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_119_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07760_ cpu.uart.div_counter\[4\] _03195_ _03190_ _03197_ _03198_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_04972_ cpu.instr_buff\[14\] _00672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06711_ _02363_ _02364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07055__I cpu.uart.divisor\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09430_ _04595_ _04607_ _04608_ _00500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07691_ _02640_ _03138_ _03139_ cpu.uart.divisor\[0\] _03140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_79_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05004__I1 _00700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06642_ _02294_ _02295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06894__I _02426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06901__A1 _02518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09361_ _04549_ cpu.startup_cycle\[0\] _04550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_63_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06573_ net1 _02229_ _02230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09292_ cpu.last_addr\[6\] cpu.last_addr\[5\] cpu.last_addr\[4\] _04486_ _04487_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_05524_ _01068_ _01078_ _01128_ _01190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
Xclkbuf_leaf_19_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_19_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_63_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08312_ _03622_ _03625_ _03626_ _00364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_19_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08243_ _03499_ _03578_ _03579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05455_ _01087_ _01120_ _01121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_62_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05386_ _01047_ _01051_ _01052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08174_ _03522_ _03523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07125_ _01616_ _02699_ _02705_ _00098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07056_ cpu.uart.receive_div_counter\[4\] cpu.uart.divisor\[4\] _02656_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_88_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06968__A1 _02186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06007_ _00944_ _00942_ _01669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_7_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05079__S0 _00770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07958_ cpu.uart.receive_div_counter\[5\] _03345_ _03354_ _03355_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_97_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07889_ cpu.uart.data_buff\[8\] _03260_ _03301_ _03302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06909_ cpu.timer_top\[3\] _02521_ _02530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xwrapped_qcpu_107 io_out[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09628_ _04755_ _02302_ _04756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09180__I _04071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09559_ _04695_ _04704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08645__A1 _02421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05003__S0 _00697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05213__I _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10265_ _00523_ clknet_leaf_49_wb_clk_i net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10196_ _00454_ clknet_leaf_65_wb_clk_i cpu.last_addr\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06187__A2 _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09125__A2 _04273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07136__A1 _01114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08884__A1 _04042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput10 io_in[18] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput21 io_in[6] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__04962__I _00661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05240_ _00909_ _00910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput32 sram_out[6] net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_109_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05171_ _00842_ _00843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_24_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08930_ _04101_ _04137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08861_ _04069_ _04070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07812_ cpu.uart.div_counter\[14\] _03239_ _03240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08792_ cpu.last_addr\[13\] _03996_ _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07743_ _03177_ _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04955_ cpu.br_rel_dest\[4\] _00655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07674_ _02655_ _03122_ cpu.uart.div_counter\[13\] _02632_ _03123_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_04886_ _00588_ _00589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08609__I _03370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09413_ _04593_ _04594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06625_ _02259_ _02279_ _02280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09344_ _01909_ _04531_ _04530_ _04535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06556_ cpu.PC\[6\] _02213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08627__B2 _00958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09275_ _04197_ _04459_ _04470_ _04199_ _04471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_62_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05507_ _01172_ _01173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06487_ _02110_ _02144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_117_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05438_ _01103_ _01104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08226_ _03555_ _03567_ _03568_ _00336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_7_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08157_ cpu.toggle_ctr\[14\] _03504_ _03505_ cpu.toggle_ctr\[13\] _03506_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_70_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05369_ _01033_ _01034_ _01007_ _01035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07108_ _01753_ _02687_ _02694_ _00092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08088_ cpu.orig_PC\[6\] _03454_ _03447_ _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07039_ cpu.uart.receive_div_counter\[1\] _02639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_31_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10050_ _00309_ clknet_leaf_63_wb_clk_i cpu.orig_PC\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05208__I cpu.base_address\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08866__A1 _00637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05224__S0 _00891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_111_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10248_ _00506_ clknet_leaf_59_wb_clk_i cpu.ROM_spi_cycle\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07357__A1 _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10179_ _00437_ clknet_leaf_78_wb_clk_i cpu.base_address\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08857__A1 _03836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06410_ _00914_ _02017_ _02066_ _00953_ _02067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_45_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07390_ _02203_ _02883_ _02884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06341_ _00954_ _00946_ _01950_ _01998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09060_ _04248_ _04255_ _04263_ _04264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_60_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06272_ _01148_ _01928_ _01929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08011_ cpu.had_int _03396_ cpu.needs_interrupt _03397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05223_ cpu.regs\[4\]\[2\] cpu.regs\[5\]\[2\] cpu.regs\[6\]\[2\] cpu.regs\[7\]\[2\]
+ _00891_ _00893_ _00894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__09034__A1 _02570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05154_ cpu.PORTB_DDR\[2\] net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XTAP_TAPCELL_ROW_77_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09962_ _00221_ clknet_leaf_38_wb_clk_i cpu.spi.data_in_buff\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05085_ _00759_ _00777_ _00778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08913_ _04109_ _04114_ _04120_ _04113_ _04121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09893_ _00152_ clknet_leaf_86_wb_clk_i cpu.regs\[6\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07348__A1 cpu.regs\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07952__B _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08844_ _02418_ _00667_ _04054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08775_ _03990_ _03970_ _03992_ _03993_ _00460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05987_ cpu.toggle_top\[4\] _01253_ _01259_ _01649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07726_ _01899_ _03169_ _03170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_34_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_34_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_04938_ _00613_ _00639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06571__A2 _02227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08339__I _03635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04869_ cpu.startup_cycle\[1\] cpu.startup_cycle\[0\] _00572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07657_ _03107_ _03101_ _03108_ _03104_ _00227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_67_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07588_ _01872_ _01879_ _03052_ _03058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_48_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06608_ _02239_ _02249_ _02263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09327_ _04482_ _04484_ _04521_ _04522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_62_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06539_ _02192_ _02195_ _02196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09258_ _04374_ _04437_ _04454_ _04404_ _04007_ _04455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09189_ _04386_ _04387_ _04388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08209_ _03472_ cpu.toggle_ctr\[0\] cpu.toggle_ctr\[1\] _03557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07036__B1 _01583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output73_I net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10102_ _00361_ clknet_leaf_103_wb_clk_i cpu.pwm_top\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10033_ _00292_ clknet_leaf_30_wb_clk_i cpu.uart.receive_div_counter\[15\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05910_ _01108_ _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06890_ _02514_ _02499_ _02515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05841_ _01248_ _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08560_ _03815_ _03817_ _03819_ _00419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05772_ _00726_ _01437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07511_ _02947_ _02969_ _02988_ _02994_ _02995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08491_ _03729_ _03761_ _03769_ _03770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07502__A1 cpu.timer_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07442_ cpu.spi.dout\[7\] _02916_ _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07373_ _02853_ _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09112_ cpu.orig_PC\[7\] _03854_ _04314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06324_ _00902_ _00896_ _00925_ _00929_ _00887_ _01950_ _01981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_29_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07105__I1 _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05116__I0 cpu.regs\[12\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05311__I _00978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06255_ cpu.mem_cycle\[1\] _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09043_ _04243_ _04242_ _04245_ _04246_ _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_111_Right_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05292__A2 _00960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05206_ _00876_ _00877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06186_ _01140_ _01268_ _01273_ _01057_ _01845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__05131__I3 cpu.regs\[11\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05137_ _00826_ _00827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09945_ _00204_ clknet_leaf_21_wb_clk_i cpu.spi.data_out_buff\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05068_ _00756_ _00758_ _00761_ _00743_ _00762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_09876_ _00135_ clknet_leaf_112_wb_clk_i cpu.regs\[8\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08827_ _01107_ _01942_ _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08758_ cpu.last_addr\[4\] _03980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08689_ _03925_ _00442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09494__A1 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07709_ _00621_ _03157_ _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08297__A2 _03613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09246__A1 _03469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05221__I _00837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07280__I0 _02753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06783__A2 _02413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10016_ _00275_ clknet_leaf_34_wb_clk_i cpu.uart.receive_buff\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07732__A1 _03007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09485__A1 cpu.pwm_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06040_ _01055_ _01699_ _01700_ _01701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_clkbuf_leaf_25_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07991_ _02658_ _03380_ _03352_ _03381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06942_ _01619_ _01006_ _01043_ _02558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_09730_ _01963_ _04837_ _04845_ _00563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09661_ _04778_ _04784_ _04787_ _03993_ _00552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09206__C _04321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06873_ _02495_ _02496_ _02497_ _02500_ _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09592_ _04600_ _02297_ _02298_ _02302_ _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_08612_ _03840_ _03863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05824_ cpu.uart.dout\[2\] _00616_ _01488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09476__A1 _04558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08543_ _03804_ _03790_ _03805_ _00416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05755_ _01419_ _01420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_82_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05686_ _01351_ _01352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08474_ cpu.timer\[11\] _03742_ _03755_ _03756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07425_ _02912_ _02913_ _02915_ _00188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_64_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09228__B2 _04162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07356_ _02851_ _02852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07287_ cpu.regs\[6\]\[7\] _02801_ _02808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06307_ _01963_ _01948_ _01964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_32_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09026_ _04176_ _04214_ _04230_ _04202_ _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06238_ _01175_ _01895_ _01896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_17_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06169_ cpu.uart.divisor\[15\] _01382_ _01827_ _00012_ _01828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_13_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08203__A2 _03551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09928_ _00187_ clknet_leaf_39_wb_clk_i cpu.spi.dout\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09859_ _00118_ clknet_leaf_112_wb_clk_i cpu.regs\[11\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09467__A1 _03079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output36_I net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06205__A1 _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_109_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput8 io_in[16] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05540_ _01183_ _01186_ _01187_ _01205_ _01206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_59_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08130__A1 cpu.toggle_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05471_ _01060_ _01137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_52_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08190_ _03491_ _03537_ _03538_ _03539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07210_ _01353_ _02761_ _00127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07141_ _02710_ _02714_ _02716_ _00103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07072_ cpu.uart.receive_counter\[1\] _02669_ _02671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06023_ _00832_ _01683_ _00845_ _01684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_2_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07944__A1 _02662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07974_ _02650_ _03360_ _03367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_58_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09713_ _01868_ _04821_ _04830_ _00561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06925_ _02523_ _02542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09644_ _02360_ _04771_ _02346_ _04772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06856_ cpu.timer\[2\] _02475_ _02486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08775__C _03993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05807_ _01270_ _01471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_2_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05022__I2 _00715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05036__I _00717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06787_ _02426_ _02427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_38_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09575_ cpu.PORTA_DDR\[1\] _04712_ _04713_ _04715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05738_ cpu.timer_div\[1\] _01400_ _01402_ _01403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08526_ cpu.timer_div\[1\] _03791_ _03774_ _03794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07251__I _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05669_ _01333_ _01335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08457_ _03741_ _03742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_37_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05486__A2 _01145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07408_ _02852_ _02900_ _02901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08388_ _02976_ _03679_ _03681_ _03683_ _03684_ _03685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_07339_ cpu.regs\[3\]\[1\] _02840_ _02842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09009_ _04213_ _04214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10281_ _00539_ clknet_leaf_13_wb_clk_i cpu.PORTA_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08360__A1 cpu.timer_capture\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05174__A1 _00843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08112__A1 _02254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04921__A1 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05477__A2 _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06977__A2 _02589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06729__A2 _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07336__I _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06240__I _01888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04971_ _00607_ _00671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06710_ _00691_ _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07690_ cpu.uart.div_counter\[0\] _03139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_69_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06641_ _00571_ _02294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09360_ _04548_ _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_06572_ _01907_ _01040_ _01921_ _02229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__05960__I0 net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09291_ cpu.last_addr\[3\] _04485_ _04486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_05523_ _01188_ _01189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_87_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08311_ cpu.timer_div_counter\[0\] cpu.timer_div_counter\[1\] cpu.timer_div_counter\[2\]
+ _03626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_63_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_35_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05454_ _00595_ _00605_ _01002_ _01117_ _01120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_74_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08242_ _03562_ _03577_ _03578_ _00342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xclkbuf_leaf_59_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_59_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_62_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05385_ _00991_ _01050_ _01051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08173_ cpu.toggle_ctr\[2\] _03522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07124_ cpu.regs\[13\]\[3\] _02703_ _02705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07055_ cpu.uart.divisor\[14\] _02655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_15_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06006_ _00938_ _00940_ _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07957_ _03352_ _03353_ _03354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06908_ _02450_ _02529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07888_ _02513_ _03236_ _03301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08342__A1 cpu.timer_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09627_ _04566_ _04560_ _04755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06839_ _02470_ _02471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xwrapped_qcpu_108 io_out[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__08077__I _03410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09558_ _04695_ _04703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08509_ _02529_ _03777_ _03782_ _00405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_108_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05003__S1 _00698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09489_ cpu.pwm_top\[1\] _03586_ _04654_ cpu.pwm_top\[2\] _04655_ _04656_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_93_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08805__I _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Left_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08026__B _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10264_ _00522_ clknet_leaf_46_wb_clk_i net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10195_ _00453_ clknet_leaf_65_wb_clk_i cpu.last_addr\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_21_Left_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07136__A2 _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08333__A1 cpu.timer_top\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08884__A2 _04091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06895__A1 _01031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput11 io_in[19] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput22 io_in[7] net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput33 sram_out[7] net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_12_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05170_ _00006_ _00842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08860_ cpu.PC\[0\] _04069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08572__A1 _02648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07811_ _03157_ _03236_ _03238_ _03239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_106_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_106_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08791_ _00686_ _04003_ _04004_ _00465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07742_ _03179_ _03183_ _02930_ _00237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_04954_ _00653_ cpu.br_rel_dest\[6\] _00654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07673_ cpu.uart.div_counter\[14\] _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_04885_ _00585_ _00587_ _00588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09412_ _02348_ _04592_ _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06886__A1 cpu.timer_capture\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06624_ net19 _02229_ _02276_ _02278_ _02279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09343_ _04534_ _00487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06555_ cpu.PC\[7\] _02212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08627__A2 _03864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09274_ cpu.orig_PC\[13\] _03863_ _04470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05506_ _01089_ _01172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06486_ _02139_ _02142_ _02143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06638__A1 _02283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05437_ _01102_ _01103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08225_ _03530_ _03566_ _03568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_99_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05368_ cpu.br_rel_dest\[6\] _01034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08156_ cpu.toggle_top\[13\] _03505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07063__A1 cpu.uart.divisor\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07107_ cpu.regs\[14\]\[5\] _02685_ _02694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08087_ _03400_ _03454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05299_ _00965_ _00966_ _00967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_113_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07038_ _02448_ _02638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_11_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08989_ _01573_ _04188_ _04193_ _04194_ _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_98_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08866__A2 _01115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05224__S1 _00893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08963__C _04169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06764__B _02406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_4_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_4_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_21_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10247_ _00505_ clknet_leaf_61_wb_clk_i cpu.ROM_spi_dat_out\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10178_ _00436_ clknet_leaf_81_wb_clk_i cpu.base_address\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_89_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06580__A3 _01118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05540__A1 _01183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06340_ _01940_ _01996_ _01997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_29_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06271_ _01154_ _01164_ _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08010_ net17 _03396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05222_ _00892_ _00893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_52_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07045__A1 _02640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05153_ cpu.PORTB_DDR\[1\] net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_77_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09961_ _00220_ clknet_leaf_38_wb_clk_i cpu.spi.data_in_buff\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05084_ cpu.regs\[12\]\[4\] cpu.regs\[13\]\[4\] cpu.regs\[14\]\[4\] cpu.regs\[15\]\[4\]
+ _00749_ _00750_ _00777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_110_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08912_ _04116_ _04118_ _04119_ _04120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08545__A1 _02467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09892_ _00151_ clknet_leaf_86_wb_clk_i cpu.regs\[6\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08843_ _02418_ _04048_ _04050_ _04052_ _04053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_08774_ _03159_ _03993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05986_ _01643_ _01645_ _01647_ _01648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07725_ _03009_ cpu.spi.counter\[1\] _01900_ _03169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_04937_ _00606_ _00638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_88_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08848__A2 _00919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07656_ cpu.uart.receive_buff\[5\] _03102_ _03108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_04868_ _00567_ _00568_ _00569_ _00570_ _00571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_07587_ _01903_ _03057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_74_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_74_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_75_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06607_ _02242_ _02260_ _02261_ _02262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09326_ _04520_ _04521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06538_ _02194_ _02195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09257_ _00769_ _04452_ _04453_ _04454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_106_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08208_ cpu.toggle_clkdiv cpu.toggle_ctr\[1\] cpu.toggle_ctr\[0\] _03556_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_16_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06469_ _02125_ _02122_ _02126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_105_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09188_ cpu.PC\[10\] _00876_ _04387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_31_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08139_ cpu.toggle_ctr\[7\] _03488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_43_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08784__A1 cpu.ROM_addr_buff\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08090__I _02455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05598__A1 _00637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10101_ _00360_ clknet_leaf_3_wb_clk_i cpu.pwm_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output66_I net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08536__A1 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05219__I _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10032_ _00291_ clknet_leaf_33_wb_clk_i cpu.uart.receive_div_counter\[14\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_4_0_wb_clk_i clknet_0_wb_clk_i clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_14_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_15_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05133__S0 _00816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08527__A1 _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05840_ _01247_ _01503_ _01504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05771_ _01435_ _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_49_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07510_ _02951_ _02966_ _02992_ _02993_ _02994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_77_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07280__S _02796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08490_ _03743_ _02508_ _03769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07441_ _02925_ _02911_ _02926_ _00694_ _00193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_clkbuf_leaf_54_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07372_ _02867_ _01351_ _01931_ _02868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09111_ _04248_ _04312_ _04313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07266__A1 _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06323_ _01944_ _01980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_29_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05116__I1 cpu.regs\[13\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06254_ _01908_ _01910_ _01911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09042_ _04106_ _04246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05205_ cpu.base_address\[2\] _00876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06185_ _01840_ _01841_ _01843_ _01844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07018__A1 _02460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05136_ _00797_ _00820_ _00825_ _00826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_40_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09944_ _00203_ clknet_leaf_21_wb_clk_i cpu.spi.data_out_buff\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08518__A1 cpu.spi.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05067_ _00759_ _00760_ _00761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09875_ _00134_ clknet_leaf_95_wb_clk_i cpu.regs\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08826_ _04027_ _04033_ _04035_ _04036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_93_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08757_ _03972_ _03978_ _03979_ _00456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05969_ cpu.uart.divisor\[12\] _01484_ _00616_ _01631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08688_ _03924_ cpu.ROM_addr_buff\[3\] _03921_ _03925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07708_ _03156_ _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07639_ cpu.uart.receive_buff\[0\] _03095_ _03096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_83_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09309_ cpu.last_addr\[6\] _04503_ _04504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_91_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07009__A1 _02447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10214__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08509__A1 _02529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07280__I1 cpu.regs\[6\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10015_ _00274_ clknet_leaf_34_wb_clk_i cpu.uart.receive_buff\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05743__A1 _01407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_4_Left_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07767__C _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07990_ _03376_ _03372_ _03380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06941_ _02556_ _02218_ _02557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09660_ _04778_ _04786_ net77 _04787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05982__A1 cpu.timer_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08611_ _03837_ _03862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06872_ _02498_ _02499_ _02500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05823_ _01485_ _01486_ _01142_ _01487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05734__A1 cpu.spi.dout\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09591_ _02540_ _04718_ _04724_ _00545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_85_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08542_ cpu.timer_div\[6\] _03799_ _03802_ _03805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05754_ _01417_ _01418_ _01172_ _01419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08473_ _02489_ _03751_ _03755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07424_ _02914_ _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_59_Left_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05685_ _01308_ _01350_ _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08119__B _03467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07355_ _02393_ _01906_ _02850_ _02851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__07239__A1 _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07286_ _01868_ _02807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06306_ _01945_ _01963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_33_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09025_ _04223_ _04227_ _04229_ _04230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06237_ _00642_ _00669_ _01895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_5_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06168_ _01818_ _01375_ _01696_ _01826_ _01382_ _01827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_40_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_68_Left_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05119_ _00797_ _00803_ _00809_ _00810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_06099_ _01758_ _01759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09927_ _00186_ clknet_leaf_83_wb_clk_i cpu.regs\[2\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06102__B net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08911__A1 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09858_ _00117_ clknet_leaf_114_wb_clk_i cpu.regs\[11\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08809_ cpu.IE _04015_ _04020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09789_ _00052_ clknet_leaf_7_wb_clk_i cpu.timer_capture\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_77_Left_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09219__A2 _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06150__B2 _00811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06150__A1 _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05964__A1 _01621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput9 io_in[17] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05470_ _01135_ _01136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05142__I cpu.PORTA_DDR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09549__I _04674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07140_ cpu.regs\[12\]\[0\] _02715_ _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07071_ _02668_ _02670_ _02365_ _00079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06022_ cpu.regs\[0\]\[6\] cpu.multiplier.a\[6\] cpu.regs\[2\]\[6\] cpu.regs\[3\]\[6\]
+ _00835_ _00969_ _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_23_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09394__A1 _02478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07973_ _03308_ _03366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09712_ cpu.regs\[9\]\[7\] _04824_ _04830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05270__I3 cpu.regs\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06924_ cpu.timer_top\[7\] _02534_ _02541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09643_ _04760_ _04762_ _04770_ _04730_ _04771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06855_ _02485_ _00048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05806_ _01168_ _01469_ _01470_ _00014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09574_ _02518_ _04711_ _04714_ _00538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08525_ _03789_ _03793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06786_ _02425_ _02426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05183__A2 _00854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05737_ _01401_ _01402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06148__I _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06132__A1 _01790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05668_ _00711_ _01333_ _01334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_18_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08456_ _01225_ _03741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07880__A1 _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07407_ _02897_ _02899_ _02900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08387_ _03651_ _03684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05599_ _01057_ _01264_ _01265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07338_ _01352_ _02839_ _02841_ _00175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07269_ _02796_ _02797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09008_ _02216_ _04212_ _04213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10280_ _00538_ clknet_leaf_99_wb_clk_i cpu.PORTA_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__06199__A1 _00826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05946__A1 _00905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07699__A1 _02648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07699__B2 _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_85_Left_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08538__I _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04921__A2 _00622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08112__A2 _03404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06123__A1 cpu.timer_capture\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05477__A3 _01142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_94_Left_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05937__A1 cpu.timer_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04970_ _00666_ _00669_ _00670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05137__I _00826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06640_ _01934_ _02292_ _02293_ _00025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06362__B2 _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05960__I1 cpu.PORTA_DDR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04912__A2 _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06571_ _01923_ _02227_ _02228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09290_ cpu.last_addr\[2\] cpu.last_addr\[1\] cpu.last_addr\[0\] _04485_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__06114__A1 _00615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05522_ _01016_ _01084_ _01188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08310_ cpu.timer_div_counter\[0\] cpu.timer_div_counter\[1\] cpu.timer_div_counter\[2\]
+ _03625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_63_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05453_ _01003_ _01118_ _01119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08241_ cpu.toggle_ctr\[12\] _03576_ _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_6_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05384_ _01049_ _01050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08172_ _03519_ _03521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08183__I cpu.toggle_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07123_ _01552_ _02699_ _02704_ _00097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07054_ _02649_ cpu.uart.receive_div_counter\[12\] _02650_ _02642_ _02653_ _02654_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
Xclkbuf_leaf_99_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_99_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_28_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_28_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06005_ net94 _00949_ _01456_ _01667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_7_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05928__A1 cpu.spi.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07956_ _03351_ _03348_ _03353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input28_I sram_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06907_ _02527_ _02520_ _02528_ _02524_ _00057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05047__I _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_106_Right_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07887_ _03291_ _03299_ _03300_ _00265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09626_ net78 _04754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_97_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06838_ _01061_ _01077_ _02469_ _02470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xwrapped_qcpu_109 io_out[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_06769_ _02393_ _02411_ _02412_ _02371_ _02413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_09557_ _02529_ _04696_ _04702_ _00533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06105__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08508_ cpu.spi.divisor\[3\] _03778_ _03782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09488_ cpu.pwm_top\[3\] cpu.pwm_counter\[3\] _04655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_38_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08439_ _03608_ _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output96_I net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10263_ _00521_ clknet_leaf_42_wb_clk_i net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10194_ _00452_ clknet_leaf_69_wb_clk_i cpu.ROM_addr_buff\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06967__I0 _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08708__I1 cpu.ROM_addr_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06592__A1 _02009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09530__A1 _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06895__A2 _02433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput12 io_in[1] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput23 io_in[8] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09349__A1 _03057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08790_ cpu.ROM_addr_buff\[12\] _03991_ _04004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07810_ _03180_ _03237_ _03238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07741_ _03139_ _03182_ _03183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09521__A1 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04953_ _00652_ _00653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_07672_ cpu.uart.divisor\[15\] _03119_ cpu.uart.div_counter\[14\] _03120_ _03121_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_04884_ _00586_ _00587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09411_ _02366_ _02345_ _04591_ _04592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06623_ _01927_ _02277_ _02278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09342_ _04531_ _04481_ _04533_ _04527_ _04534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_90_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06554_ cpu.PC\[8\] _02211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_118_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05505_ _01086_ _01171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09273_ _04462_ _04468_ _04346_ _04469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06485_ _02033_ _02141_ _02142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05436_ _00618_ _00583_ _01095_ _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_08224_ _03530_ _03566_ _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_28_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05367_ _00653_ _01033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08155_ cpu.toggle_top\[14\] _03504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07106_ _02693_ _00091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08086_ _03452_ _03453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05298_ cpu.regs\[0\]\[5\] cpu.multiplier.a\[5\] cpu.regs\[2\]\[5\] cpu.regs\[3\]\[5\]
+ _00898_ _00899_ _00966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_07037_ _02628_ _02629_ _02630_ _02448_ _02636_ _02637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_11_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08988_ _04154_ _04194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07939_ cpu.uart.receive_div_counter\[1\] _03328_ _03339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09609_ cpu.ROM_addr_buff\[0\] _04738_ _04739_ _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08866__A3 _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08079__A1 _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07126__I0 _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06780__B _00685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07595__C _02506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10246_ _00504_ clknet_leaf_61_wb_clk_i cpu.ROM_spi_dat_out\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08554__A2 _03813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07357__A3 _01932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10177_ _00435_ clknet_leaf_78_wb_clk_i cpu.base_address\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_89_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09503__A1 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_44_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04879__A1 net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07293__A2 _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06270_ _01923_ _01926_ _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_114_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05221_ _00837_ _00892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_25_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05152_ cpu.PORTB_DDR\[0\] net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_80_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08461__I _03739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09960_ _00219_ clknet_leaf_41_wb_clk_i cpu.spi.data_in_buff\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05083_ _00775_ _00776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_40_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07077__I _02456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08911_ _01430_ _04115_ _04119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09742__A1 _03442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09891_ _00150_ clknet_leaf_90_wb_clk_i cpu.regs\[7\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07805__I _02390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08842_ _02070_ _04051_ _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_83_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08773_ cpu.ROM_addr_buff\[7\] _03991_ _03992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05985_ _01646_ _01647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07724_ _02440_ _03168_ _00233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04936_ _00636_ _00637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06308__A1 _01952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07655_ cpu.uart.dout\[5\] _03107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_88_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_04867_ cpu.ROM_spi_cycle\[3\] cpu.ROM_spi_cycle\[2\] _00570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_67_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06606_ _02238_ _02252_ _02261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XPHY_EDGE_ROW_40_Left_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07586_ _01879_ _03052_ _03054_ _03056_ _00208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_48_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09325_ _04493_ _04495_ _04519_ _04520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06537_ _01969_ _02170_ _02193_ _02194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09256_ _04452_ _04437_ _04453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06468_ _02097_ _02123_ _02124_ _02125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__08481__A1 _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06156__I _01815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_43_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_43_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_105_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05419_ _01030_ _01084_ _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_63_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08207_ _03552_ _03555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09187_ cpu.PC\[10\] _00876_ _04386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06399_ _02046_ _02054_ _02055_ _02056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_99_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08138_ _02467_ _03481_ _03487_ _00329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08069_ _03439_ _03434_ _03440_ _00307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10100_ _00359_ clknet_leaf_3_wb_clk_i cpu.pwm_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10031_ _00290_ clknet_leaf_30_wb_clk_i cpu.uart.receive_div_counter\[13\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09733__A1 _01942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output59_I net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05235__I _00905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08775__A2 _03970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05133__S1 _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09724__A1 _04043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10229_ _00487_ clknet_leaf_56_wb_clk_i cpu.mem_cycle\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_72_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05770_ _01434_ _01435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_0_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05145__I cpu.PORTB_DDR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07440_ cpu.spi.data_in_buff\[6\] _02921_ _02926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08456__I _01225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07371_ net1 _02855_ _02866_ _02867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09110_ _02423_ _04188_ _04311_ _04194_ _04312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06322_ _01977_ _01978_ _01979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09041_ cpu.orig_PC\[5\] _04244_ _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07266__A2 _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06253_ _01909_ _01910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_13_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05204_ _00875_ net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06184_ _00650_ _01057_ _01273_ _01173_ _01842_ _01843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_102_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05135_ _00804_ _00822_ _00824_ _00797_ _00825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__06777__A1 _02419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09943_ _00202_ clknet_leaf_18_wb_clk_i cpu.spi.data_out_buff\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05066_ cpu.regs\[12\]\[3\] cpu.regs\[13\]\[3\] cpu.regs\[14\]\[3\] cpu.regs\[15\]\[3\]
+ _00752_ _00753_ _00760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05764__B _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09874_ _00133_ clknet_leaf_97_wb_clk_i cpu.regs\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09715__A1 _04070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08825_ _04034_ _01937_ _04035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input10_I io_in[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08756_ cpu.ROM_addr_buff\[3\] _03976_ _03979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05968_ _01375_ _01627_ _01629_ _01630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08687_ _03446_ _03917_ _03923_ _03924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07707_ _03154_ _03155_ _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04919_ _00620_ _00621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_05899_ _01555_ _01559_ _01561_ _01562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06701__A1 cpu.ROM_addr_buff\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07638_ _03092_ _03095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07270__I _02796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07569_ _03028_ _03040_ _03042_ _00205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05060__S0 _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09308_ cpu.last_addr\[5\] _03980_ _04486_ _04503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_63_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09239_ _04433_ _04435_ _04436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10014_ _00273_ clknet_leaf_35_wb_clk_i cpu.uart.receive_buff\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07445__I _02929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08142__B1 cpu.toggle_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_27_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_75_Right_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06208__B1 _01866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08879__C _00657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_105_Left_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06940_ _02216_ _02556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input2_I io_in[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06871_ _02472_ _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05822_ cpu.uart.divisor\[10\] _01484_ _01486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08610_ _03857_ _03861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07184__A1 _02684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_84_Right_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09570__I _04710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09590_ cpu.PORTA_DDR\[7\] _04719_ _04720_ _04724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08541_ _02462_ _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_49_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05753_ _01086_ _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05684_ net26 _01310_ _01311_ _01349_ _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_49_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08472_ _03740_ _03753_ _03754_ _00396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07423_ _00692_ _02914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_114_Left_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07354_ _02324_ _02319_ _02395_ _02850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_85_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05759__B _00904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07285_ _02806_ _00157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06305_ _01961_ _01958_ _01962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06236_ _01893_ _01894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_93_Right_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09024_ _04010_ _04214_ _04228_ _04158_ _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06998__A1 _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06167_ net14 _01121_ _01823_ _01825_ _01826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06098_ _01757_ _01758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05118_ _00804_ _00806_ _00808_ _00797_ _00809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_05049_ _00713_ _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09926_ _00185_ clknet_leaf_83_wb_clk_i cpu.regs\[2\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09857_ _00116_ clknet_leaf_115_wb_clk_i cpu.regs\[11\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08808_ _04016_ _04019_ _03395_ _00467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09788_ _00051_ clknet_leaf_7_wb_clk_i cpu.timer_capture\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06922__A1 _02538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08739_ _02331_ _03964_ _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08675__A1 _03439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09155__A2 _04273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05272__S0 _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08666__A1 _00911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07070_ cpu.uart.receive_counter\[0\] _02667_ _02669_ _02670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_54_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05652__A1 _00908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06021_ _00842_ _01681_ _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_30_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07972_ cpu.uart.receive_div_counter\[9\] _03365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09711_ _04829_ _00560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06923_ _02466_ _02540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09642_ _04520_ _04769_ _04770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06854_ cpu.timer_capture\[1\] _02471_ _02482_ _02484_ _02485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06904__A1 _02525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06785_ _01356_ _02425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09573_ cpu.PORTA_DDR\[0\] _04712_ _04713_ _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05805_ cpu.regs\[15\]\[1\] _01354_ _01470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08524_ _01174_ _03790_ _03792_ _03648_ _00410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05736_ _01025_ _00997_ _01062_ _01401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_26_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05667_ _00864_ _00869_ _01333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08455_ _03739_ _03740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05598_ _00637_ _01263_ _01264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08386_ _02498_ _03682_ _03683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_46_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07406_ _01926_ _02223_ _02898_ _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_18_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07337_ cpu.regs\[3\]\[0\] _02840_ _02841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07268_ _02795_ _02796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_103_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06219_ _01875_ cpu.spi.divisor\[4\] _01876_ cpu.spi.div_counter\[7\] _01877_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09007_ _03445_ _04132_ _04212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07199_ _02754_ _00123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_103_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09909_ _00168_ clknet_leaf_86_wb_clk_i cpu.regs\[4\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09424__B _04603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08896__A1 _04043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output41_I net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05254__S0 _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08648__A1 _03885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06783__B _00685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_3_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06802__I cpu.uart.divisor\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06023__B _00845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05153__I cpu.PORTB_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08639__B2 _01733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06570_ _01939_ _02201_ _02202_ _02226_ _02227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__09300__A2 cpu.ROM_addr_buff\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05521_ net6 _01053_ _01185_ _01187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_87_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07311__A1 _02807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04992__I net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05452_ _01117_ _01118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_74_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08240_ cpu.toggle_ctr\[12\] _03576_ _03577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08171_ cpu.toggle_ctr\[4\] _03517_ _03518_ _03519_ _03520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_27_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05383_ cpu.IO_addr_buff\[3\] _01048_ _01049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07122_ cpu.regs\[13\]\[2\] _02703_ _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07053_ _02651_ cpu.uart.receive_div_counter\[15\] _02652_ cpu.uart.divisor\[14\]
+ _02653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_88_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_93_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06004_ _00878_ _01665_ _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_11_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_68_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_68_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07955_ _03330_ _03352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06906_ cpu.timer_top\[2\] _02521_ _02528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09625_ _03618_ _04753_ _00550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07543__I _01897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07886_ cpu.uart.data_buff\[8\] _03288_ _03289_ _03300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_37_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06837_ _01063_ _02432_ _02469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07550__A1 _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06768_ _02333_ _02411_ _02412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09556_ cpu.PORTB_DDR\[3\] _04697_ _04698_ _04702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06699_ cpu.ROM_spi_dat_out\[7\] _02351_ _02352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05719_ _01379_ _01383_ _00012_ _01384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08507_ _02527_ _03777_ _03781_ _00404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09487_ _03589_ _04654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_38_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08438_ cpu.timer\[13\] _03692_ _03656_ _03725_ _03726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_92_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05864__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09055__A1 _02570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08369_ _03654_ _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08802__A1 _04007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10262_ _00520_ clknet_leaf_42_wb_clk_i net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA_output89_I net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10193_ _00451_ clknet_leaf_70_wb_clk_i cpu.ROM_addr_buff\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09154__B _04324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_34_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08284__I _03607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05855__A1 _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput13 io_in[20] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput24 io_in[9] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_12_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05148__I cpu.PORTA_DDR\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_73_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07740_ _03181_ _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04952_ cpu.br_rel_dest\[7\] _00652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_74_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07671_ _02655_ _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07532__A1 _02427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04883_ cpu.IO_addr_buff\[0\] _00586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09410_ _04555_ _04589_ _04590_ _04591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06622_ _02262_ _02275_ _02277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09341_ _04482_ _04521_ _04532_ _04533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06553_ _02209_ _02210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_114_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05504_ _01155_ _01170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06707__I _02359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09272_ _04340_ _04466_ _04467_ _04468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_74_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_115_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_115_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06484_ _02065_ _02140_ _02141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__05846__A1 cpu.toggle_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09037__A1 _02570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05435_ _01034_ _01101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_7_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08223_ cpu.toggle_ctr\[5\] cpu.toggle_ctr\[4\] _03559_ _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_99_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05366_ _01027_ _01031_ _01032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08154_ _03496_ _03498_ _03502_ _03503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_70_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08085_ cpu.PC\[6\] _03452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07105_ cpu.regs\[14\]\[4\] _01678_ _02692_ _02693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07036_ cpu.uart.receive_div_counter\[7\] _02631_ _01583_ cpu.uart.receive_div_counter\[3\]
+ _02635_ _02636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_70_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05259__S _00830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_rebuffer13_I _00870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05297_ _00831_ _00965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06023__A1 _00832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08987_ _04189_ _04177_ _04191_ _04192_ _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05621__I1 cpu.multiplier.a\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07938_ _03338_ _00278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07869_ _02489_ _03278_ _03286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09608_ _02318_ _02319_ _02337_ _04739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09539_ _03798_ _04688_ _04691_ _00526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07126__I1 cpu.regs\[13\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_118_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05837__A1 cpu.timer_capture\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08832__I _01952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06352__I _00783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10245_ _00503_ clknet_leaf_65_wb_clk_i cpu.ROM_spi_dat_out\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10176_ _00434_ clknet_leaf_50_wb_clk_i cpu.IO_addr_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06014__A1 net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07514__A1 _02944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05828__A1 cpu.spi.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09019__A1 cpu.PC\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08490__A2 _02508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05220_ _00890_ _00891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_25_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05151_ cpu.PORTA_DDR\[2\] net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XTAP_TAPCELL_ROW_77_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05082_ cpu.regs\[8\]\[4\] cpu.regs\[9\]\[4\] cpu.regs\[10\]\[4\] cpu.regs\[11\]\[4\]
+ _00749_ _00750_ _00775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08910_ _03436_ _03848_ _04117_ _04118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09890_ _00149_ clknet_leaf_110_wb_clk_i cpu.regs\[7\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08841_ _02271_ _00768_ _04051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06005__A1 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08772_ _03969_ _03991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05984_ cpu.pwm_top\[4\] _01505_ _01086_ _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07723_ _01900_ _03162_ _03167_ _03161_ _03168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_109_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04935_ _00600_ _00636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06308__A2 _01963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07654_ _03105_ _03101_ _03106_ _03104_ _00226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_88_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04866_ cpu.ROM_spi_cycle\[0\] _00569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_95_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06605_ _02251_ _02260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07585_ _03055_ _03056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09258__A1 _04374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09324_ _04496_ _04497_ _04498_ _04518_ _04519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_48_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06536_ _01941_ _02171_ _02193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09255_ _04103_ _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_63_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06467_ _02088_ _02094_ _02124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05418_ _00588_ _01050_ _01084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__05295__A2 _00960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08206_ _03553_ _03554_ _00330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09186_ _04243_ _04383_ _04384_ _04246_ _04385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_71_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06398_ _02037_ _02044_ _02055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_16_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05349_ _00595_ _00604_ _01002_ _01006_ _01015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_16_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08137_ cpu.toggle_top\[7\] _03482_ _03484_ _03487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08068_ cpu.orig_PC\[1\] _03428_ _03430_ _03440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_83_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_83_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_101_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_12_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_12_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_12_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07019_ cpu.toggle_top\[14\] _02621_ _02623_ _02625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10030_ _00289_ clknet_leaf_29_wb_clk_i cpu.uart.receive_div_counter\[12\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06900__I _02523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09432__B _04571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09249__A1 _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08562__I _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06483__A1 _01730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06483__B2 _01797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10228_ _00486_ clknet_leaf_56_wb_clk_i cpu.mem_cycle\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_72_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09724__A2 _00985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10159_ _00418_ clknet_leaf_55_wb_clk_i cpu.rom_data_dist vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05161__I _00832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07370_ _02859_ _02865_ _02852_ _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06321_ _01941_ _01975_ _01976_ _01978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_29_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06252_ cpu.mem_cycle\[4\] _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09040_ _03840_ _04244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05203_ _00855_ _00874_ _00875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_5_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06183_ cpu.toggle_top\[15\] _01842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_13_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05029__A2 _00722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05134_ _00804_ _00823_ _00824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09942_ _00201_ clknet_leaf_19_wb_clk_i cpu.spi.data_out_buff\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05065_ _00702_ _00759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07816__I _03213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09873_ _00132_ clknet_leaf_95_wb_clk_i cpu.regs\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08824_ _00665_ _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08755_ cpu.last_addr\[3\] _03967_ _03978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05336__I _01001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05967_ _01628_ _01377_ _01381_ _01629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07706_ cpu.uart.counter\[3\] cpu.uart.counter\[2\] _03155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08686_ _03909_ _00748_ _03923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__04960__A1 cpu.uart.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07551__I _03010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04918_ _00619_ _00620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05898_ _01099_ _01560_ _01561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07637_ _03093_ _03094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07568_ cpu.spi.data_out_buff\[6\] _03011_ _03041_ _03042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05060__S1 _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09307_ _03990_ cpu.ROM_addr_buff\[7\] _04487_ _04502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_63_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06519_ _02173_ _02176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_90_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07499_ _02979_ _02981_ _02982_ _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09238_ _03469_ _04434_ _04435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_8_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09169_ _03461_ _03849_ _04342_ _04368_ _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_50_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output71_I net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07717__A1 _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10013_ _00272_ clknet_leaf_35_wb_clk_i cpu.uart.receive_buff\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08557__I _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07461__I _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09642__A1 _04520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08445__A2 _03621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08292__I _03602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06870_ cpu.timer\[4\] _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05821_ _01482_ _01483_ _01484_ _01485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07184__A2 _02729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06931__A2 _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04995__I _00693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08540_ _03801_ _03793_ _03803_ _00415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05752_ cpu.toggle_top\[1\] _01417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08133__A1 cpu.toggle_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05683_ _01313_ _01348_ _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08471_ cpu.timer_capture\[10\] _03746_ _03727_ _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07422_ cpu.spi.data_in_buff\[1\] _02907_ _02913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07353_ _02807_ _02840_ _02849_ _00182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07284_ _02756_ cpu.regs\[6\]\[6\] _02796_ _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06304_ _00746_ _01961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_33_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06235_ _01892_ _01893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09023_ cpu.orig_PC\[4\] _03854_ _04228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06998__A2 _02609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08930__I _04101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06166_ _01824_ _01189_ _01204_ _01825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06097_ _01755_ _01756_ _01757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05117_ _00790_ _00807_ _00808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05048_ _00742_ net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_09925_ _00184_ clknet_leaf_83_wb_clk_i cpu.regs\[2\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09856_ _00115_ clknet_leaf_114_wb_clk_i cpu.regs\[11\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08807_ cpu.orig_flags\[3\] _04017_ _04014_ _04018_ _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09787_ _00050_ clknet_leaf_7_wb_clk_i cpu.timer_capture\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06999_ _02610_ _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08738_ cpu.mem_cycle\[1\] _01914_ _03964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_68_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08124__A1 cpu.toggle_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08377__I _03608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08669_ _03908_ _03909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08675__A2 _00649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09624__B2 _04752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09001__I _04007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06610__A1 _02186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06020_ cpu.regs\[4\]\[6\] cpu.regs\[5\]\[6\] cpu.regs\[6\]\[6\] cpu.regs\[7\]\[6\]
+ _00968_ _00969_ _01681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_42_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05652__A2 _01116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07971_ _03327_ _03364_ _00285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06922_ _02538_ _02533_ _02539_ _02531_ _00061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09710_ _02821_ cpu.regs\[9\]\[6\] _04819_ _04829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09581__I _04710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09641_ _02328_ _04764_ _04766_ _04768_ _04769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_93_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06853_ _02483_ _02484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06784_ _02388_ _02415_ _02424_ _00038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09572_ _02378_ _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05804_ _01468_ _01469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08523_ _00986_ _03791_ _03792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05735_ _00589_ _01027_ _01063_ _01400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_77_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08454_ _01076_ _02469_ _03739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_05666_ _01329_ _01331_ _01332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07405_ _02882_ _02222_ _02207_ _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05597_ _01110_ _01034_ _01263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08385_ _02490_ _03667_ _03682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07336_ _02838_ _02840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07093__A1 _01113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09006_ cpu.PC\[4\] _04073_ _04211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07267_ _02684_ _02777_ _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06218_ cpu.spi.divisor\[7\] _01876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08660__I _00882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07198_ _02753_ cpu.regs\[10\]\[4\] _02745_ _02754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06149_ _01341_ _01808_ _01456_ _01435_ _01809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_41_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09908_ _00167_ clknet_leaf_86_wb_clk_i cpu.regs\[4\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08896__A2 _04103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09839_ _00098_ clknet_leaf_107_wb_clk_i cpu.regs\[13\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_24_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05254__S1 _00837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09440__B _04603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08835__I _04042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08820__A2 _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08570__I _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06831__A1 _02463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05634__A2 _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05190__S0 _00858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_114_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_63_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08336__A1 cpu.timer_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09334__C _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05520_ _01185_ _01186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_87_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05451_ _00600_ _00609_ _00611_ _01004_ _01117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__07311__A2 _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08170_ cpu.toggle_ctr\[3\] _03519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05382_ cpu.IO_addr_buff\[2\] _01048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_07121_ _02697_ _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07052_ cpu.uart.receive_div_counter\[14\] _02652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__06822__A1 cpu.uart.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_93_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06003_ _01660_ _01560_ _01663_ _01665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07954_ cpu.uart.receive_div_counter\[5\] _03351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06905_ _02446_ _02527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07885_ cpu.uart.data_buff\[7\] _03260_ _03298_ _03299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09624_ net76 _04735_ _04737_ _04752_ _04753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06836_ _02467_ _02442_ _02468_ _00046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06767_ _01918_ _02324_ _02410_ _02411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xclkbuf_leaf_37_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_37_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09555_ _03823_ _04696_ _04701_ _00532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06698_ _02295_ _02351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09260__B _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05718_ cpu.uart.divisor\[9\] _01382_ _01383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08506_ cpu.spi.divisor\[2\] _03778_ _03781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_108_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09486_ _04647_ cpu.pwm_counter\[0\] _03589_ _04651_ _04652_ _04653_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_92_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05649_ _01314_ _01315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08437_ cpu.timer\[13\] _03724_ _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08368_ _02978_ _02977_ _02980_ _03667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_33_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08802__A2 _04008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07319_ _02783_ _02826_ _02829_ _00168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08299_ _02463_ _03613_ _03617_ _00360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_34_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05172__S0 _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10261_ _00519_ clknet_leaf_44_wb_clk_i net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__08566__A1 _02640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10192_ _00450_ clknet_leaf_70_wb_clk_i cpu.ROM_addr_buff\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_6_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09294__A2 cpu.last_addr\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput14 io_in[21] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput25 rst_n net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_25_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06813__I _00933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04951_ _00650_ _00651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08676__S _03813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07670_ cpu.uart.div_counter\[15\] _03119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_04882_ cpu.IO_addr_buff\[1\] _00585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07532__A2 _03007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06621_ _02262_ _02275_ _02276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09340_ _04531_ _02410_ _04532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06552_ cpu.PC\[9\] _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08475__I _03607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09271_ _04183_ _04458_ _04366_ _04467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05503_ cpu.br_rel_dest\[0\] _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_75_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08222_ _03563_ _03565_ _00335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_23_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06483_ _01730_ _02018_ _02066_ _01797_ _02140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05434_ _00988_ _01092_ _01097_ _01099_ _01100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_7_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05365_ _01028_ _01030_ _01031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_55_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08153_ _03499_ _01723_ _02620_ _03489_ _03501_ _03502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_7_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08084_ _02214_ _03449_ _03451_ _00311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07104_ _01114_ _02684_ _02692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07035_ _02632_ cpu.uart.receive_div_counter\[13\] cpu.uart.receive_div_counter\[6\]
+ _02633_ _02634_ _02635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_05296_ _00962_ _00963_ _00964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08548__A1 _00674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08986_ _04152_ _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07937_ _02677_ _03337_ _03338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input33_I sram_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05082__I0 cpu.regs\[8\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05621__I2 cpu.regs\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07523__A2 cpu.spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07868_ _03273_ _03284_ _03285_ _00261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05074__I cpu.multiplier.a\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09607_ _01912_ _02317_ _02318_ _02319_ _04738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__05534__A1 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07799_ _03115_ _03195_ _03182_ _03228_ _03229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06819_ _00619_ _02455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09538_ net55 _04689_ _04690_ _04691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05802__I _01466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09469_ _04558_ _04638_ _00509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_100_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08787__A1 cpu.ROM_addr_buff\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05249__I _00918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10244_ _00502_ clknet_leaf_65_wb_clk_i cpu.ROM_spi_dat_out\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10175_ _00433_ clknet_leaf_50_wb_clk_i cpu.IO_addr_buff\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07464__I cpu.timer_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06808__I _00905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08295__I _03608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09267__A2 _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05128__I1 _00815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05150_ cpu.PORTA_DDR\[1\] net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05159__I _00830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05081_ _00772_ _00773_ _00759_ _00774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08840_ _01267_ _04049_ _04050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06005__A2 _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08771_ cpu.last_addr\[7\] _03990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_109_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05983_ _01505_ _01644_ _01645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07722_ _01900_ _03165_ _03167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_04934_ cpu.uart.busy cpu.spi.busy _00635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07653_ cpu.uart.receive_buff\[4\] _03102_ _03106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_04865_ cpu.ROM_spi_cycle\[1\] _00568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_88_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06308__A3 _00916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06604_ _01935_ _02259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09323_ _04500_ _04501_ _04502_ _04517_ _04518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_07584_ _00692_ _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_87_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06535_ _02105_ _02191_ _02192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09254_ _04137_ _04437_ _04450_ _04162_ _04451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_62_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06466_ _02088_ _02094_ _02123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09185_ cpu.orig_PC\[10\] _03863_ _04384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05417_ _01026_ _01083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08205_ _03472_ _03528_ _03554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06397_ _02037_ _02044_ _02054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08136_ _02463_ _03481_ _03486_ _00328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_99_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05348_ cpu.IO_addr_buff\[1\] _00586_ _01013_ _01014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08067_ _03438_ _03439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05279_ _00947_ _00948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07018_ _02460_ _02611_ _02624_ _00072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08941__A1 _04138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08969_ _04169_ _04175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_52_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_52_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_86_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09004__I _02929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10227_ _00485_ clknet_leaf_63_wb_clk_i cpu.mem_cycle\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05994__A1 _00958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08932__A1 cpu.PC\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10158_ _00417_ clknet_leaf_19_wb_clk_i cpu.timer_div\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10089_ _00348_ clknet_leaf_102_wb_clk_i cpu.pwm_counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09342__C _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06171__A1 cpu.spi.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05442__I _01107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08999__A1 _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06320_ _01975_ _01976_ _01941_ _01977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_45_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06251_ cpu.mem_cycle\[5\] _01908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05202_ _00856_ _00873_ _00874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09412__A2 _04592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06182_ cpu.toggle_top\[7\] _01254_ _01260_ _01841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05133_ cpu.regs\[12\]\[7\] cpu.regs\[13\]\[7\] cpu.regs\[14\]\[7\] cpu.regs\[15\]\[7\]
+ _00816_ _00817_ _00823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09941_ _00200_ clknet_leaf_17_wb_clk_i cpu.spi.data_out_buff\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05064_ _00757_ _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09176__A1 _00715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05037__I0 cpu.regs\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09872_ _00131_ clknet_leaf_97_wb_clk_i cpu.regs\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08823_ _01542_ _01566_ _04028_ _04032_ _04033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_29_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08754_ _03972_ _03975_ _03977_ _00455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05966_ cpu.uart.divisor\[4\] _01628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07705_ cpu.uart.counter\[0\] cpu.uart.counter\[1\] _03154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_04917_ _00618_ _00619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08685_ _03922_ _00441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__04960__A2 cpu.spi.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05897_ _01555_ _01559_ _01560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08151__A2 cpu.toggle_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07636_ _03092_ _03093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07567_ _03025_ _03041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09306_ cpu.last_addr\[8\] cpu.ROM_addr_buff\[8\] _04488_ _04501_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__09100__A1 _03433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06518_ _02174_ _02175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_90_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09237_ _02206_ _04408_ _04434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07498_ cpu.timer_top\[3\] _02975_ _02980_ cpu.timer_top\[2\] _02982_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_35_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06449_ _02105_ _00883_ _02106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09168_ _03848_ _04357_ _04368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09099_ _03453_ _04240_ _04301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08119_ cpu.toggle_top\[0\] _03475_ _03467_ _03476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output64_I net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07717__A2 _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10012_ _00271_ clknet_leaf_35_wb_clk_i cpu.uart.receive_buff\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_106_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06153__A1 net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05262__I _00931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06821__I _02456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05820_ _01380_ _01484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_19_Left_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05751_ _01171_ _01415_ _01416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_85_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05682_ _01315_ net90 _01347_ _01348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08470_ _02959_ _03742_ _03752_ _03753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07421_ cpu.spi.dout\[1\] _02911_ _02912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07352_ cpu.regs\[3\]\[7\] _02843_ _02849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08483__I _03739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06303_ _01949_ _01953_ _01959_ _01960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_72_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07283_ _02791_ _02798_ _02805_ _00156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Left_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06234_ cpu.spi.counter\[0\] _01891_ _01892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09022_ _00662_ _04226_ _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06165_ net5 _01824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_96_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_3_0_wb_clk_i clknet_0_wb_clk_i clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_05116_ cpu.regs\[12\]\[6\] cpu.regs\[13\]\[6\] cpu.regs\[14\]\[6\] cpu.regs\[15\]\[6\]
+ _00799_ _00800_ _00807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_40_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06096_ _01294_ _01292_ _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05047_ _00741_ _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09924_ _00183_ clknet_leaf_83_wb_clk_i cpu.regs\[2\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09855_ _00114_ clknet_leaf_115_wb_clk_i cpu.regs\[11\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08806_ _00933_ _04017_ _04018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_37_Left_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06998_ _01258_ _02609_ _02610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_clkbuf_leaf_14_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09786_ _00049_ clknet_leaf_8_wb_clk_i cpu.timer_capture\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08737_ cpu.last_addr\[0\] _03963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05949_ _01573_ _01170_ _01611_ _01306_ _01612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_95_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08668_ _00648_ _03908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_68_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06135__A1 _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07619_ cpu.spi.data_in_buff\[1\] _01894_ _03078_ cpu.spi.data_in_buff\[2\] _03082_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_49_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08599_ _03850_ _03851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_52_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Left_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05949__A1 _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_53_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_55_Left_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06374__B2 _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_101_Right_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08115__A2 _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09620__C _03993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_64_Left_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06429__A2 _01757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_92_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07970_ _02650_ _03309_ _03342_ _03363_ _03364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_73_Left_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06921_ cpu.timer_top\[6\] _02534_ _02539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09551__A1 _03815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09640_ _00578_ _04767_ _04541_ _04768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06852_ _00626_ _02483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_109_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_109_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06783_ _02423_ _02413_ _00685_ _02424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09571_ _04710_ _04712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05803_ _01467_ _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_89_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06117__A1 cpu.spi.divisor\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05734_ cpu.spi.dout\[1\] _01177_ _01398_ _01399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08522_ _03789_ _03791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08453_ _03738_ _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07865__A1 _00906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05665_ _00882_ _01330_ _01331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07404_ _02895_ _02174_ _02896_ _02897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_85_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05596_ cpu.toggle_top\[8\] _01260_ _01261_ _01262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05630__I _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08384_ _03680_ _03681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07617__A1 _03043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07335_ _02838_ _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07266_ _02742_ _02781_ _02794_ _00150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07093__A2 _02684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06217_ cpu.spi.div_counter\[4\] _01875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09005_ _04174_ _04209_ _04210_ _00473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_61_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07197_ _01677_ _02753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06148_ _01799_ _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_111_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06079_ _00796_ _01740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09907_ _00166_ clknet_leaf_88_wb_clk_i cpu.regs\[5\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05077__I _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09542__A1 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09838_ _00097_ clknet_leaf_101_wb_clk_i cpu.regs\[13\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09769_ _00032_ clknet_leaf_81_wb_clk_i cpu.br_rel_dest\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_1_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05190__S1 _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_7_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_7_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_9_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09533__A1 net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06320__B _01941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05450_ cpu.br_rel_dest\[0\] _01116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__06546__I _01938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05381_ _01046_ _01047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_28_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07120_ _01469_ _02699_ _02702_ _00096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_112_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07051_ cpu.uart.divisor\[15\] _02651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XPHY_EDGE_ROW_81_Left_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06002_ _01660_ _01560_ _01663_ _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_07953_ _03349_ _03350_ _00281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07884_ _02508_ _03236_ _03298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06904_ _02525_ _02520_ _02526_ _02524_ _00056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09623_ _04750_ _04751_ _04742_ _04752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06835_ cpu.uart.divisor\[7\] _02435_ _02457_ _02468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06766_ _02338_ _01916_ _02410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09554_ cpu.PORTB_DDR\[2\] _04697_ _04698_ _04701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06697_ net54 _02349_ _02350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05717_ _01381_ _01382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08505_ _02525_ _03777_ _03780_ _00403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09485_ cpu.pwm_top\[6\] cpu.pwm_counter\[6\] _04652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_108_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05648_ _00910_ _01098_ _01314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06510__A1 _01963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08436_ _02965_ _03719_ _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08367_ _03666_ _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05579_ _01242_ _01244_ _01245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07318_ cpu.regs\[4\]\[1\] _02827_ _02829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08298_ cpu.pwm_top\[6\] _03603_ _03615_ _03617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07249_ cpu.regs\[7\]\[1\] _02781_ _02784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10260_ _00518_ clknet_leaf_42_wb_clk_i net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05172__S1 _00839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10191_ _00449_ clknet_leaf_70_wb_clk_i cpu.ROM_addr_buff\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_6_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09515__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08869__A3 _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput15 io_in[23] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput26 sram_out[0] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07925__I _03213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06568__A1 _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09506__A1 _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04950_ _00637_ _00650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_74_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04881_ net25 _00583_ _00584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06620_ _02264_ _02274_ _02275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06551_ cpu.PC\[10\] _02208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_114_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09270_ cpu.PC\[13\] _00912_ _04465_ _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_47_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06482_ _01961_ _01758_ _01955_ _02138_ _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_05502_ _01167_ _01168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05433_ _01098_ _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08221_ cpu.toggle_ctr\[5\] _03564_ _03565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_23_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05364_ _01029_ _01030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08152_ cpu.toggle_ctr\[10\] _01512_ _03500_ _03501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08083_ cpu.orig_PC\[5\] _03443_ _03447_ _03451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05295_ _00951_ _00960_ _00963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07103_ _01616_ _02686_ _02691_ _00090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07034_ cpu.uart.divisor\[9\] _02629_ cpu.uart.receive_div_counter\[5\] _01695_ _02634_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_70_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08985_ _04173_ _04190_ _04191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07936_ _02639_ _03334_ _03336_ _03337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input26_I sram_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07867_ cpu.uart.data_buff\[4\] _03276_ _03041_ _03285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09606_ _04736_ _04734_ _04737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07798_ _03115_ _03227_ _03228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06818_ _02453_ _02454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08720__A2 cpu.regs\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09537_ _04674_ _04690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06749_ _02395_ _02396_ _02397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_78_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09468_ _04631_ _04637_ _04638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_100_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08484__A1 cpu.timer_capture\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09399_ _04546_ _04579_ _04580_ _04581_ _04582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_93_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08419_ _02960_ cpu.timer\[8\] _03698_ _03710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_74_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output94_I net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06798__A1 cpu.uart.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10243_ _00501_ clknet_leaf_65_wb_clk_i cpu.ROM_spi_dat_out\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10174_ _00432_ clknet_leaf_50_wb_clk_i cpu.IO_addr_buff\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05128__I2 cpu.regs\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06824__I _00981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05080_ cpu.regs\[4\]\[4\] cpu.regs\[5\]\[4\] cpu.regs\[6\]\[4\] cpu.regs\[7\]\[4\]
+ _00749_ _00750_ _00773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_110_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07655__I cpu.uart.dout\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08770_ _03984_ _03987_ _03989_ _00459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05982_ cpu.timer_top\[12\] _01598_ _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07721_ _03160_ _03164_ _03166_ _00232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_109_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04933_ _00631_ _00633_ _00634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07652_ cpu.uart.dout\[4\] _03105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_04864_ cpu.ROM_spi_cycle\[4\] _00567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_88_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07583_ cpu.spi.div_counter\[2\] _03045_ _03053_ _03002_ _03054_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06603_ _01752_ _01936_ _02235_ _02258_ _00023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09322_ _03936_ _04504_ _04514_ _04516_ _04517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_87_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06534_ _01732_ _02131_ _02040_ _01798_ _02191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09253_ _04439_ _04449_ _04450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06465_ _02112_ _02118_ _02121_ _02122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_90_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09184_ _04382_ _04383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05416_ _01061_ _01063_ _01067_ _01081_ _01082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_08204_ _03552_ _03553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06396_ _02030_ _02051_ _02052_ _02053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05347_ _00591_ cpu.IO_addr_buff\[2\] _01013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_08135_ cpu.toggle_top\[6\] _03482_ _03484_ _03486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_99_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08066_ _03437_ _03438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05278_ _00946_ _00947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07017_ _01723_ _02621_ _02623_ _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08968_ _04173_ _04073_ _04174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06952__A1 _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07919_ cpu.uart.receive_buff\[6\] _03321_ _03315_ cpu.uart.receive_buff\[5\] _03324_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08899_ _00910_ _04080_ _04107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_92_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_92_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06704__B2 cpu.ROM_addr_buff\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05063__S0 _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_21_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_21_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_39_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05443__A1 _01108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09709__A1 _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09185__A2 _03863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10226_ _00484_ clknet_leaf_63_wb_clk_i cpu.mem_cycle\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08393__B1 _03681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10157_ _00416_ clknet_leaf_19_wb_clk_i cpu.timer_div\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10088_ _00347_ clknet_leaf_104_wb_clk_i cpu.pwm_counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08696__A1 _02214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06250_ cpu.rom_data_dist _01907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_5_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05201_ _00872_ _00873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_108_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06181_ cpu.pwm_top\[7\] _01249_ _01839_ _01171_ _01840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08620__B2 _03870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05132_ _00821_ _00822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_110_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09940_ _00199_ clknet_leaf_17_wb_clk_i cpu.spi.data_out_buff\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05063_ cpu.regs\[8\]\[3\] cpu.regs\[9\]\[3\] cpu.regs\[10\]\[3\] cpu.regs\[11\]\[3\]
+ _00752_ _00753_ _00757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_115_Right_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05037__I1 _00728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09871_ _00130_ clknet_leaf_94_wb_clk_i cpu.regs\[0\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08822_ _01862_ _04024_ _04029_ _04031_ _04032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_08753_ _03920_ _03976_ _03977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05965_ net10 _01626_ _01053_ _01627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_04916_ net25 _00618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07704_ cpu.uart.data_buff\[0\] _03152_ _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08684_ _03919_ _03920_ _03921_ _03922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08687__A1 _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05896_ _00763_ _01558_ _01559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07635_ _02679_ _02678_ _03092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07566_ cpu.spi.data_out_buff\[7\] _03008_ _03039_ _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09305_ cpu.last_addr\[9\] cpu.ROM_addr_buff\[9\] _04499_ _04500_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__06892__C _02506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06517_ _02173_ _02157_ _02174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_106_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09236_ _02204_ _02206_ _04408_ _04433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_61_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07497_ cpu.timer_top\[1\] _02977_ _02980_ cpu.timer_top\[2\] _02981_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_106_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06448_ _00813_ _02105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09167_ _04340_ _04357_ _04365_ _04366_ _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06379_ _02033_ _02034_ _02035_ _02036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09098_ _04101_ _04300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08118_ _03473_ _03475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_43_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08049_ _01427_ _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10011_ _00270_ clknet_leaf_35_wb_clk_i cpu.uart.receive_buff\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output57_I net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05900__A2 _00931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_82_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07169__A1 _02717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10209_ _00467_ clknet_leaf_58_wb_clk_i cpu.TIE vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06916__A1 _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09353__C _03398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05750_ cpu.pwm_top\[1\] _01252_ _01415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05027__S0 _00703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06144__A2 _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05681_ _01316_ _01322_ _01323_ _01346_ _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_07420_ _02910_ _02911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07351_ _02848_ _00181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_116_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06302_ _01940_ _01958_ _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08841__A1 _02271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07282_ cpu.regs\[6\]\[5\] _02801_ _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06233_ _01888_ _01890_ _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09021_ _02416_ _04188_ _04225_ _04194_ _04226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_72_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05655__A1 _00711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06164_ _01055_ _01821_ _01822_ _01823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_13_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05115_ _00805_ _00806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06095_ _01288_ _01290_ _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05046_ _00713_ _00734_ _00740_ _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09923_ _00182_ clknet_leaf_94_wb_clk_i cpu.regs\[3\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_4_12_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09854_ _00113_ clknet_leaf_115_wb_clk_i cpu.regs\[11\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08805_ _04012_ _04017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06907__A1 _02527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06997_ _01093_ _00669_ _02609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09785_ _00048_ clknet_leaf_6_wb_clk_i cpu.timer_capture\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08736_ _03962_ _00452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05948_ _01170_ _01610_ _01611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08667_ _02388_ _03900_ _03907_ _00438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05879_ _01329_ _01331_ _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07332__A1 _02807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07618_ _02364_ _03081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_71_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08598_ _01159_ _03849_ _03850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_52_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09085__A1 _02421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07549_ cpu.spi.data_out_buff\[2\] _03016_ _03026_ _03027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_101_Left_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09219_ cpu.PC\[11\] _01099_ _04417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_51_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_80_Right_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08899__A1 _00910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05257__S0 _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_109_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06832__I _01761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05448__I _01113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08759__I _03966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06920_ _02462_ _02538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06988__B _02558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07663__I _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06851_ _02480_ _02473_ _02474_ _02481_ _02482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06782_ _01110_ _02423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09570_ _04710_ _04711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05802_ _01466_ _01467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09303__A2 cpu.ROM_addr_buff\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08521_ _03789_ _03790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05733_ _01397_ _01398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08452_ cpu.timer_capture\[15\] _03714_ _03737_ _03722_ _03738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05664_ _01157_ _01330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__05876__A1 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07403_ _02895_ _02174_ _01925_ _02896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05595_ _01060_ _01261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08383_ _03655_ _03680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08814__A1 _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07334_ _02837_ _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_45_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07265_ cpu.regs\[7\]\[7\] _02786_ _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09004_ _02929_ _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06216_ _01872_ cpu.spi.divisor\[3\] cpu.spi.divisor\[7\] _01873_ _01874_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06742__I _02390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09258__C _04007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07196_ _02722_ _02746_ _02752_ _00122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06147_ _01802_ _01806_ _01807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_13_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06078_ _01736_ _01738_ _01739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06053__A1 cpu.timer_capture\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05800__A1 net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09906_ _00165_ clknet_leaf_91_wb_clk_i cpu.regs\[5\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05029_ _00702_ _00722_ _00724_ _00003_ _00725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__08669__I _03908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09837_ _00096_ clknet_leaf_101_wb_clk_i cpu.regs\[13\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09768_ _00031_ clknet_leaf_81_wb_clk_i cpu.br_rel_dest\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_57_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05093__I _00770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08719_ _03908_ _03949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_68_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09699_ cpu.regs\[9\]\[1\] _04821_ _04823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_1_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09230__A1 _00748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06044__A1 _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09049__A1 _04138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05858__A1 _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05380_ _00594_ _00604_ _01001_ _01005_ _01046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_15_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07050_ cpu.uart.receive_div_counter\[8\] _02650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07658__I cpu.uart.dout\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06001_ _00780_ _01662_ _01663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_2_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07952_ cpu.uart.receive_div_counter\[4\] _03347_ _03234_ _03350_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07883_ _03291_ _03296_ _03297_ _00264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06903_ cpu.timer_top\[1\] _02521_ _02526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09622_ _03936_ _02355_ _02356_ cpu.ROM_addr_buff\[10\] _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06834_ _02466_ _02467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_37_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09553_ _03820_ _04696_ _04700_ _00531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08504_ cpu.spi.divisor\[1\] _03778_ _03780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06765_ _02388_ _02402_ _02409_ _00034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06696_ _02344_ _02346_ _02348_ _02349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05716_ _01380_ _01381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09484_ cpu.pwm_top\[2\] _04651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_93_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05647_ _01312_ _01309_ _01313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__05849__A1 _01512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08435_ _03723_ _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_34_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08366_ cpu.timer_capture\[1\] _03663_ _03665_ _03257_ _03666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_18_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05578_ cpu.timer_top\[0\] _01243_ _01244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07317_ _02776_ _02826_ _02828_ _00167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08297_ _02460_ _03613_ _03616_ _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_46_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_46_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_61_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07248_ _01467_ _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07179_ _01816_ cpu.regs\[11\]\[6\] _02731_ _02741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10190_ _00448_ clknet_leaf_69_wb_clk_i cpu.ROM_addr_buff\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05088__I _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09279__A1 _00784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput16 io_in[26] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_107_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput27 sram_out[1] net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09179__B _04324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07478__I cpu.timer_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05068__A2 _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06568__A2 _02223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05791__A3 _01329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04880_ _00566_ _00582_ _00583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05623__S0 _01285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06557__I cpu.PC\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06550_ _02206_ _02207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_114_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06481_ _01758_ _01956_ _01961_ _02138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05501_ _01166_ _01167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08772__I _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05432_ cpu.base_address\[2\] _01098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09690__A1 _01303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08220_ cpu.toggle_ctr\[4\] _03559_ _03564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_31_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05363_ cpu.IO_addr_buff\[4\] _00593_ _01029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08151_ _03490_ cpu.toggle_top\[11\] _03500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08082_ _02556_ _03449_ _03450_ _00310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_82_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05294_ _00936_ _00950_ _00962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07102_ cpu.regs\[14\]\[3\] _02685_ _02691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07033_ _01771_ _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_113_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08721__B _03950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07756__A1 _03088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08548__A3 _01041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08984_ _04149_ _04190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07935_ _02639_ _03328_ _03335_ _03336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05082__I2 cpu.regs\[10\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09605_ _02315_ _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_98_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07866_ cpu.uart.data_buff\[3\] _03282_ _03283_ _03284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input19_I io_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07797_ cpu.uart.div_counter\[11\] _03221_ _03227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06817_ _01694_ _02453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09536_ _04680_ _04689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06748_ _01908_ _01910_ _02325_ _02396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09467_ _03079_ _04636_ _04637_ _00508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06679_ _02331_ _00578_ _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_65_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08418_ _03709_ _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09398_ _04546_ _04577_ _00693_ _04581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_81_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08349_ _00589_ _01013_ _01079_ _02431_ _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_6_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10242_ _00500_ clknet_leaf_65_wb_clk_i cpu.ROM_spi_dat_out\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07747__A1 _02677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10173_ _00431_ clknet_leaf_14_wb_clk_i cpu.IO_addr_buff\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06022__I1 cpu.multiplier.a\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05281__I _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07683__B1 _01583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06840__I _01220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07720_ _01889_ _03165_ _03161_ _03166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_109_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05981_ _01620_ _01243_ _01411_ _01642_ _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_04932_ _00625_ _00632_ _00633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07651_ _03100_ _03101_ _03103_ _03104_ _00225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_88_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04863_ cpu.instr_cycle\[2\] _00566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07582_ cpu.spi.div_counter\[2\] _03048_ _03044_ _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06602_ net12 _01923_ _02237_ _02253_ _02255_ _02257_ _02258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
X_09321_ cpu.last_addr\[5\] cpu.ROM_addr_buff\[5\] _04515_ _04516_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_75_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06533_ _00815_ _00948_ _02190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08716__B _03946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09663__A1 _02419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09252_ _04346_ _04445_ _04448_ _04449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06464_ net128 _02092_ _02120_ _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09183_ _02208_ _04381_ _04382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05415_ _01074_ _01075_ _01080_ _01081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_44_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06395_ _02047_ _02050_ _02052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08203_ _00621_ _03551_ _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05346_ _00993_ _00999_ _01011_ _01012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_71_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08134_ _02460_ _03481_ _03485_ _00327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_99_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06324__S1 _01950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_33_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08065_ _03436_ _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_70_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05277_ _00945_ _00946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07016_ _02456_ _02623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08967_ _02217_ _04173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07918_ _03320_ _03323_ _00273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09282__B _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08898_ _00659_ _04106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07849_ cpu.uart.data_buff\[0\] _03249_ _03269_ _03270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_79_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05063__S1 _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09519_ net66 _04673_ _04675_ _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_61_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_61_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_72_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06925__I _02523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05443__A2 _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10225_ _00483_ clknet_4_15_0_wb_clk_i cpu.PC\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_72_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10156_ _00415_ clknet_leaf_19_wb_clk_i cpu.timer_div\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10087_ _00346_ clknet_leaf_104_wb_clk_i cpu.pwm_counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05682__A2 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05200_ _00871_ _00872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06180_ _01836_ _01837_ _01838_ _01839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_111_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05131_ cpu.regs\[8\]\[7\] cpu.regs\[9\]\[7\] cpu.regs\[10\]\[7\] cpu.regs\[11\]\[7\]
+ _00816_ _00817_ _00821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_05062_ _00735_ _00756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05434__A2 _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09870_ _00129_ clknet_leaf_97_wb_clk_i cpu.regs\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08821_ _01744_ _04030_ _04031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_0_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_117_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05037__I2 _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06934__A2 _01906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08752_ _03969_ _03976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05964_ _01621_ _01188_ _01624_ _01625_ _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08136__A1 _02463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08683_ _03812_ _03921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_04915_ net71 _00617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07703_ _03151_ _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07634_ cpu.uart.dout\[0\] _03091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05895_ _01156_ _01557_ _01558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07565_ _02513_ _03038_ _03039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09304_ cpu.last_addr\[8\] _04488_ _04499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07496_ cpu.timer\[2\] _02980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_8_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06516_ _02160_ _02168_ _02172_ _02173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_09235_ _02205_ _04379_ _04432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06447_ _02081_ _02102_ _02103_ _02104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_8_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09166_ _04147_ _04366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05673__A2 _01333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06378_ _01950_ _00978_ _02034_ _01967_ _02035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_43_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09097_ _04169_ _04299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05329_ _00994_ _00995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08117_ _03473_ _03474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08048_ _01303_ _03423_ _03424_ _00302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05425__A2 _01056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10010_ _00269_ clknet_leaf_35_wb_clk_i cpu.uart.receive_buff\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09999_ _00258_ clknet_leaf_24_wb_clk_i cpu.uart.data_buff\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05029__C _00003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08127__A1 _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_55_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08850__A2 _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06613__A1 _01759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08366__A1 cpu.timer_capture\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10208_ _00466_ clknet_leaf_69_wb_clk_i cpu.last_addr\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10139_ _00398_ clknet_leaf_4_wb_clk_i cpu.timer_capture\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05680_ _01332_ _01334_ _01338_ _01345_ _01346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__05027__S1 _00704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07350_ _02821_ cpu.regs\[3\]\[6\] _02838_ _02848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06301_ _00861_ net125 net117 _00866_ _01957_ _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_09020_ _04189_ _04213_ _04224_ _04192_ _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08841__A2 _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07281_ _02804_ _00155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06232_ cpu.spi.counter\[3\] cpu.spi.counter\[2\] cpu.spi.counter\[4\] _01889_ _01890_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_5_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06163_ net67 _01018_ _01822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05114_ cpu.regs\[8\]\[6\] cpu.regs\[9\]\[6\] cpu.regs\[10\]\[6\] cpu.regs\[11\]\[6\]
+ _00799_ _00800_ _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06094_ _01354_ _01753_ _01754_ _00018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09922_ _00181_ clknet_leaf_90_wb_clk_i cpu.regs\[3\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05045_ _00735_ _00737_ _00739_ _00713_ _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_40_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06080__A2 _00979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09853_ _00112_ clknet_leaf_113_wb_clk_i cpu.regs\[11\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08804_ _00687_ _04015_ _04016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09784_ _00047_ clknet_leaf_8_wb_clk_i cpu.timer_capture\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08735_ _03961_ cpu.ROM_addr_buff\[13\] _03952_ _03962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06996_ cpu.toggle_top\[8\] _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_05947_ _00687_ _01298_ _01608_ _01609_ _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__05591__A1 cpu.toggle_top\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08666_ _00911_ _03901_ _03904_ _03907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05878_ _01541_ _01540_ _01542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07617_ _03043_ _03080_ _00215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08597_ _03848_ _03849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_105_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07548_ _03025_ _03026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_24_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07479_ _02962_ cpu.timer\[11\] _02959_ _02958_ _02963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_106_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08690__I _03908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09218_ _01327_ _04192_ _04415_ _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09149_ _04166_ _04328_ _04350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08348__A1 _02540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08899__A2 _04080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05257__S1 _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07020__A1 _02463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05193__S0 _00858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08105__I _03456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06850_ cpu.timer\[1\] _02475_ _02481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07011__A1 _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05801_ _01429_ _01433_ _01464_ _01465_ _01466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_117_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06781_ _02385_ _02415_ _02422_ _00037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_89_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08520_ _01395_ _02469_ _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05732_ _01396_ _01397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05663_ _01328_ _01329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_26_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08451_ _02998_ _03736_ _03662_ _03737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07402_ _02885_ _02887_ _02895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_73_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05594_ _01259_ _01260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08382_ _03668_ _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07333_ _01165_ _02543_ _02837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_118_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_118_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07264_ _02793_ _00149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06215_ cpu.spi.div_counter\[7\] _01873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09003_ _04175_ _04203_ _04208_ _04209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07195_ cpu.regs\[10\]\[3\] _02750_ _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06146_ _01736_ _01738_ _01805_ _01806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__06589__B1 _02040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06077_ _01737_ _01665_ _01738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09905_ _00164_ clknet_leaf_88_wb_clk_i cpu.regs\[5\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05028_ _00707_ _00723_ _00724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09836_ _00095_ clknet_leaf_101_wb_clk_i cpu.regs\[13\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09767_ _00030_ clknet_leaf_54_wb_clk_i cpu.instr_buff\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_57_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06979_ _02584_ _02592_ _02593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08718_ _03948_ _00448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09698_ _01352_ _04820_ _04822_ _00554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08649_ cpu.orig_IO_addr_buff\[7\] _03842_ _03845_ _01297_ _03894_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08502__A1 cpu.spi.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06816__A1 _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05175__S0 _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08569__A1 _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07004__I _02610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06807__A1 _02440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08544__B _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06000_ _00880_ _01661_ _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_93_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07951_ cpu.uart.receive_div_counter\[4\] _03345_ _03346_ _03348_ _03349_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06902_ _02443_ _02525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05794__A1 _00726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05408__B _01073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07882_ cpu.uart.data_buff\[7\] _03288_ _03289_ _03297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09621_ _03920_ _04738_ _04739_ _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07535__A2 _03007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06833_ _02465_ _02466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09552_ cpu.PORTB_DDR\[1\] _04697_ _04698_ _04700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06764_ _01573_ _02400_ _02406_ _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05715_ _01008_ _01210_ _01380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_77_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08503_ _02518_ _03777_ _03779_ _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06695_ cpu.spi_clkdiv _02347_ _02348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09483_ _04645_ _04646_ _04648_ _04649_ _04650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_TAPCELL_ROW_102_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05646_ _01139_ _01312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05849__A2 _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08434_ cpu.timer_capture\[12\] _03714_ _03721_ _03722_ _03723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_34_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05577_ _01235_ _01243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08365_ _02998_ _03664_ _03662_ _03665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08799__A1 _01041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06753__I _02400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07316_ cpu.regs\[4\]\[0\] _02827_ _02828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08296_ cpu.pwm_top\[5\] _03603_ _03615_ _03616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07247_ _02776_ _02780_ _02782_ _00143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07178_ _02725_ _02733_ _02740_ _00116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06129_ cpu.toggle_top\[14\] _01172_ _01137_ _01789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06026__A2 _00843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08971__A1 _04173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_86_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_86_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_15_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_15_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_6_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09819_ _00078_ clknet_leaf_80_wb_clk_i _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_69_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08348__C _03648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput17 io_in[28] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput28 sram_out[2] net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_64_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05528__A1 _01190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08539__B _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05623__S1 _01286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05500_ _01114_ _01165_ _01166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06480_ _02129_ _02136_ _02137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_05431_ _01096_ _01097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05700__A1 cpu.PORTB_DDR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08150_ cpu.toggle_ctr\[13\] _03499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_23_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05362_ _00992_ _01013_ _01028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_7_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07101_ _01552_ _02686_ _02690_ _00089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08081_ cpu.orig_PC\[4\] _03443_ _03447_ _03450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05293_ _00961_ net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07032_ cpu.uart.divisor\[13\] _02632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA_clkbuf_leaf_23_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08983_ _04150_ _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07934_ _03329_ _03335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05082__I3 cpu.regs\[11\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07865_ _00906_ _03278_ _03283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_39_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09604_ _04734_ _04735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07796_ _03214_ _03226_ _00248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06816_ _02451_ _02436_ _02452_ _00042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09535_ _04680_ _04688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06747_ _01913_ _02316_ _02395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_78_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06678_ net130 _02331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09466_ _04632_ _00568_ _04627_ _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA_clkbuf_leaf_62_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07692__A1 _02640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09681__A2 _00958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05629_ _01288_ _01290_ _01292_ _01294_ _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_08417_ cpu.timer_capture\[9\] _03678_ _03708_ _03690_ _03709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09397_ _04547_ _04572_ _04569_ _04580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_108_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08348_ _02540_ _03643_ _03649_ _03648_ _00377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_104_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08279_ _03603_ _03604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10241_ _00499_ clknet_leaf_62_wb_clk_i cpu.ROM_spi_dat_out\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10172_ _00430_ clknet_leaf_14_wb_clk_i cpu.IO_addr_buff\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05758__A1 _01335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06022__I2 cpu.regs\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05930__A1 cpu.spi.dout\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_66_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07435__A1 _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06238__A2 _01895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_107_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05980_ cpu.timer_capture\[12\] _01233_ _01641_ _01236_ _01642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_04931_ cpu.IE cpu.needs_interrupt _00632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07650_ _03055_ _03104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_88_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07581_ _03048_ _03044_ _03052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05921__A1 _01583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06601_ _02256_ _02257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09320_ _03980_ _04486_ _04515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06532_ _02186_ _01758_ _02014_ _02188_ _02189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_09251_ _00936_ _04256_ _04447_ _04262_ _04448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06463_ _02119_ _00872_ _02093_ _02120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08202_ _03472_ _03550_ _03551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_28_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09182_ _02221_ _04212_ _04381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05414_ _01078_ _01079_ _01080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06394_ _02047_ _02050_ _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05345_ _01010_ _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_50_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08133_ cpu.toggle_top\[5\] _03482_ _03484_ _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_99_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08064_ cpu.PC\[1\] _03436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_113_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05988__A1 cpu.toggle_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05276_ _00938_ _00940_ _00942_ _00944_ _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_07015_ _02454_ _02615_ _02622_ _00071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_101_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09718__A3 _04834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input31_I sram_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08958__I _04091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08966_ _03885_ _04172_ _00472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07917_ cpu.uart.receive_buff\[5\] _03321_ _03315_ cpu.uart.receive_buff\[4\] _03323_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08897_ _04103_ _04099_ _04104_ _04105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07848_ _03265_ _03269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05912__A1 net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09518_ _03801_ _04672_ _04677_ _00519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07779_ _02363_ _03213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09449_ _04609_ _04622_ _04623_ _00504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_66_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07417__A1 cpu.spi.dout\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_30_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_30_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05979__A1 _01638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10224_ _00482_ clknet_leaf_74_wb_clk_i cpu.PC\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10155_ _00414_ clknet_leaf_9_wb_clk_i cpu.timer_div\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09590__A1 cpu.PORTA_DDR\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10086_ _00345_ clknet_leaf_117_wb_clk_i cpu.toggle_ctr\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07012__I cpu.toggle_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05130_ _00818_ _00819_ _00804_ _00820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_111_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05061_ _00751_ _00754_ _00735_ _00755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_111_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08820_ _01659_ _01670_ _04030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05037__I3 cpu.regs\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08751_ cpu.last_addr\[2\] _03967_ _03975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07615__C _03079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05963_ net63 _01017_ _01188_ _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08682_ cpu.ROM_addr_buff\[2\] _03920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04914_ _00616_ _00012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07702_ _03150_ _03151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05894_ _00956_ _01556_ _01557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07633_ _03088_ _03090_ _00221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07564_ _03006_ _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09303_ cpu.last_addr\[11\] cpu.ROM_addr_buff\[11\] _04490_ _04498_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_07495_ cpu.timer_top\[1\] _02977_ _02978_ cpu.timer_top\[0\] _02979_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06515_ _00747_ _02171_ _02172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08018__I _03400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09234_ _04407_ _04430_ _04431_ _00481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_63_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06446_ _02098_ _02101_ _02103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09165_ _04362_ _04363_ _04364_ _04365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04881__A1 net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08116_ _01085_ _02433_ _03473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06377_ _01946_ _01797_ _02034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09096_ _02596_ _04273_ _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05328_ cpu.IO_addr_buff\[1\] _00994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07078__B _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08047_ cpu.orig_flags\[0\] _03418_ _03421_ _03424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05259_ _00927_ _00928_ _00830_ _00929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_102_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07806__B _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09998_ _00257_ clknet_leaf_25_wb_clk_i cpu.uart.counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06386__A1 _00783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08949_ _00661_ _04148_ _04155_ _04156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07541__B _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08063__A1 _03433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10207_ _00465_ clknet_leaf_69_wb_clk_i cpu.last_addr\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07435__C _00694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10138_ _00397_ clknet_leaf_5_wb_clk_i cpu.timer_capture\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06129__A1 cpu.toggle_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10069_ _00328_ clknet_leaf_3_wb_clk_i cpu.toggle_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_82_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06846__I _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07280_ _02753_ cpu.regs\[6\]\[4\] _02796_ _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06300_ _01955_ _01956_ _01957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_116_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06231_ cpu.spi.counter\[0\] cpu.spi.counter\[1\] _01889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_73_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06162_ _01364_ _01819_ _01820_ _01476_ _01821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06581__I _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05113_ _00756_ _00804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06093_ cpu.regs\[15\]\[5\] _01553_ _01754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05044_ _00735_ _00738_ _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09921_ _00180_ clknet_leaf_94_wb_clk_i cpu.regs\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09852_ _00111_ clknet_leaf_112_wb_clk_i cpu.regs\[11\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08803_ _03403_ _04014_ _04015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09783_ _00046_ clknet_leaf_26_wb_clk_i cpu.uart.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09306__A1 cpu.last_addr\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08734_ _02254_ _03949_ _03960_ _03961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06995_ _02552_ _02606_ _02607_ _00066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05946_ _00905_ _01282_ _01298_ _01609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08665_ _02385_ _03900_ _03906_ _00437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05877_ _00742_ _00904_ _01541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07616_ cpu.spi.data_in_buff\[0\] _01894_ _03078_ cpu.spi.data_in_buff\[1\] _03080_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08596_ _03847_ _03848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_105_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07547_ _02455_ _03025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_24_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07478_ cpu.timer_top\[11\] _02962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_118_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09217_ _04342_ _04414_ _04415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06429_ _01946_ _01757_ _01967_ _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07587__I _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09148_ _04300_ _04329_ _04348_ _04317_ _04349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09079_ _04279_ _04280_ _04281_ _04282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_15_Left_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output62_I net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09545__A1 _03833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06359__A1 cpu.multiplier.a\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05582__A2 _01073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_24_Left_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06531__A1 _02009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09042__I _04106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Left_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05193__S1 _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07446__B _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08121__I _03456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05800_ net27 _01310_ _01311_ _01465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_42_Left_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06780_ _02421_ _02413_ _00685_ _02422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05731_ _01395_ _01009_ _01224_ _01396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_05662_ _01327_ cpu.base_address\[2\] _01328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08450_ cpu.timer\[15\] _03735_ _03736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08381_ _03677_ _03678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07401_ _02854_ _02893_ _02894_ _00185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05593_ _01011_ _01258_ _01259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07332_ _02807_ _02827_ _02836_ _00174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_51_Left_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07263_ _02756_ cpu.regs\[7\]\[6\] _02779_ _02793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06214_ _01871_ _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09002_ _02389_ _04178_ _04205_ _04206_ _04207_ _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_5_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07194_ _02719_ _02746_ _02751_ _00121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06145_ net95 _01735_ _01805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06589__A1 _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06076_ _00780_ _01662_ _01737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_41_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09527__A1 net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09904_ _00163_ clknet_leaf_91_wb_clk_i cpu.regs\[5\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05027_ cpu.regs\[12\]\[1\] cpu.regs\[13\]\[1\] cpu.regs\[14\]\[1\] cpu.regs\[15\]\[1\]
+ _00703_ _00704_ _00723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09835_ _00094_ clknet_leaf_97_wb_clk_i cpu.regs\[14\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09766_ _00029_ clknet_leaf_52_wb_clk_i cpu.instr_buff\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_57_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06761__A1 _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06978_ _02257_ _02586_ _02591_ _02592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08717_ _03947_ cpu.ROM_addr_buff\[9\] _03937_ _03948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_83_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05929_ _01587_ _01590_ _01591_ _01592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09697_ cpu.regs\[9\]\[0\] _04821_ _04822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08648_ _03885_ _03893_ _00433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_1_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08579_ _03804_ _03826_ _03832_ _00425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07069__A2 net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05175__S1 _00839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05627__I0 cpu.regs\[8\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09518__A1 _03801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05252__A1 _00913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07780__I _03213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05555__A2 _01220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04909__I _00611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_2_0_wb_clk_i clknet_0_wb_clk_i clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_86_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06504__A1 _02105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09500__I _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_13_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07950_ cpu.uart.receive_div_counter\[4\] _03347_ _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09509__A1 net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06901_ _02518_ _02520_ _02522_ _02524_ _00055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05794__A2 _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07881_ cpu.uart.data_buff\[6\] _03282_ _03295_ _03296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09620_ _04745_ _04735_ _04749_ _03993_ _00549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06743__A1 _02389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06832_ _01761_ _02465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_37_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09551_ _03815_ _04696_ _04699_ _00530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06763_ _02385_ _02402_ _02408_ _00033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05714_ _01376_ _01378_ _01208_ _01379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08502_ cpu.spi.divisor\[0\] _03778_ _03779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06694_ _00569_ _02294_ _02347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09482_ cpu.pwm_top\[5\] cpu.pwm_counter\[5\] _04649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_102_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08433_ _00627_ _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_77_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_52_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05645_ _01104_ _01311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05849__A3 _01126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08364_ cpu.timer\[1\] _03658_ _03664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_46_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05576_ _01241_ _01242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08248__A1 _02478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07315_ _02825_ _02827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08295_ _03608_ _03615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07246_ cpu.regs\[7\]\[0\] _02781_ _02782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07177_ cpu.regs\[11\]\[5\] _02736_ _02740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09748__A1 _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06128_ cpu.toggle_top\[6\] _01253_ _01259_ _01788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_113_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06059_ cpu.pwm_top\[5\] _01505_ _01418_ _01720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_6_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08184__B1 cpu.toggle_top\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06734__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_91_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09818_ _00077_ clknet_leaf_94_wb_clk_i _00006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xclkbuf_leaf_55_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_55_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09749_ _04837_ _04861_ _04862_ _00565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_68_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput18 io_in[29] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput29 sram_out[3] net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05776__A2 _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08175__B1 cpu.toggle_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06025__I0 cpu.regs\[12\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05084__S0 _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05430_ _00618_ _01093_ _01095_ _01096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_28_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05361_ _01026_ _01027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_31_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07100_ cpu.regs\[14\]\[2\] _02687_ _02690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08080_ _03403_ _03449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08650__A1 _02423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05292_ _00951_ _00960_ _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_3_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07031_ _01818_ _02631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__05464__A1 _01031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08982_ _04116_ _04188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07933_ _03333_ _03331_ _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07864_ _03207_ _03282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_39_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09603_ _01000_ _00580_ _02343_ _04734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__06716__A1 _00579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06815_ cpu.uart.divisor\[3\] _02437_ _02391_ _02452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07795_ cpu.uart.div_counter\[11\] _03178_ _03182_ _03225_ _03226_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_64_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06746_ _02393_ _02394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09534_ _03796_ _04681_ _04687_ _00525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08469__A1 _00906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06677_ _02323_ _02329_ _02330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09465_ _04630_ _04628_ _04632_ _04636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05628_ _01284_ _01293_ _01294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08416_ _02990_ _03679_ _03681_ _03707_ _03684_ _03708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_09396_ _02360_ _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_74_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05559_ _01066_ _01224_ _01225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08347_ cpu.timer_top\[15\] _03644_ _03649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08278_ _03602_ _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_102_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_102_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07229_ _02719_ _02765_ _02770_ _00137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06713__B _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10240_ _00498_ clknet_leaf_61_wb_clk_i cpu.ROM_spi_dat_out\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10171_ _00429_ clknet_leaf_15_wb_clk_i cpu.IO_addr_buff\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05302__S1 _00969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_110_Right_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05066__S0 _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09050__I _04147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_7_Left_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08632__B2 _00950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08935__A2 _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06946__A1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04930_ _00624_ _00631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06849__I _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05057__S0 _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07371__A1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07580_ _03049_ _03051_ _02930_ _00207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06600_ _01926_ _02256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09112__A2 _03854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06531_ _02009_ _02187_ _02188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09250_ _04257_ _04436_ _04446_ _04342_ _04447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xclkbuf_leaf_0_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_0_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_90_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08871__A1 _01303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08201_ _03510_ _03525_ _03535_ _03549_ _03550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_06462_ _02105_ _02119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09181_ _02882_ _04379_ _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05413_ cpu.IO_addr_buff\[4\] _00593_ _01079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_50_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06393_ _02011_ _02048_ _02049_ _02050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05344_ _01009_ _01010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08623__A1 _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08132_ _03456_ _03484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_99_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08063_ _03433_ _03434_ _03435_ _00306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_71_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05275_ _00943_ _00006_ _00944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_71_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05988__A2 _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07014_ _02620_ _02621_ _02616_ _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_24_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08304__I _02944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08926__A2 _03433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08965_ _04131_ _04072_ _04171_ _03836_ _04172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07916_ _03320_ _03322_ _00272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input24_I io_in[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08896_ _04043_ _04103_ _04104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07847_ cpu.uart.data_buff\[1\] _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07362__A1 _02856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07778_ _03088_ _03212_ _00244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09517_ net64 _04673_ _04675_ _04677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_108_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06729_ _02373_ _02376_ _02380_ _00027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09103__A2 _01034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09448_ cpu.ROM_spi_dat_out\[6\] _04594_ _04603_ _04623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09379_ _04565_ _00492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output92_I net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10223_ _00481_ clknet_leaf_74_wb_clk_i cpu.PC\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_70_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_70_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10154_ _00413_ clknet_leaf_20_wb_clk_i cpu.timer_div\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_72_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09045__I _04108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10085_ _00344_ clknet_leaf_117_wb_clk_i cpu.toggle_ctr\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07353__A1 _02807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05903__A2 _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04917__I _00618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08605__A1 _03850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09648__C _03398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06353__B _02009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05060_ cpu.regs\[4\]\[3\] cpu.regs\[5\]\[3\] cpu.regs\[6\]\[3\] cpu.regs\[7\]\[3\]
+ _00752_ _00753_ _00754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06919__A1 _02536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08750_ _03972_ _03973_ _03974_ _00454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05962_ _01364_ _01622_ _01623_ _01198_ _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08681_ _03442_ _03917_ _03918_ _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04913_ _00615_ _00616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07701_ _03124_ _03149_ _03150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05893_ _01325_ _01107_ _01556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07632_ cpu.spi.data_in_buff\[6\] _01893_ _03085_ cpu.spi.data_in_buff\[7\] _03090_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09302_ cpu.last_addr\[10\] cpu.ROM_addr_buff\[10\] _04489_ _04497_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_88_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07563_ _03028_ _03036_ _03037_ _00204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07494_ cpu.timer\[0\] _02978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_48_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06514_ _01968_ _02170_ _02171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09233_ _00693_ _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_61_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06445_ _02101_ _02098_ _02102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_4_15_0_wb_clk_i clknet_0_wb_clk_i clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_90_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09164_ _04362_ _04363_ _04108_ _04364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04881__A2 _00583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08115_ _03472_ _02365_ _00321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06376_ _01967_ _02033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09095_ _04274_ _04297_ _04210_ _00476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05327_ _00989_ _00992_ _00993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__05658__I _00908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08046_ _03401_ _03423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05258_ cpu.regs\[0\]\[3\] cpu.multiplier.a\[3\] cpu.regs\[2\]\[3\] cpu.regs\[3\]\[3\]
+ _00889_ _00926_ _00928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_43_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08969__I _04169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09021__A1 _02416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05830__A1 cpu.spi.dout\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05189_ _00857_ _00860_ _00861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_101_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09997_ _00256_ clknet_leaf_25_wb_clk_i cpu.uart.counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08948_ _01525_ _04116_ _04153_ _04154_ _04155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_98_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08879_ _04078_ _04083_ _04087_ _00657_ _04088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__07822__B _03242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_88_Left_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09088__A1 _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_97_Left_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_74_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10206_ _00464_ clknet_leaf_69_wb_clk_i cpu.last_addr\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06377__A2 _01797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10137_ _00396_ clknet_leaf_5_wb_clk_i cpu.timer_capture\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10068_ _00327_ clknet_leaf_117_wb_clk_i cpu.toggle_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_85_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06230_ _01874_ _01877_ _01881_ _01887_ _01888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_72_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06161_ net47 _01021_ _01820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09251__A1 _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05112_ _00801_ _00802_ _00790_ _00803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06092_ _01752_ _01753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05043_ cpu.regs\[12\]\[2\] cpu.regs\[13\]\[2\] cpu.regs\[14\]\[2\] cpu.regs\[15\]\[2\]
+ _00716_ _00717_ _00738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_09920_ _00179_ clknet_leaf_95_wb_clk_i cpu.regs\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_40_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06811__B _02391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07565__A1 _02513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09851_ _00110_ clknet_leaf_102_wb_clk_i cpu.regs\[12\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08802_ _04007_ _04008_ _04013_ _04014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_09782_ _00045_ clknet_leaf_17_wb_clk_i cpu.uart.divisor\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06994_ _02271_ _02567_ _02607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09306__A2 cpu.ROM_addr_buff\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08733_ _03916_ cpu.regs\[3\]\[5\] _03960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05945_ _01471_ _01606_ _01607_ _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_96_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08664_ _00913_ _03901_ _03904_ _03906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05876_ net92 _00917_ _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07615_ _03076_ _01894_ _03078_ _02906_ _03079_ _00214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08595_ cpu.base_address\[5\] _00935_ _01161_ _03847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__05879__A1 _01329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08029__I _03410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07546_ cpu.spi.data_out_buff\[3\] _03021_ _03023_ _03024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09216_ _04258_ _04409_ _04413_ _04414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07477_ _02958_ _02959_ _02960_ _02955_ _02961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06428_ _02084_ _00782_ _02085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_44_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09147_ _04331_ _04347_ _04348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06359_ cpu.multiplier.a\[5\] _02015_ _02016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09078_ _02213_ _02421_ _04281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06056__A1 _01716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08029_ _03410_ _03411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_116_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07556__A1 _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output55_I net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06047__A1 cpu.spi.divisor\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06631__B _02070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09661__C _03993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09233__I _00693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05730_ _00995_ _01076_ _01395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_clkbuf_leaf_42_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05661_ _01326_ _01327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_58_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08380_ _03650_ _03677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07400_ _00729_ _02869_ _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05592_ _01079_ _01051_ _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_58_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07331_ cpu.regs\[4\]\[7\] _02830_ _02836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07262_ _02791_ _02781_ _02792_ _00148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06213_ cpu.spi.div_counter\[3\] _01871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09001_ _04007_ _04207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09224__A1 _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07193_ cpu.regs\[10\]\[2\] _02750_ _02751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06144_ _01337_ _01692_ _01802_ _01543_ _01803_ _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_5_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06075_ _00796_ _01735_ _01736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09903_ _00162_ clknet_leaf_88_wb_clk_i cpu.regs\[5\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05026_ _00721_ _00722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__07538__A1 _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09834_ _00093_ clknet_leaf_96_wb_clk_i cpu.regs\[14\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_81_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05013__A2 _00706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09765_ _00028_ clknet_leaf_79_wb_clk_i cpu.base_address\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_57_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06977_ _02237_ _02589_ _02590_ _02256_ _02591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08716_ _03461_ _03933_ _03946_ _03947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05928_ cpu.spi.divisor\[3\] _01133_ _01591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09696_ _04819_ _04821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08647_ cpu.IO_addr_buff\[6\] _03858_ _03892_ _03883_ _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05859_ cpu.IE _01299_ _01520_ _01522_ _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_1_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08578_ _02655_ _03827_ _03830_ _03832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08915__C _04106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07529_ _03009_ _01898_ _03010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_92_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05252__A2 _00919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09053__I _04150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06504__A2 _00955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04925__I _00626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09206__A1 _04374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_9_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08132__I _03456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06900_ _02523_ _02524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07880_ _02503_ _03236_ _03295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06831_ _02463_ _02442_ _02464_ _00045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09550_ cpu.PORTB_DDR\[0\] _04697_ _04698_ _04699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06762_ _01525_ _02400_ _02406_ _02408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05713_ cpu.uart.divisor\[1\] _01377_ _01378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08501_ _03776_ _03778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09481_ _04647_ cpu.pwm_counter\[0\] _03586_ cpu.pwm_top\[1\] _04648_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06693_ _00622_ _02345_ _02346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09693__A1 _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08432_ _02965_ _03668_ _03680_ _03720_ _03677_ _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_05644_ _01309_ _01310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_34_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05575_ _01027_ _01240_ _01241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08248__A2 _03551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08363_ _03662_ _03663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07314_ _02825_ _02826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08294_ _02454_ _03613_ _03614_ _00358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_116_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07245_ _02779_ _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_33_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07176_ _02739_ _00115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06127_ cpu.pwm_top\[6\] _01249_ _01786_ _01418_ _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_113_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06058_ cpu.timer_top\[13\] _01411_ _01251_ _01719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05009_ _00705_ _00706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_6_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09817_ _00076_ clknet_leaf_95_wb_clk_i _00005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09748_ _00747_ _04835_ _04862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_69_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08926__B _03442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09679_ _04803_ _04804_ _01542_ _04805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_95_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_95_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_96_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_24_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_24_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_92_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput19 io_in[2] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_107_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_70_Left_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06025__I1 cpu.regs\[13\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05084__S1 _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09511__I _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07686__B1 _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05360_ _01025_ _01026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05291_ _00922_ _00956_ _00959_ _00960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_43_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07030_ cpu.uart.receive_div_counter\[2\] _02630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_11_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08981_ _04179_ _04177_ _04185_ _04186_ _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_11_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07932_ _03308_ _03333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08797__I _03839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07863_ _03273_ _03280_ _03281_ _00260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_39_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09602_ _03618_ _04733_ _00547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06814_ _02450_ _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09533_ net82 _04682_ _04683_ _04687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07794_ cpu.uart.div_counter\[11\] _03221_ _03225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06745_ cpu.rom_data_dist _02393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06676_ _02321_ _00578_ _01920_ _02329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_09464_ _04630_ _04628_ _04635_ _03398_ _00507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__05527__I0 net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09395_ _04576_ _04578_ _00495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05627_ cpu.regs\[8\]\[7\] cpu.regs\[9\]\[7\] cpu.regs\[10\]\[7\] cpu.regs\[11\]\[7\]
+ _01285_ _01286_ _01293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_08415_ _02960_ _03706_ _03707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08346_ _02462_ _03643_ _03647_ _03648_ _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_116_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05558_ _00591_ _00590_ _01068_ _01224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08277_ _01073_ _02432_ _03602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05489_ _01145_ _01155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07228_ cpu.regs\[8\]\[2\] _02769_ _02770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07159_ cpu.regs\[12\]\[7\] _02720_ _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10170_ _00428_ clknet_leaf_50_wb_clk_i cpu.IO_addr_buff\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08500__I _03776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05066__S1 _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06955__I cpu.PC\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_69_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08632__A2 _03864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_78_Right_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06946__A2 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04957__A1 _00654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10299_ _00557_ clknet_leaf_108_wb_clk_i cpu.regs\[9\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_108_Left_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05057__S1 _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_87_Right_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06530_ _01296_ _02015_ _02187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06461_ net124 _02117_ _02118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_44_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05412_ _01077_ _01071_ _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08200_ _03536_ _03541_ _03548_ _03510_ _03549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XPHY_EDGE_ROW_117_Left_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09180_ _04071_ _04379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06392_ _02020_ _02026_ _02049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05343_ _01008_ _01009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08131_ _02454_ _03481_ _03483_ _00326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08062_ cpu.orig_PC\[0\] _03428_ _03430_ _03435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05274_ cpu.regs\[12\]\[4\] cpu.regs\[13\]\[4\] cpu.regs\[14\]\[4\] cpu.regs\[15\]\[4\]
+ _00890_ _00838_ _00943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_113_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_96_Right_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05988__A3 _01126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07013_ _02610_ _02621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_113_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08964_ _02389_ _04135_ _04164_ _04170_ _04171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07915_ cpu.uart.receive_buff\[4\] _03321_ _03316_ cpu.uart.receive_buff\[3\] _03322_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08895_ _01330_ _01937_ _04103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07846_ _03263_ _03267_ _03242_ _00257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input17_I io_in[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_04989_ _00687_ cpu.needs_timer_interrupt _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07777_ _03146_ _03209_ _03211_ _03212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09516_ _03798_ _04672_ _04676_ _00518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_108_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06728_ _00936_ _02377_ _02379_ _02380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09447_ cpu.ROM_spi_dat_out\[5\] _04579_ _04606_ _04621_ _04622_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_93_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06659_ cpu.startup_cycle\[3\] _02312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09378_ _03057_ _04561_ _04564_ _04565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__06873__A1 _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08329_ cpu.timer_top\[8\] _03637_ _03638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08378__A1 cpu.timer_capture\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10222_ _00480_ clknet_leaf_74_wb_clk_i cpu.PC\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__04939__A1 _00637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10153_ _00412_ clknet_leaf_16_wb_clk_i cpu.timer_div\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09326__I _04520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10084_ _00343_ clknet_leaf_118_wb_clk_i cpu.toggle_ctr\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08853__A2 _01273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06864__A1 cpu.timer_capture\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input9_I io_in[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07700_ _03125_ _03126_ _03143_ _03148_ _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_05961_ net43 _01020_ _01623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08680_ _03909_ _00729_ _03918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_04912_ _00584_ _00599_ _00614_ _00615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_05892_ _00741_ _01534_ _01536_ _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07631_ _03088_ _03089_ _00220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07562_ cpu.spi.data_out_buff\[5\] _03011_ _03026_ _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08296__B _03615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09301_ cpu.last_addr\[13\] _04491_ _04496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06513_ _02065_ _02169_ _02170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07493_ cpu.timer\[1\] _02977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_09232_ _04206_ _04426_ _04427_ _04429_ _03836_ _04430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_06444_ _02077_ _02099_ _02100_ _02101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_29_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09163_ _02209_ _03903_ _04363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06375_ _00745_ _02031_ _02032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_16_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05326_ _00991_ _00992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08114_ cpu.toggle_clkdiv _03472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09094_ _04175_ _04293_ _04296_ _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08045_ _03420_ _03413_ _03422_ _00301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06083__A2 _00979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05257_ cpu.regs\[4\]\[3\] cpu.regs\[5\]\[3\] cpu.regs\[6\]\[3\] cpu.regs\[7\]\[3\]
+ _00834_ _00926_ _00927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_31_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05188_ cpu.regs\[4\]\[0\] cpu.regs\[5\]\[0\] cpu.regs\[6\]\[0\] cpu.regs\[7\]\[0\]
+ _00858_ _00859_ _00860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_09996_ _00255_ clknet_leaf_23_wb_clk_i cpu.uart.counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08947_ _04113_ _04154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08878_ _04084_ _04085_ _04086_ _04078_ _04087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_07829_ cpu.uart.counter\[3\] _03252_ _03151_ _03253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08532__A1 _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10205_ _00463_ clknet_leaf_69_wb_clk_i cpu.last_addr\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06901__C _02524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10136_ _00395_ clknet_leaf_5_wb_clk_i cpu.timer_capture\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10067_ _00326_ clknet_leaf_117_wb_clk_i cpu.toggle_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__08523__A1 _00986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_32_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06534__B1 _02040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06160_ net58 cpu.PORTA_DDR\[7\] _01192_ _01819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_25_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09675__B _00913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05111_ cpu.regs\[4\]\[6\] cpu.regs\[5\]\[6\] cpu.regs\[6\]\[6\] cpu.regs\[7\]\[6\]
+ _00799_ _00800_ _00802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_13_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06091_ _01751_ _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_111_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05042_ _00736_ _00737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07565__A2 _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09850_ _00109_ clknet_leaf_104_wb_clk_i cpu.regs\[12\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08801_ _04010_ _04012_ _04013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09781_ _00044_ clknet_leaf_26_wb_clk_i cpu.uart.divisor\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06993_ _02283_ _02554_ _02605_ _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08732_ _03959_ _00451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05944_ _00949_ _01276_ _01518_ _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08663_ _02382_ _03900_ _03905_ _00436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08514__A1 cpu.spi.divisor\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05875_ _01537_ _01538_ _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07614_ _03001_ _03079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08594_ cpu.orig_IO_addr_buff\[0\] _03842_ _03845_ _00986_ _03846_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_105_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07545_ _02489_ _03022_ _03023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07476_ cpu.timer\[9\] _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09215_ _02207_ _04150_ _04413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06427_ _00952_ _02017_ _02001_ _00945_ _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_106_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05669__I _01333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05500__A1 _01114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09146_ _04339_ _04341_ _04345_ _04346_ _04347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_16_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06358_ cpu.multiplier.a\[3\] _00767_ _02015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09077_ _03453_ _01058_ _04280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05309_ _00974_ _00976_ _00977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06289_ cpu.multiplier.a\[0\] _01946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_49_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_49_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08028_ _02455_ _03410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_116_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09979_ _00238_ clknet_leaf_29_wb_clk_i cpu.uart.div_counter\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05111__S0 _00799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08505__A1 _02525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_105_Right_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08664__B _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_116_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06631__C _01761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10119_ _00378_ clknet_leaf_10_wb_clk_i cpu.timer\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09514__I _04674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05660_ _01325_ _01326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05591_ cpu.toggle_top\[0\] _01171_ _01173_ _01256_ _01257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_58_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07330_ _02835_ _00173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09000_ _04034_ _04206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05489__I _01145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07261_ cpu.regs\[7\]\[5\] _02786_ _02792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07192_ _02744_ _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06212_ _01354_ _01869_ _01870_ _00020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06143_ _01451_ _01691_ _01803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06074_ _01156_ _01734_ _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09902_ _00161_ clknet_leaf_87_wb_clk_i cpu.regs\[5\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05025_ cpu.regs\[8\]\[1\] cpu.regs\[9\]\[1\] cpu.regs\[10\]\[1\] cpu.regs\[11\]\[1\]
+ _00697_ _00698_ _00721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05549__A1 cpu.uart.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09833_ _00092_ clknet_leaf_100_wb_clk_i cpu.regs\[14\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09764_ _00027_ clknet_leaf_79_wb_clk_i cpu.base_address\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_57_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05952__I _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06976_ net19 _02558_ _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05927_ cpu.uart.dout\[3\] _01022_ _01589_ _01590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09695_ _04819_ _04820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08715_ _03942_ cpu.regs\[3\]\[1\] _03946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08646_ _03838_ _03890_ _03891_ _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05858_ _01450_ _01521_ _01298_ _01522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_1_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08577_ _03801_ _03826_ _03831_ _00424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05721__A1 _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05789_ _01435_ _01454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_37_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07528_ cpu.spi.counter\[0\] _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07459_ cpu.timer_div\[6\] _02941_ cpu.timer_div_counter\[7\] _02935_ _02942_ _02943_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_118_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09129_ cpu.orig_PC\[8\] _04244_ _04330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09215__A2 _04150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07226__A1 _02717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06732__B _02379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06958__I _01938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09151__A1 _00696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09454__A2 _04592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08965__B2 _03836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05779__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06291__I2 _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06830_ cpu.uart.divisor\[6\] _02435_ _02457_ _02464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05772__I _00726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06761_ _02382_ _02402_ _02407_ _00032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06692_ cpu.spi_clkdiv _02294_ _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05712_ _01374_ _01377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09142__A1 _03848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08500_ _03776_ _03777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09480_ cpu.pwm_top\[0\] _04647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05643_ _01094_ _01309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09693__A2 _02729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08431_ cpu.timer\[12\] _03719_ _03720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_102_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05574_ _01239_ _01030_ _01240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_62_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08362_ _03651_ _03662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07313_ _02824_ _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08293_ cpu.pwm_top\[4\] _03603_ _03609_ _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07244_ _02779_ _02780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_33_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07175_ _01679_ cpu.regs\[11\]\[4\] _02731_ _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08956__B2 _04162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06126_ _01783_ _01784_ _01785_ _01786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_113_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06057_ _01713_ _01715_ _01717_ _01718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05008_ cpu.regs\[8\]\[0\] cpu.regs\[9\]\[0\] cpu.regs\[10\]\[0\] cpu.regs\[11\]\[0\]
+ _00703_ _00704_ _00705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_6_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09816_ _00075_ clknet_leaf_94_wb_clk_i _00004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_06959_ _02573_ _02574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09747_ _01613_ _02555_ _04860_ _04861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08993__I _04106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08731__I1 cpu.ROM_addr_buff\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09678_ _00712_ _00873_ _01459_ _04804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09684__A2 _01733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08629_ _03862_ _03876_ _03877_ _03878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_65_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_64_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_64_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_64_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05305__S0 _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09372__A1 _04558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08175__A2 cpu.toggle_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06186__A1 _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05933__A1 _01593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__04936__I _00636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05290_ _00911_ _00958_ _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08143__I cpu.toggle_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06413__A2 cpu.multiplier.a\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08980_ _04154_ _04186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07931_ _03327_ _03332_ _00277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07862_ cpu.uart.data_buff\[3\] _03276_ _03041_ _03281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09601_ net75 _04727_ _04732_ _04583_ _04733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06813_ _00933_ _02450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05224__I0 cpu.regs\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09532_ _03823_ _04681_ _04686_ _00524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07793_ _03214_ _03224_ _00247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06744_ _02373_ _02388_ _02392_ _00030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06675_ _02320_ _02323_ _02327_ _02328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08713__I1 cpu.ROM_addr_buff\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09463_ _04628_ _04634_ _04630_ _04635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05527__I1 cpu.PORTA_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09394_ _02478_ _04577_ _04578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05626_ _00857_ _01291_ _00887_ _01292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_08414_ _03702_ _03698_ _03706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08345_ _03159_ _03648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05557_ _01222_ _01223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_80_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08276_ _03585_ _03601_ _00353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05488_ _01153_ _01154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_116_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07227_ _02763_ _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08053__I _03407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07158_ _02727_ _00109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06109_ net13 _01370_ _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07089_ _02381_ _02683_ _02420_ _00084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_100_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_111_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_111_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_4_4_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05391__A2 _00657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05230__I3 cpu.regs\[11\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06891__A2 _02513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08093__A1 _02597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06904__C _02524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09593__A1 cpu.ROM_spi_mode vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10298_ _00556_ clknet_leaf_108_wb_clk_i cpu.regs\[9\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07307__I _01814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05271__B _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06460_ _01945_ _02116_ _02117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_34_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07042__I _01209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05411_ _00585_ _01076_ _01077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_44_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06391_ _02020_ _02026_ _02048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08130_ cpu.toggle_top\[4\] _03482_ _03477_ _03483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08084__A1 _02214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05342_ _00606_ _01007_ _01008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08061_ _03401_ _03434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05273_ _00831_ _00941_ _00848_ _00942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_99_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07012_ cpu.toggle_top\[12\] _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_70_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09584__A1 cpu.PORTA_DDR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08963_ _00728_ _04166_ _04168_ _04169_ _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07914_ _03312_ _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08894_ _00679_ _04101_ _04102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07198__I0 _02753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07845_ cpu.uart.counter\[3\] _03264_ _03266_ _03267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04988_ cpu.TIE _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07776_ _03146_ _03210_ _03204_ _03211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__06570__A1 _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09515_ net63 _04673_ _04675_ _04676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06727_ _02378_ _02379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09446_ _04562_ _04571_ _04621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_108_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06658_ _02306_ _02311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09377_ _04562_ _04563_ _02313_ _04564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05609_ _01272_ _01274_ _01275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_47_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06589_ _01799_ _02131_ _02040_ _01296_ _02245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_105_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08328_ _03635_ _03637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_105_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07822__A1 _03094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08259_ _03584_ cpu.pwm_counter\[1\] _03589_ _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10221_ _00479_ clknet_leaf_75_wb_clk_i cpu.PC\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10152_ _00411_ clknet_leaf_9_wb_clk_i cpu.timer_div\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08511__I _03776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10083_ _00342_ clknet_leaf_113_wb_clk_i cpu.toggle_ctr\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06031__I _01691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_22_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08302__A2 _03613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06313__A1 _01952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09566__A1 _02538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_61_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05960_ net55 cpu.PORTA_DDR\[4\] _01192_ _01622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_04911_ _00601_ _00606_ _00613_ _00614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_49_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05891_ _01168_ _01552_ _01554_ _00015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07630_ cpu.spi.data_in_buff\[5\] _03083_ _03085_ cpu.spi.data_in_buff\[6\] _03089_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06876__I _00981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07561_ cpu.spi.data_out_buff\[6\] _03021_ _03035_ _03036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09300_ cpu.last_addr\[12\] cpu.ROM_addr_buff\[12\] _04494_ _04495_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_75_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06512_ _01798_ _02018_ _02066_ _01295_ _02169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07492_ cpu.timer\[4\] _02976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09231_ _00680_ _04410_ _04428_ _04404_ _04429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06443_ _02062_ net126 _02100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09162_ _04334_ _04335_ _04361_ _04362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_8_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06374_ _00953_ _01992_ _01994_ _00945_ _02031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_28_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08113_ _02440_ _03396_ _00320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05325_ cpu.IO_addr_buff\[1\] _00990_ _00991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09093_ _04267_ _04276_ _04295_ _04235_ _04207_ _04296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_71_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08044_ cpu.orig_IO_addr_buff\[7\] _03418_ _03421_ _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05020__I _00703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05256_ _00005_ _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09557__A1 _02529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05187_ _00838_ _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__08780__A2 _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09995_ _00254_ clknet_leaf_25_wb_clk_i cpu.uart.counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08946_ _04150_ _04134_ _04151_ _04152_ _04153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_71_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08877_ cpu.br_rel_dest\[0\] _04084_ _04086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07828_ cpu.uart.counter\[2\] _03252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05346__A2 _00999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06786__I _02425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07759_ cpu.uart.div_counter\[4\] _03196_ _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_106_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08296__A1 cpu.pwm_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09429_ cpu.ROM_spi_dat_out\[2\] _04598_ _04603_ _04608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_81_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08048__A1 _01303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05282__A1 _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10204_ _00462_ clknet_leaf_68_wb_clk_i cpu.last_addr\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05585__A2 _01073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10135_ _00394_ clknet_leaf_5_wb_clk_i cpu.timer_capture\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10066_ _00325_ clknet_leaf_2_wb_clk_i cpu.toggle_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_82_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05105__I _00796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08287__A1 _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06837__A2 _02432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05110_ cpu.regs\[0\]\[6\] _00798_ cpu.regs\[2\]\[6\] cpu.regs\[3\]\[6\] _00799_
+ _00800_ _00801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_96_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06090_ _01307_ _01729_ _01748_ _01750_ _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__07262__A2 _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09539__A1 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05041_ cpu.regs\[8\]\[2\] cpu.regs\[9\]\[2\] cpu.regs\[10\]\[2\] cpu.regs\[11\]\[2\]
+ _00716_ _00731_ _00736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_40_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06222__B1 cpu.spi.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08800_ _04011_ _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09780_ _00043_ clknet_leaf_17_wb_clk_i cpu.uart.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06773__A1 _02416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06992_ _02584_ _02604_ _02605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07923__C _02439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08731_ _03958_ cpu.ROM_addr_buff\[12\] _03952_ _03959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05943_ _00918_ _01516_ _01605_ _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08662_ _03903_ _03901_ _03904_ _03905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07613_ _03077_ _03078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05874_ _01528_ _01530_ _01535_ _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_88_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08593_ _03844_ _03845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05443__C _00911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07544_ _03006_ _03022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05015__I _00711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07325__I0 _02818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07475_ cpu.timer\[10\] _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09214_ _04197_ _04410_ _04411_ _04199_ _04412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_48_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06426_ _00746_ _02082_ _02083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05500__A2 _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09145_ _00661_ _04346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06357_ _00744_ _00767_ _02014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09076_ _04277_ _04278_ _04279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05308_ _00843_ _00975_ _00849_ _00976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06288_ _01944_ _01945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_31_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05264__A1 _00911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08027_ _01048_ _03402_ _03409_ _00296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05239_ _00908_ _00909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_116_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08061__I _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09978_ _00237_ clknet_leaf_29_wb_clk_i cpu.uart.div_counter\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06764__A1 _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05111__S1 _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_89_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_89_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08929_ _00664_ _00612_ _04136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_18_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_18_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08992__A2 _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10118_ _00377_ clknet_leaf_11_wb_clk_i cpu.timer_top\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10049_ _00308_ clknet_leaf_63_wb_clk_i cpu.orig_PC\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09016__B _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_11_Left_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05590_ _01246_ _01250_ _01255_ _01256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_85_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07260_ _01751_ _02791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07191_ _02717_ _02746_ _02749_ _00120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06211_ cpu.regs\[15\]\[7\] _01553_ _01870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06142_ _00810_ _01801_ _01802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_53_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06073_ _01326_ _01733_ _01734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09901_ _00160_ clknet_leaf_86_wb_clk_i cpu.regs\[5\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05024_ _00718_ _00719_ _00707_ _00720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06994__A1 _02271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09832_ _00091_ clknet_leaf_100_wb_clk_i cpu.regs\[14\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09763_ _00026_ clknet_leaf_43_wb_clk_i net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08714_ _03945_ _00447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_4_9_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06975_ _02030_ _02588_ _02589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05926_ _01588_ _01589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09694_ _04818_ _04819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xrebuffer10 _02114_ net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08645_ _02421_ _03851_ _03891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05857_ _01518_ _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_1_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07171__A1 cpu.regs\[11\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08576_ cpu.uart.divisor\[13\] _03827_ _03830_ _03831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05721__A2 _01142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07527_ _03006_ _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05788_ _01340_ _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08671__A1 _03433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08056__I _03410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07458_ _01496_ cpu.timer_div_counter\[2\] _02941_ cpu.timer_div\[6\] _02942_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_118_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07389_ _02882_ _02222_ _02883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_45_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06409_ _02001_ _02066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_118_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09128_ _04328_ _04329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09059_ _02419_ _04256_ _04261_ _04262_ _04263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05627__I3 cpu.regs\[11\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06985__A1 _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output60_I net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07162__A1 _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06907__C _02524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06268__A3 _00663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08662__A1 _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05476__A1 _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07217__A2 _01813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05079__I1 _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06976__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09525__I _04680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput90 net90 sram_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06728__A1 _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07940__A3 cpu.uart.receive_div_counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06760_ _01430_ _02401_ _02406_ _02407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06691_ _02295_ _02343_ _02344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05711_ _01372_ _01373_ _01375_ _01376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05642_ _01169_ _01170_ _01301_ _01305_ _01307_ _01308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_08430_ cpu.timer\[11\] _03715_ _03719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_102_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05573_ _01019_ _01239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_62_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08361_ _03653_ _03659_ _03661_ _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08653__A1 _03885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07312_ _02711_ _02777_ _02824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08292_ _03602_ _03613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07243_ _02778_ _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05011__S0 _00703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07174_ _02722_ _02732_ _02738_ _00114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06125_ cpu.timer_top\[14\] _01598_ _01251_ _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_68_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06056_ _01716_ _01243_ _01598_ _01717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_113_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05007_ _00001_ _00704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09815_ _00011_ clknet_leaf_57_wb_clk_i cpu.instr_cycle\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09746_ _02584_ _04859_ _04860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06958_ _01938_ _02573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_69_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05909_ net29 _01310_ _01311_ _01572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09677_ _01437_ _00884_ _04803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_68_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08628_ _01573_ _03867_ _03877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07144__A1 _02717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06889_ cpu.timer\[7\] _02514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_96_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08559_ cpu.uart.divisor\[8\] _03818_ _03802_ _03819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08644__B2 _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05458__A1 _01121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05002__S0 _00697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06743__B _02391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05305__S1 _00899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_33_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_33_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_20_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08389__C _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08883__A1 _04070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer1 _02058_ net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_11_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07930_ _03328_ _03309_ _03331_ _03332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09255__I _04103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07861_ cpu.uart.data_buff\[2\] _03264_ _03279_ _03280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07374__A1 _00696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09600_ _04568_ _04728_ _02311_ _04731_ _04732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_07792_ cpu.uart.div_counter\[10\] _03178_ _03222_ _03223_ _03224_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06812_ _02447_ _02436_ _02449_ _00041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_39_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09531_ net81 _04682_ _04683_ _04686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06743_ _02389_ _02377_ _02391_ _02392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06674_ _02316_ _02324_ _02326_ _02327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_09462_ _00567_ _04633_ _04634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_47_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09393_ _04547_ _04555_ _04572_ _04577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_46_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05625_ cpu.regs\[12\]\[7\] cpu.regs\[13\]\[7\] cpu.regs\[14\]\[7\] cpu.regs\[15\]\[7\]
+ _01285_ _01286_ _01291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_08413_ _03663_ _03704_ _03705_ _00386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05556_ _01221_ _01222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08344_ cpu.timer_top\[14\] _03644_ _03647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05487_ _00650_ _01103_ _01152_ _00882_ _01153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_6_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08275_ cpu.pwm_counter\[7\] _03599_ _03601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07226_ _02717_ _02765_ _02768_ _00136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08334__I _02523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05860__A1 _01304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_1_0_wb_clk_i clknet_0_wb_clk_i clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07157_ _01816_ cpu.regs\[12\]\[6\] _02713_ _02727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06108_ _01122_ _01766_ _01767_ _01052_ _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_30_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07088_ _02375_ _02683_ _02417_ _00083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06039_ net64 _01195_ _01700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_12_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09729_ _01466_ _02554_ _04835_ _04844_ _04845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_97_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08865__A1 _04070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05223__S0 _00891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08617__A1 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09593__A2 _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_51_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05603__A1 _01257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10297_ _00555_ clknet_leaf_109_wb_clk_i cpu.regs\[9\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04947__I net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08856__A1 _04008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05410_ _00990_ _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_68_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08608__A1 _03585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06390_ _02037_ _02044_ _02046_ _02047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_05341_ _01003_ _01006_ _01007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_clkbuf_leaf_90_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08060_ _03432_ _03433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_70_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05272_ cpu.regs\[8\]\[4\] cpu.regs\[9\]\[4\] cpu.regs\[10\]\[4\] cpu.regs\[11\]\[4\]
+ _00834_ _00892_ _00941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_99_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07011_ _02451_ _02615_ _02619_ _00070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05842__A1 cpu.timer_top\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08962_ _00666_ _04169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07913_ _03213_ _03320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08893_ _04100_ _02430_ _04101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07844_ _03265_ _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07198__I1 cpu.regs\[10\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_3_Left_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_04987_ _00649_ _00623_ _00684_ _00629_ _00686_ _00008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_07775_ _03200_ _03210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09514_ _04674_ _04675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06726_ _00620_ _02378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08847__A1 _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09445_ _04620_ _00503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_108_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06657_ _02300_ _02306_ _02309_ _02310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_94_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05608_ _00636_ _01273_ _01274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09376_ _04548_ _04543_ _04563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06588_ _02192_ _02195_ _02243_ _02244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05539_ net21 _01189_ _01201_ _01204_ _01205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_08327_ _03635_ _03636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08064__I cpu.PC\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Left_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08258_ cpu.pwm_counter\[2\] _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09024__A1 _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07209_ _02760_ _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_76_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10220_ _00478_ clknet_leaf_75_wb_clk_i cpu.PC\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08189_ _03499_ _01723_ _02620_ _03489_ _03538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_100_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10151_ _00410_ clknet_leaf_16_wb_clk_i cpu.timer_div\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10082_ _00341_ clknet_leaf_112_wb_clk_i cpu.toggle_ctr\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_58_Left_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07338__A1 _01352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06010__A1 _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06313__A2 _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_67_Left_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_65_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_76_Left_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04910_ _00609_ _00612_ _00613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__06001__A1 _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05890_ cpu.regs\[15\]\[2\] _01553_ _01554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07560_ _02508_ _03022_ _03035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08829__A1 _01108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06511_ _02161_ _02164_ _02167_ _02168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_118_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09230_ _00748_ _04351_ _04428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09689__B _04814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07491_ cpu.timer\[3\] _02975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07501__A1 _01716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06442_ _02062_ net126 _02099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09161_ _04336_ _04361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_56_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06373_ _02008_ _02028_ _02029_ _02030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_16_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08112_ _02254_ _03404_ _03471_ _00319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09254__B2 _04162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09092_ _00798_ _04232_ _04294_ _04295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05324_ _00586_ _00990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06068__A1 _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05815__A1 net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08043_ _03410_ _03421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05301__I _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09006__A1 cpu.PC\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05255_ _00923_ _00924_ _00830_ _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_101_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05186_ _00835_ _00858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09994_ _00253_ clknet_leaf_17_wb_clk_i cpu.uart.has_byte vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08945_ _04115_ _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_71_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input22_I io_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08876_ _03432_ _03847_ _04085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_98_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07827_ _03248_ _03152_ _03251_ _03158_ _00254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07758_ _03117_ _03191_ _03196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08059__I cpu.PC\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06709_ _02349_ _02352_ _02361_ _02362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_94_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07689_ cpu.uart.div_counter\[10\] _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09428_ cpu.ROM_spi_dat_out\[1\] _04579_ _04605_ _04606_ _04607_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_66_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09359_ cpu.startup_cycle\[1\] _04548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_81_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06059__A1 cpu.pwm_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output90_I net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05282__A2 _00950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10203_ _00461_ clknet_leaf_68_wb_clk_i cpu.last_addr\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10134_ _00393_ clknet_leaf_3_wb_clk_i cpu.timer\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10065_ _00324_ clknet_leaf_2_wb_clk_i cpu.toggle_top\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05121__I _00811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05040_ _00707_ _00735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_84_Left_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09691__C _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06991_ _02579_ _02599_ _02603_ _02604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08730_ _03469_ _03949_ _03957_ _03958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05942_ _01602_ _01603_ _01604_ _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08661_ _03829_ _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05873_ _01098_ _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07612_ _01896_ _01892_ _03077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_93_Left_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08592_ _00667_ _03843_ _03844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09475__A1 net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07543_ _01897_ _03021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_52_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07474_ cpu.timer_top\[10\] _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_118_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09213_ cpu.orig_PC\[11\] _03841_ _04411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06425_ _01730_ _01992_ _01994_ _01797_ _02082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_98_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09144_ _00984_ _04192_ _04344_ _04154_ _04345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_8_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05031__I _00726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06356_ _02011_ _02012_ _02003_ _02013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09075_ cpu.PC\[5\] _00636_ _04251_ _04278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05307_ cpu.regs\[12\]\[5\] cpu.regs\[13\]\[5\] cpu.regs\[14\]\[5\] cpu.regs\[15\]\[5\]
+ _00891_ _00893_ _00975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_06287_ _01943_ _01944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05966__I cpu.uart.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08026_ cpu.orig_IO_addr_buff\[2\] _03408_ _03303_ _03409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05238_ cpu.base_address\[3\] _00908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_116_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05169_ _00833_ _00840_ _00841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_40_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09977_ _00236_ clknet_leaf_26_wb_clk_i cpu.uart.busy vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06764__A2 _02400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08928_ _04134_ _04135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08859_ _04068_ _00469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_4_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_58_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_58_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_79_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_14_0_wb_clk_i clknet_0_wb_clk_i clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_91_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10117_ _00376_ clknet_leaf_11_wb_clk_i cpu.timer_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10048_ _00307_ clknet_leaf_55_wb_clk_i cpu.orig_PC\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08680__A2 _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06210_ _01868_ _01869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07190_ cpu.regs\[10\]\[1\] _02747_ _02749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06141_ _00880_ _01800_ _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_5_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08162__I cpu.toggle_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06072_ _01732_ _01733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05023_ cpu.regs\[4\]\[1\] cpu.regs\[5\]\[1\] cpu.regs\[6\]\[1\] cpu.regs\[7\]\[1\]
+ _00697_ _00698_ _00719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_09900_ _00159_ clknet_leaf_86_wb_clk_i cpu.regs\[5\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09831_ _00090_ clknet_leaf_102_wb_clk_i cpu.regs\[14\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06974_ _02587_ _02051_ _02588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09762_ _00025_ clknet_leaf_82_wb_clk_i cpu.regs\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_08713_ _03944_ cpu.ROM_addr_buff\[8\] _03937_ _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08111__B _03467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05925_ _00992_ _00997_ _01025_ _00989_ _01588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_57_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08499__A2 _01040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09693_ _02546_ _02729_ _04818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xrebuffer11 _00863_ net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08644_ cpu.orig_IO_addr_buff\[6\] _03842_ _03845_ _01808_ _03890_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05856_ _01471_ _01517_ _01519_ _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08575_ _03829_ _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_95_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05787_ _01437_ _01449_ _01452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_1_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07526_ _03006_ _03007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08120__A1 _02427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08671__A2 _00649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07457_ cpu.timer_div_counter\[6\] _02941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_118_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07388_ _02208_ _02882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06408_ _00782_ _02065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_118_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09127_ _04325_ _04327_ _04328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06339_ _00853_ _01993_ _01995_ _00914_ _01996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_105_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_105_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07397__B _02890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08072__I _03407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09058_ _04113_ _04262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06434__A1 _00854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08009_ _03392_ _03394_ _03395_ _00292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06985__A2 _02569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04996__B2 _00694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06737__A2 _02385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05096__S1 _00786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output53_I net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07698__B1 _02441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07162__A2 _02729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05476__A2 _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06425__A1 _01730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05079__I2 _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06425__B2 _01797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06976__A2 _02558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04987__A1 _00649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08710__I _03908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput80 net80 io_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput91 net91 sram_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05400__A2 _01065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_qcpu_98 io_oeb[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_06690_ _02304_ _02310_ _02315_ _02342_ _02343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__07770__B _00645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05710_ _01374_ _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05641_ _01306_ _01307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_77_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08360_ cpu.timer_capture\[0\] _03660_ _03615_ _03661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_102_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05572_ _01231_ _01234_ _01237_ _01238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07311_ _02807_ _02812_ _02823_ _00166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_3_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_3_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_34_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08291_ _02451_ _03604_ _03612_ _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_73_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07242_ _01165_ _02777_ _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05011__S1 _00704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07173_ cpu.regs\[11\]\[3\] _02736_ _02738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09602__A1 _03618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08106__B _03467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06124_ cpu.timer_top\[6\] _01500_ _01241_ _01784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06416__B2 _00854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06055_ cpu.timer_top\[5\] _01716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_113_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06341__S _01950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05006_ _00000_ _00703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07664__C _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09814_ _00010_ clknet_leaf_54_wb_clk_i cpu.instr_cycle\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_6_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06957_ _02570_ _02571_ _02572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09669__B2 _01041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09745_ _02574_ _04855_ _04858_ _04859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_68_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06888_ _02465_ _02513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09676_ _01862_ _04029_ _04802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05908_ _01463_ _01570_ _01571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_68_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08627_ cpu.orig_IO_addr_buff\[3\] _03864_ _03865_ _00958_ _03876_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05839_ cpu.timer_top\[2\] _01243_ _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05155__A1 net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08558_ _03816_ _03818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07509_ _02956_ cpu.timer\[8\] _02947_ _02968_ _02993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_37_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08489_ _03760_ _03767_ _03768_ _00399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_107_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05002__S1 _00698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_30_Left_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_41_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_73_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_73_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_99_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05394__A1 _01057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08332__A1 _02525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08883__A2 _04091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_80_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer2 _02238_ net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_51_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09536__I _04680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07860_ _02480_ _03278_ _03279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07791_ _03138_ _03219_ _03223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06811_ _02448_ _02437_ _02391_ _02449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_39_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09530_ _03820_ _04681_ _04685_ _00523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06742_ _02390_ _02391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_64_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09461_ _04631_ _04632_ _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06673_ _01913_ _02325_ _02326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_19_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09392_ _04556_ _04572_ _04547_ _04576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_65_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_47_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05624_ _00857_ _01289_ _00897_ _01290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08412_ cpu.timer_capture\[8\] _03652_ _03675_ _03705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05555_ _01010_ _01220_ _01221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_46_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08343_ _02459_ _03643_ _03646_ _03641_ _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_74_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08274_ _03598_ _03600_ _00352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_116_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05486_ _01151_ _01145_ _01102_ _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_61_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07225_ cpu.regs\[8\]\[1\] _02766_ _02768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07156_ _02725_ _02715_ _02726_ _00108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06107_ net4 _01199_ _01767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07087_ _02414_ _02683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06038_ _01364_ _01697_ _01698_ _01198_ _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08350__I _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05376__A1 _01040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07989_ cpu.uart.receive_div_counter\[12\] _03376_ _03372_ _03379_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_2
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09728_ _04838_ _04843_ _02553_ _04844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09659_ _04785_ _04783_ _04786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_69_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_8_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05223__S1 _00893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07053__B2 cpu.uart.divisor\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10296_ _00554_ clknet_leaf_109_wb_clk_i cpu.regs\[9\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08305__A1 _02390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06316__B1 _01971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05340_ _01005_ _01006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05271_ _00831_ _00939_ _00007_ _00940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_99_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07010_ cpu.toggle_top\[11\] _02612_ _02616_ _02619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07044__B2 cpu.uart.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07044__A1 cpu.uart.divisor\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08961_ _04167_ _04135_ _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07912_ _03243_ _03319_ _00271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08892_ _00651_ _00638_ _00639_ _00635_ _04100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_07843_ _03156_ _03151_ _03265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_04986_ _00685_ _00686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07774_ _03157_ _03207_ _03200_ _03208_ _03209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_79_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09513_ _03607_ _04674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06725_ _02372_ _02377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08847__A2 _01694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09444_ cpu.ROM_spi_dat_out\[5\] _04609_ _04619_ _04527_ _04620_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06656_ _02296_ _02308_ _02309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_108_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06858__A1 cpu.timer_capture\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_74_Right_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05607_ _01059_ _01273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09375_ _02359_ _04562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05530__A1 cpu.PORTB_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06587_ _00815_ _00948_ _02196_ _02243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05538_ _01203_ _01204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08345__I _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08326_ _01240_ _02433_ _03635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_104_Left_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08257_ _03001_ _03588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05469_ _00993_ _01125_ _01135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_61_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06086__A2 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08188_ _03493_ _03498_ _03501_ _03537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07208_ _01148_ _01154_ _02759_ _02543_ _02760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_104_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07139_ _02713_ _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07035__B2 _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_83_Right_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08080__I _03403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05597__A1 _01110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10150_ _00409_ clknet_leaf_12_wb_clk_i cpu.spi.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08013__C _03398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10081_ _00340_ clknet_leaf_114_wb_clk_i cpu.toggle_ctr\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_113_Left_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_87_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06561__A3 cpu.PC\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_92_Right_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_84_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05521__A1 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10279_ _00537_ clknet_leaf_14_wb_clk_i cpu.PORTB_DDR\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08858__C _02439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04958__I _00657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08829__A2 _01942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07490_ cpu.timer\[5\] _02974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_06510_ _01963_ _02141_ _02166_ _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_29_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06441_ _02088_ _02094_ _02097_ _02098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_29_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_100_Right_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_84_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09160_ _04243_ _04358_ _04359_ _04246_ _04360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06372_ _02027_ _02010_ _02013_ _02029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08111_ cpu.orig_PC\[13\] _03464_ _03467_ _03471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09091_ _04268_ _04276_ _04294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05323_ _00598_ _00989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07002__C _02542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08042_ cpu.IO_addr_buff\[7\] _03420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05254_ cpu.regs\[8\]\[3\] cpu.regs\[9\]\[3\] cpu.regs\[10\]\[3\] cpu.regs\[11\]\[3\]
+ _00889_ _00837_ _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_43_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07017__A1 _01723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05185_ _00842_ _00857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09993_ _00252_ clknet_leaf_28_wb_clk_i cpu.uart.div_counter\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08944_ _04131_ _04149_ _04151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_71_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08517__A1 _02538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08875_ _00678_ _00672_ _04084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07826_ _03248_ _03249_ _03250_ _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07244__I _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input15_I io_in[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07757_ _03177_ _03195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04969_ _00639_ _00668_ _00669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06708_ _02353_ _02358_ _02310_ _02360_ _02361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_39_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07688_ cpu.uart.div_counter\[0\] _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09427_ _02351_ _04596_ _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06639_ cpu.regs\[2\]\[7\] _01933_ _02293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09358_ _02299_ _04547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08309_ _03623_ _03624_ _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09289_ _01915_ _04483_ _04484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10202_ _00460_ clknet_leaf_68_wb_clk_i cpu.last_addr\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05114__S0 _00799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10133_ _00392_ clknet_leaf_2_wb_clk_i cpu.timer\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08508__A1 cpu.spi.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05990__B2 _01137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05990__A1 _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10064_ _00323_ clknet_leaf_2_wb_clk_i cpu.toggle_top\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07154__I _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06926__C _02542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06222__A2 cpu.spi.divisor\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06990_ _02256_ _02600_ _02602_ _02603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input7_I io_in[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05941_ cpu.toggle_top\[11\] _01259_ _01261_ _01604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08660_ _00882_ _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05872_ _01528_ _01530_ _01535_ _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07611_ net16 _03076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08591_ _00651_ _01618_ _03843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09475__A2 _03551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07542_ _03013_ _03019_ _03020_ _00200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07473_ _02955_ cpu.timer\[9\] cpu.timer\[8\] _02956_ _02957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_118_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08109__B _03467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09212_ _04409_ _04410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06424_ _02053_ _02079_ _02080_ _02081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09143_ _02856_ _03849_ _04342_ _04343_ _04344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05312__I _00979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07238__A1 cpu.regs\[8\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06355_ _01997_ _02000_ _02012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_8_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05306_ _00965_ _00973_ _00974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_44_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09074_ cpu.PC\[5\] _00636_ _04277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06286_ _00714_ _01943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05237_ _00907_ net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08025_ _03407_ _03408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05264__A3 _00933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05168_ cpu.regs\[0\]\[1\] cpu.multiplier.a\[1\] cpu.regs\[2\]\[1\] cpu.regs\[3\]\[1\]
+ _00836_ _00839_ _00840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_40_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09976_ _00235_ clknet_leaf_39_wb_clk_i cpu.spi.counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05099_ cpu.regs\[8\]\[5\] cpu.regs\[9\]\[5\] cpu.regs\[10\]\[5\] cpu.regs\[11\]\[5\]
+ _00770_ _00786_ _00791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05272__I0 cpu.regs\[8\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05972__A1 cpu.spi.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08927_ _04132_ _04133_ _04134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08858_ _01427_ _03870_ _04036_ _04067_ _02439_ _04068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_07809_ cpu.uart.div_counter\[14\] _03230_ _03231_ _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_4_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08789_ cpu.last_addr\[12\] _03996_ _04003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09403__B _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_98_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_98_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_109_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_27_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_27_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_109_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06762__B _02406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06452__A2 _02072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07149__I _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05963__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10116_ _00375_ clknet_leaf_11_wb_clk_i cpu.timer_top\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10047_ _00306_ clknet_leaf_54_wb_clk_i cpu.orig_PC\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08901__A1 _04108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08968__A1 _04173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06140_ _01326_ _01799_ _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06071_ _01731_ _01732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05022_ cpu.regs\[0\]\[1\] _00714_ _00715_ cpu.regs\[3\]\[1\] _00716_ _00717_ _00718_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09830_ _00089_ clknet_leaf_100_wb_clk_i cpu.regs\[14\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09761_ _00024_ clknet_leaf_82_wb_clk_i cpu.regs\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_06973_ _02052_ _02587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08712_ _02856_ _03933_ _03943_ _03944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05924_ _01582_ _01584_ _01586_ _01587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_57_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09692_ _04817_ _00553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xrebuffer12 _02075_ net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05706__A1 _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08643_ _03885_ _03889_ _00432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05855_ _00957_ _01276_ _01518_ _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08574_ _03607_ _03829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05786_ _01342_ _01451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_1_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07525_ _01896_ _03006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07456_ cpu.timer_div\[1\] _02933_ _02934_ cpu.timer_div\[5\] _02939_ _02940_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__06138__I _01797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06131__A1 _00979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06407_ _02063_ _02036_ _02064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07387_ _02854_ _02880_ _02881_ _00184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_118_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09126_ _03432_ _02857_ _04327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06338_ _01994_ _01995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08353__I _02944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_31_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07631__A1 _03088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09057_ _04257_ _04241_ _04259_ _04260_ _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06269_ _01925_ _01926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06434__A2 _02072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08008_ _02929_ _03395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08187__A2 _01842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09959_ _00218_ clknet_leaf_40_wb_clk_i cpu.spi.data_in_buff\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output46_I net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06757__B _02404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09439__A2 _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_70_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06122__A1 _01779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05887__I _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05079__I3 cpu.regs\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput70 net70 io_out[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06189__A1 _01335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08178__A2 _01417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput81 net81 io_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput92 net92 sram_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06189__B2 _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05936__A1 cpu.timer_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09678__A2 _00873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05127__I _00786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_qcpu_99 io_oeb[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_37_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05640_ _01097_ _01306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_86_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05571_ _01236_ _01237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_102_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_13_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07310_ cpu.regs\[5\]\[7\] _02815_ _02823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06113__A1 cpu.uart.divisor\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08290_ cpu.pwm_top\[3\] _03605_ _03609_ _03612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07241_ _01100_ _01105_ _01112_ _02777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_27_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07172_ _02719_ _02732_ _02737_ _00113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06123_ cpu.timer_capture\[14\] _01233_ _01782_ _01236_ _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__06416__A2 _02072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06054_ _01500_ _01714_ _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_113_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_115_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05005_ _00002_ _00702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07517__I net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09813_ _00009_ clknet_leaf_57_wb_clk_i cpu.instr_cycle\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09118__A1 _02271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06956_ _02556_ _02218_ _02571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09744_ _02574_ _04857_ _04858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09675_ _00827_ _01854_ _00913_ _04801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06887_ _02512_ _00053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05907_ _01436_ _00765_ _01569_ _01570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06027__S1 _00969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08626_ _03860_ _03875_ _00429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05838_ _01498_ _01499_ _01501_ _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05155__A2 cpu.ROM_spi_mode vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08557_ _03816_ _03817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05769_ _00610_ _01434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_91_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06104__A1 cpu.PORTB_DDR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07152__I0 _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07508_ _02954_ _02963_ _02957_ _02991_ _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_08488_ cpu.timer_capture\[13\] _03764_ _03758_ _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07439_ cpu.spi.dout\[6\] _02925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09109_ _04257_ _04302_ _04310_ _04260_ _04311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_17_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07604__A1 _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05918__A1 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06591__A1 _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_42_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_42_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_68_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08096__A1 _02856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer3 _00868_ net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_11_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05909__A1 net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07790_ _03210_ _03221_ _03222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06810_ cpu.uart.divisor\[2\] _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05224__I3 cpu.regs\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06741_ _00620_ _02390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09520__A1 _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09460_ cpu.ROM_spi_cycle\[2\] _04632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06672_ _01917_ _01919_ _02325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08168__I cpu.toggle_top\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08411_ _03702_ _03692_ _03656_ _03703_ _03704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09391_ _04575_ _00494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06885__A2 _02508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05623_ cpu.regs\[4\]\[7\] cpu.regs\[5\]\[7\] cpu.regs\[6\]\[7\] cpu.regs\[7\]\[7\]
+ _01285_ _01286_ _01289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_05554_ _00997_ _01062_ _01220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08342_ cpu.timer_top\[13\] _03644_ _03646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05485_ _01150_ _01151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08273_ _02478_ _03599_ _03600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07224_ _02710_ _02765_ _02767_ _00135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07021__B _02623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07155_ cpu.regs\[12\]\[5\] _02720_ _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09587__A1 _02536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07086_ _02682_ _00082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_112_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06106_ _01476_ _01764_ _01765_ _01766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06037_ net44 _01020_ _01698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07988_ _03371_ _03378_ _00288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05376__A2 _01041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06573__A1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_114_Right_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06939_ _02548_ _02555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09727_ _02574_ _04842_ _04843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09658_ _04596_ _04590_ _04785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08609_ _03370_ _03860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09589_ _02538_ _04718_ _04723_ _00544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_53_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09578__A1 _02527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10295_ _00553_ clknet_leaf_79_wb_clk_i cpu.C vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08553__A2 _03813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06996__I cpu.toggle_top\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08305__A2 _03621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06316__A1 _01942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08069__A1 _03439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05270_ cpu.regs\[0\]\[4\] cpu.multiplier.a\[4\] cpu.regs\[2\]\[4\] cpu.regs\[3\]\[4\]
+ _00834_ _00926_ _00939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_3_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09547__I _04695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08792__A2 _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08960_ _04165_ _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_110_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07911_ cpu.uart.receive_buff\[3\] _03313_ _03316_ cpu.uart.receive_buff\[2\] _03319_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08891_ _04098_ _04099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07842_ _03207_ _03264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05358__A2 _01007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09512_ _04664_ _04673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07773_ _03146_ cpu.uart.div_counter\[6\] _03201_ _03208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_04985_ _00621_ _00685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05315__I _00982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06724_ _02375_ _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08847__A3 _00981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06307__A1 _01963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09443_ _04594_ _04618_ _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06655_ _02307_ _02308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_108_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09374_ _04560_ _04548_ _04544_ _02295_ _04561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_87_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05606_ _01139_ _00657_ _01272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05530__A2 _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07530__I _03010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08325_ _03623_ _03634_ _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06586_ _02185_ _02240_ _02241_ _02242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05537_ _01202_ _01087_ _01203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_61_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05468_ _01133_ _01134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08256_ _03585_ _03587_ _00347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05294__A1 _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07207_ _01431_ _01163_ _02759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08187_ _03494_ _01842_ _03536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05399_ _00587_ _01065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07138_ _02713_ _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07069_ cpu.uart.receiving net15 _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_100_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05597__A2 _01034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10080_ _00339_ clknet_leaf_118_wb_clk_i cpu.toggle_ctr\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_87_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08299__A1 _02463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07346__I0 _02818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08471__A1 cpu.timer_capture\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10278_ _00536_ clknet_leaf_98_wb_clk_i cpu.PORTB_DDR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09723__A1 _00873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06537__A1 _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04974__I _00663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06440_ _02074_ _02095_ _02096_ _02097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06371_ _02010_ _02013_ _02027_ _02028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08110_ _03469_ _03404_ _03470_ _00318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_83_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09090_ _04176_ _04276_ _04292_ _04202_ _04293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_71_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05322_ cpu.br_rel_dest\[2\] _00988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08041_ _03417_ _03413_ _03419_ _00300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_71_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05253_ cpu.regs\[12\]\[3\] cpu.regs\[13\]\[3\] cpu.regs\[14\]\[3\] cpu.regs\[15\]\[3\]
+ _00889_ _00837_ _00923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_101_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05184_ cpu.base_address\[0\] _00856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09992_ _00251_ clknet_leaf_26_wb_clk_i cpu.uart.div_counter\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08943_ _04149_ _04150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08874_ _04069_ _04082_ _04083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07525__I _01896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07825_ _03151_ _03250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07756_ _03088_ _03194_ _00240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_04968_ _00667_ _00656_ _00668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06707_ _02359_ _02360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09426_ _04566_ _04561_ _04605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07687_ cpu.uart.div_counter\[1\] _03136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_04899_ cpu.br_rel_dest\[6\] _00602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_109_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07260__I _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06638_ _02283_ _01936_ _02291_ _02292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09357_ _02305_ _04546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06569_ _02203_ _02224_ _02225_ _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09288_ _02337_ _02396_ _04483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08308_ _02936_ cpu.timer_div_counter\[1\] _03624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_34_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08239_ _03562_ _03575_ _03576_ _00341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_105_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08091__I _03456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10201_ _00459_ clknet_leaf_67_wb_clk_i cpu.last_addr\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__06216__B1 cpu.spi.divisor\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05114__S1 _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10132_ _00391_ clknet_leaf_5_wb_clk_i cpu.timer\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09705__A1 _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10063_ _00322_ clknet_leaf_2_wb_clk_i cpu.toggle_top\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_89_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08692__A1 _02556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09097__I _04169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06758__A1 _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05430__A1 _00618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05940_ cpu.toggle_top\[3\] _01418_ _01172_ _01603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05871_ _00741_ _01534_ _01535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07183__A1 _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07610_ _03074_ _03075_ _02930_ _00213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08590_ _03841_ _03842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07541_ cpu.spi.data_out_buff\[1\] _03016_ _02675_ _03020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07080__I _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07472_ cpu.timer_top\[8\] _02956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09211_ _03466_ _04408_ _04409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_63_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05497__A1 _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06423_ _02056_ _02078_ _02080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05041__S0 _00716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09950__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09142_ _03848_ _04328_ _04343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06354_ _01997_ _02000_ _02011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_16_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05305_ cpu.regs\[8\]\[5\] cpu.regs\[9\]\[5\] cpu.regs\[10\]\[5\] cpu.regs\[11\]\[5\]
+ _00898_ _00899_ _00973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_114_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09073_ _04275_ _04276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_21_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06285_ _01941_ _01942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_31_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08024_ _03399_ _03407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05236_ _00878_ _00886_ _00906_ _00907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_116_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05167_ _00838_ _00839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_12_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09975_ _00234_ clknet_leaf_39_wb_clk_i cpu.spi.counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05098_ _00759_ _00790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08926_ _03438_ _03433_ _03442_ _04133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07255__I _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09163__A2 _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08857_ _03836_ _04066_ _04067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07808_ _03176_ _03236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08910__A2 _03848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08788_ _00686_ _04001_ _04002_ _00464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06921__A1 cpu.timer_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07739_ _03180_ _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_60_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09409_ _04549_ _04543_ _01037_ _01038_ _04590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_109_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_67_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_67_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_63_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08729__A2 cpu.regs\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05099__S0 _00770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10115_ _00374_ clknet_leaf_11_wb_clk_i cpu.timer_top\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10046_ _00305_ clknet_leaf_53_wb_clk_i cpu.orig_flags\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08665__A1 _02385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05479__A1 _00654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05023__S0 _00697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06140__A2 _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07640__A2 _03094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_1 _03908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06070_ _01730_ _01731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_111_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05021_ _00704_ _00717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_111_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_105_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06972_ _02585_ _02569_ _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09760_ _00023_ clknet_leaf_94_wb_clk_i cpu.regs\[2\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05923_ _00615_ _01585_ _01586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09691_ _04788_ _04815_ _04816_ _00628_ _04817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08711_ _03942_ cpu.regs\[3\]\[0\] _03943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_83_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08499__A4 _00999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08642_ cpu.IO_addr_buff\[5\] _03858_ _03888_ _03883_ _03889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_89_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05854_ _01281_ _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xrebuffer13 _00870_ net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08573_ _03798_ _03826_ _03828_ _00423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06847__C _02478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05785_ _01449_ _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07524_ _00694_ _02907_ _03005_ _00197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_65_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07455_ cpu.timer_div\[5\] _02934_ cpu.timer_div_counter\[7\] _02935_ _02938_ _02939_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06406_ _02032_ _02063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05190__I0 cpu.regs\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07386_ _00715_ _02869_ _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_118_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09125_ _04325_ _04273_ _04326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06337_ _01954_ _01956_ _01994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_114_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09056_ _04152_ _04260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06268_ _00983_ _01312_ _00663_ _01924_ _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_0_114_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08007_ _03393_ cpu.uart.receive_div_counter\[14\] _03346_ _03385_ _03394_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__05642__A1 _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05219_ _00889_ _00890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06199_ _00826_ _01854_ _01857_ _01858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_12_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09958_ _00217_ clknet_leaf_40_wb_clk_i cpu.spi.data_in_buff\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_90_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08909_ _03847_ _04098_ _04117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_114_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_114_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09889_ _00148_ clknet_leaf_90_wb_clk_i cpu.regs\[7\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07713__I _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05253__S0 _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output39_I net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06773__B _02406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09375__I _02359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06999__I _02610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput60 net60 io_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07386__A1 _00715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput71 net71 io_out[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput82 net82 io_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput93 net93 sram_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_37_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10029_ _00288_ clknet_leaf_29_wb_clk_i cpu.uart.receive_div_counter\[11\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08719__I _03908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06239__I _01896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05570_ _01235_ _01236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_102_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07240_ _01351_ _02776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07171_ cpu.regs\[11\]\[2\] _02736_ _02737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06122_ _01779_ _01780_ _01781_ _01782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08810__A1 _00905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06053_ cpu.timer_capture\[13\] _01233_ _01714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05004_ _00699_ _00700_ _00002_ _00701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09812_ _00008_ clknet_leaf_57_wb_clk_i net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_6_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07019__B _02623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05318__I _00873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06955_ cpu.PC\[5\] _02570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09743_ _02218_ _04856_ _04857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07533__I _03010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09234__B _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09674_ _00827_ _01854_ _01857_ _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06886_ cpu.timer_capture\[6\] _02494_ _02511_ _02506_ _02512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05906_ _01315_ _01562_ _01564_ _01568_ _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_68_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08625_ _00590_ _03861_ _03874_ _03870_ _03875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05837_ cpu.timer_capture\[10\] _01228_ _01500_ _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08556_ _01210_ _02609_ _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_77_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05768_ _01430_ _01431_ _01432_ _01433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07507_ cpu.timer_top\[10\] _02989_ _02990_ cpu.timer_top\[9\] _02991_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_92_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05699_ _01363_ _01364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07152__I1 cpu.regs\[12\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08487_ cpu.timer\[13\] _03761_ _03766_ _03767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07438_ _02923_ _02924_ _02915_ _00192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_92_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07369_ _02862_ _02863_ _02864_ _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_9_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09108_ _02596_ _04190_ _04310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08801__A1 _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09039_ _04009_ _04243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_99_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_82_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_82_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_31_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_11_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_11_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_82_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer4 _00896_ net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05606__A1 _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08020__A2 _03404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06740_ _00679_ _02389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06671_ cpu.mem_cycle\[5\] _01910_ _02324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_64_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05622_ _01284_ _01287_ _01288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06334__A2 _01990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08410_ _03702_ _03698_ _03703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09390_ _04573_ _04574_ _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_47_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05553_ _01174_ _01217_ _01218_ _01219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_59_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08341_ _02453_ _03643_ _03645_ _03641_ _00374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_74_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05484_ _01149_ _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_46_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08272_ cpu.pwm_counter\[6\] _03597_ _03599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09036__A1 _04070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05601__I _01115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07223_ cpu.regs\[8\]\[0\] _02766_ _02767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07154_ _01751_ _02725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07085_ _02677_ _02681_ _02682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06105_ net66 _01197_ _01765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06036_ net56 cpu.PORTA_DDR\[5\] _01192_ _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_66_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06270__A1 _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08011__A2 _03396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07987_ _03376_ _03366_ _03346_ _03377_ _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06573__A2 _02229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06938_ _02553_ _02554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09726_ _02236_ _04839_ _04841_ _02578_ _04842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_69_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09657_ _04742_ _02335_ _04783_ _04784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_69_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06869_ _02470_ _02497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_96_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08608_ _03585_ _03859_ _00427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09588_ cpu.PORTA_DDR\[6\] _04719_ _04720_ _04723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08539_ cpu.timer_div\[5\] _03799_ _03802_ _03803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08094__I _03403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10294_ _00552_ clknet_leaf_61_wb_clk_i net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08978__B _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_88_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06010__C _01434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05827__A1 _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07910_ _03243_ _03318_ _00270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08890_ _03437_ _04069_ _04098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07841_ _03248_ cpu.uart.counter\[1\] _03252_ cpu.uart.counter\[3\] _03263_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__07284__S _02796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09741__A2 _04854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07772_ _03176_ _03207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09511_ _04664_ _04672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_04984_ _00644_ _00676_ _00683_ _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06723_ net1 _02374_ _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06654_ cpu.startup_cycle\[3\] cpu.startup_cycle\[2\] _02307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09442_ cpu.ROM_spi_dat_out\[4\] _04562_ _04612_ _04618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_108_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08847__A4 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09373_ cpu.startup_cycle\[2\] _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_93_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09257__A1 _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05605_ _01036_ _01270_ _01271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_19_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06585_ _02239_ _02197_ _02241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05536_ _01016_ _01202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08324_ cpu.timer_div_counter\[7\] _03633_ _03634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_47_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05467_ _00998_ _01125_ _01133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08255_ _03584_ _03586_ _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05398_ _00585_ _01064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05294__A2 _00950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07206_ _02742_ _02747_ _02758_ _00126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08186_ _03527_ _03529_ _03534_ _03535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_104_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07137_ _02712_ _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_18_Left_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07068_ cpu.uart.receive_counter\[0\] _02667_ _02668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__06794__A2 _02433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06019_ _01680_ _00017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09496__A1 net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09709_ _01752_ _04821_ _04828_ _00559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_27_Left_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08299__A2 _03613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07346__I1 cpu.regs\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05809__A1 net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05241__I _00910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08552__I _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_36_Left_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_103_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10277_ _00535_ clknet_leaf_13_wb_clk_i cpu.PORTB_DDR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06800__I _02390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09723__A2 _01971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07734__A1 _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_45_Left_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_4_0_0_wb_clk_i clknet_0_wb_clk_i clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_75_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06370_ _02020_ _02026_ _02011_ _02027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__05151__I cpu.PORTA_DDR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05321_ _00987_ net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08040_ cpu.orig_IO_addr_buff\[6\] _03418_ _03411_ _03419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05252_ _00913_ _00919_ _00921_ _00922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09558__I _04695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_54_Left_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_11_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09411__A1 _02366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05183_ _00829_ _00854_ _00855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_24_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09991_ _00250_ clknet_leaf_26_wb_clk_i cpu.uart.div_counter\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08942_ _01162_ _04149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06710__I _00691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09714__A2 _02425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08873_ _01116_ _04081_ _04082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_63_Left_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07824_ _00599_ _01895_ _03249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07755_ cpu.uart.div_counter\[3\] _03178_ _03182_ _03193_ _03194_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_04967_ _00654_ _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06706_ _01000_ _02359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07686_ _03133_ cpu.uart.divisor\[5\] _02448_ _03134_ _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09425_ _04595_ _04602_ _04604_ _00499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_04898_ _00600_ _00601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_50_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06637_ _02259_ _02290_ _02291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09356_ _04544_ _04545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06568_ _02205_ _02223_ _02225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09287_ _04480_ _04482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05519_ _01024_ _01184_ _01185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_72_Left_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08307_ cpu.timer_div_counter\[0\] _03623_ _00362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06499_ _02137_ _02143_ _02156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_35_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08238_ cpu.toggle_ctr\[11\] _03497_ _03573_ _03576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_62_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10200_ _00458_ clknet_leaf_67_wb_clk_i cpu.last_addr\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_08169_ cpu.toggle_top\[3\] _03518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_101_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10131_ _00390_ clknet_leaf_2_wb_clk_i cpu.timer\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output69_I net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08321__B _03621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10062_ _00321_ clknet_leaf_2_wb_clk_i cpu.toggle_clkdiv vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09469__A1 _04558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06207__A1 _01852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05870_ _00879_ _01533_ _01534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_89_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__04985__I _00621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07540_ cpu.spi.data_out_buff\[2\] _03007_ _03018_ _03019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07471_ cpu.timer_top\[9\] _02955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_118_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09210_ _03463_ _04381_ _04408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__05497__A2 _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06422_ _02056_ _02078_ _02079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__05041__S1 _00731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09141_ _04152_ _04342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06353_ _00872_ _02002_ _02009_ _02010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_17_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09072_ _02213_ _04240_ _04275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_16_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05304_ _00967_ _00971_ _00972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08023_ _00995_ _03402_ _03406_ _00295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06284_ _01940_ _01941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_31_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05235_ _00905_ _00906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_4_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05166_ _00837_ _00838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_116_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09974_ _00233_ clknet_leaf_39_wb_clk_i cpu.spi.counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07536__I _03010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05097_ _00787_ _00788_ _00756_ _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08925_ _04131_ _03436_ cpu.PC\[0\] _04132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__05272__I2 cpu.regs\[10\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input20_I io_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08856_ _04008_ _04064_ _04065_ _04035_ _04066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05056__I _00731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07807_ _03233_ _03235_ _00250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08787_ cpu.ROM_addr_buff\[11\] _03988_ _04002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05999_ _01325_ _00948_ _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_84_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07738_ _03154_ _03155_ _03150_ _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08123__A1 _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07669_ _02651_ cpu.uart.div_counter\[15\] _03117_ cpu.uart.divisor\[3\] _03118_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__08674__A2 _00715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09408_ _04587_ _04588_ _01037_ _04589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_109_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09339_ _01917_ _04531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_109_Right_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07937__A1 _02677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05099__S1 _00786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_36_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_36_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10114_ _00373_ clknet_leaf_3_wb_clk_i cpu.timer_top\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10045_ _00304_ clknet_leaf_53_wb_clk_i cpu.orig_flags\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_59_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07181__I _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05023__S1 _00698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05020_ _00703_ _00716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_22_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07356__I _02851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06971_ _02213_ _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05922_ cpu.uart.divisor\[11\] _01380_ _01585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09690_ _01303_ _04788_ _04816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08710_ _03908_ _03942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08641_ _03838_ _03886_ _03887_ _03888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05853_ _01261_ _01511_ _01513_ _01516_ _00884_ _01517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__09571__I _04710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer14 _02090_ net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_107_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08572_ _02648_ _03827_ _03821_ _03828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05784_ _00888_ _01446_ _01448_ _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_07523_ _02364_ cpu.spi.busy _03005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_65_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07454_ cpu.timer_div\[0\] _02936_ cpu.timer_div_counter\[2\] _01496_ _02937_ _02938_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06405_ net115 _02061_ _02062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_45_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07385_ _01466_ _02234_ _02879_ _02880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_118_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09124_ cpu.PC\[8\] _04325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_17_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06336_ _01992_ _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09055_ _02570_ _04258_ _04259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06267_ _01336_ _01434_ _01924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08006_ cpu.uart.receive_div_counter\[15\] _03393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_102_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05218_ _00004_ _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06198_ _01855_ _01806_ _01856_ _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_13_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05149_ cpu.PORTA_DDR\[0\] net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_09957_ _00216_ clknet_leaf_41_wb_clk_i cpu.spi.data_in_buff\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_90_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08908_ _04115_ _04116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09888_ _00147_ clknet_leaf_109_wb_clk_i cpu.regs\[7\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08344__A1 cpu.timer_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08839_ _01033_ _01101_ _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_56_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05253__S1 _00837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput61 net61 io_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput50 net50 io_oeb[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput72 net72 io_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput94 net94 sram_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput83 net83 sram_addr[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10028_ _00287_ clknet_leaf_31_wb_clk_i cpu.uart.receive_div_counter\[10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08335__A1 _02527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07170_ _02730_ _02736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06121_ cpu.timer_capture\[6\] _01401_ _01226_ _01781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06052_ _01710_ _01711_ _01712_ _01713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05003_ cpu.regs\[4\]\[0\] cpu.regs\[5\]\[0\] cpu.regs\[6\]\[0\] cpu.regs\[7\]\[0\]
+ _00697_ _00698_ _00700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_113_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09811_ _00074_ clknet_leaf_116_wb_clk_i cpu.toggle_top\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09742_ _03442_ _03438_ _03446_ _04856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07814__I _02929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06954_ _02219_ _02569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08326__A1 _01240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09673_ _01266_ _04008_ _04798_ _04799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05905_ _01457_ _01565_ _01567_ _01568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06885_ _02496_ _02508_ _02497_ _02510_ _02511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_68_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08624_ _03862_ _03872_ _03873_ _03874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05836_ _01032_ _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08555_ _02426_ _03815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05767_ _01097_ _01432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_77_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07506_ cpu.timer\[9\] _02990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05698_ _01019_ _01120_ _01363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_49_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08486_ _02503_ _03751_ _03766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07437_ cpu.spi.data_in_buff\[5\] _02908_ _02924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_4_13_0_wb_clk_i clknet_0_wb_clk_i clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_9_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07368_ _02862_ _02863_ _02573_ _02864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_33_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09107_ _04179_ _04302_ _04308_ _04186_ _04309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_60_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06319_ _00841_ _00846_ _00850_ _00852_ _01957_ _01976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_33_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08801__A2 _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06812__A1 _02447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07299_ _02785_ _02811_ _02816_ _00161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09038_ _04241_ _04242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08380__I _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05379__A1 _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output51_I net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07540__A2 _03007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05551__A1 cpu.spi.dout\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08555__I _02426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer5 _02053_ net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_51_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_51_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_11_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05606__A2 _00657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05790__A1 _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06670_ _02321_ _01920_ _02322_ _02323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_59_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05621_ cpu.regs\[0\]\[7\] cpu.multiplier.a\[7\] cpu.regs\[2\]\[7\] cpu.regs\[3\]\[7\]
+ _01285_ _01286_ _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_86_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05542__A1 _01065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__04993__I _00691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05552_ _00589_ _01063_ _01129_ _01218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_58_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08340_ cpu.timer_top\[12\] _03644_ _03645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05483_ cpu.br_rel_dest\[1\] _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_58_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08271_ cpu.pwm_counter\[6\] _03597_ _03598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07222_ _02764_ _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09036__A2 _02569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07153_ _02724_ _00107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06104_ cpu.PORTB_DDR\[6\] _01202_ _01239_ _01363_ _01762_ _01763_ _01764_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
X_07084_ _02678_ _02680_ _02681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_2_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06035_ _01128_ _01184_ _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08547__A1 _00650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07986_ _03376_ _03372_ _03377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06937_ _02547_ _02553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09725_ _04043_ _01970_ _04840_ _04841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09656_ _04729_ _04781_ _04782_ _04783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_69_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08607_ _03836_ _03853_ _03858_ _01065_ _03859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06868_ _02472_ _02496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_96_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05819_ cpu.uart.divisor\[2\] _01377_ _01483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06799_ _02427_ _02436_ _02438_ _00039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09587_ _02536_ _04718_ _04722_ _00543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08538_ _03757_ _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_64_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08469_ _00906_ _03751_ _03752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07589__A2 _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10293_ _00551_ clknet_leaf_59_wb_clk_i net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05239__I _00908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09266__A2 _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08285__I _03608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07403__B _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06324__I0 _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05827__A2 _00999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08777__A1 cpu.ROM_addr_buff\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05149__I cpu.PORTA_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07840_ _03158_ _03262_ _00256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07771_ _03205_ _03206_ _00243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09510_ _03796_ _04665_ _04671_ _00517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_04983_ _00677_ _00682_ _00683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06722_ _00579_ _02374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08701__A1 _03453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09441_ _04595_ _04616_ _04617_ _00502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_40_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06653_ _02305_ _02299_ _02306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_65_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09372_ _04558_ _04559_ _00491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05604_ _01035_ _01270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06584_ _02239_ _02197_ _02240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05535_ _01194_ _01196_ _01200_ _01201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08323_ cpu.timer_div_counter\[6\] _03630_ _03633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05612__I _00884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05466_ _01082_ _01126_ _01130_ _01131_ _01132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_08254_ cpu.pwm_counter\[1\] _03586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05397_ _01062_ _01063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07205_ cpu.regs\[10\]\[7\] _02750_ _02758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08185_ _03531_ _03533_ _03534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07136_ _01114_ _02711_ _02712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07067_ cpu.uart.receiving _02666_ _02667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_76_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05059__I _00717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06018_ _01679_ cpu.regs\[15\]\[4\] _01167_ _01680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05349__A4 _01006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07969_ _02650_ _03360_ _03363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09708_ cpu.regs\[9\]\[5\] _04824_ _04828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05754__A1 _01417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09639_ _02339_ _02396_ _04767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_41_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08833__I _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_70_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10276_ _00534_ clknet_leaf_14_wb_clk_i cpu.PORTB_DDR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07734__A2 _01895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07498__A1 cpu.timer_top\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05320_ _00984_ _00986_ _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_61_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05251_ _00920_ _00921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_101_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05182_ _00853_ _00854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07359__I _02851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_7_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06225__A2 cpu.spi.divisor\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09990_ _00249_ clknet_leaf_25_wb_clk_i cpu.uart.div_counter\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08941_ _04138_ _04145_ _04146_ _04147_ _04148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08872_ _01327_ _04080_ _04081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08922__A1 _03057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07823_ cpu.uart.counter\[0\] _03248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_71_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07754_ _03117_ _03191_ _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_04966_ _00665_ _00666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06705_ _02320_ _02354_ _02357_ _02358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07685_ cpu.uart.div_counter\[2\] _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07489__A1 cpu.timer_top\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09424_ cpu.ROM_spi_dat_out\[1\] _04598_ _04603_ _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_04897_ cpu.br_rel_dest\[5\] _00600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06636_ net20 _02229_ _02287_ _02289_ _02290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06161__A1 net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09355_ _04543_ _04544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_90_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06567_ _02205_ _02223_ _02224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09286_ _04480_ _04481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08989__A1 _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05518_ _00587_ _01075_ _01184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08306_ _03622_ _03623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06498_ _02137_ _02143_ _02155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05449_ _01036_ _01115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08237_ _03497_ _03573_ cpu.toggle_ctr\[11\] _03575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_105_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07269__I _02796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08168_ cpu.toggle_top\[4\] _03517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_108_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_108_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_42_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08099_ _03461_ _03459_ _03462_ _00315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06216__A2 cpu.spi.divisor\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07119_ cpu.regs\[13\]\[1\] _02700_ _02702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05975__A1 _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10130_ _00389_ clknet_leaf_1_wb_clk_i cpu.timer\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10061_ _00320_ clknet_leaf_58_wb_clk_i cpu.had_int vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08321__C _02404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05517__I cpu.uart.divisor\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05027__I0 cpu.regs\[12\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09152__C _04321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09157__B2 _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10259_ _00517_ clknet_leaf_46_wb_clk_i net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05427__I _00583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Left_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05718__A1 cpu.uart.divisor\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05194__A2 _00865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07470_ cpu.timer_top\[12\] _02952_ _02953_ cpu.timer_top\[11\] _02954_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06421_ _02062_ _02075_ _02077_ _02078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_09140_ _04340_ _04328_ _04254_ _04341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_6_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_6_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_8_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06352_ _00783_ _02009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09071_ _02585_ _04273_ _04274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06283_ _00745_ _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_05303_ _00842_ _00970_ _00845_ _00971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_44_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08022_ cpu.orig_IO_addr_buff\[1\] _03404_ _03303_ _03406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05234_ _00904_ _00905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05165_ _00005_ _00837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_116_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09973_ _00232_ clknet_leaf_34_wb_clk_i cpu.spi.counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06721__I _02372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05096_ cpu.regs\[4\]\[5\] cpu.regs\[5\]\[5\] cpu.regs\[6\]\[5\] cpu.regs\[7\]\[5\]
+ _00785_ _00786_ _00788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_40_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08924_ cpu.PC\[2\] _04131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05272__I3 cpu.regs\[11\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08855_ _03425_ _04008_ _04065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08786_ cpu.last_addr\[11\] _03996_ _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07806_ _03230_ _03231_ _03234_ _03235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input13_I io_in[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07737_ _03137_ _03178_ _03179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05998_ _00764_ _01558_ _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_04949_ _00648_ _00649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_84_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07668_ cpu.uart.div_counter\[3\] _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__06134__A1 _01733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09407_ _01038_ _02308_ _04563_ _02309_ _04588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_07599_ _03065_ _03045_ _03066_ _03002_ _03067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_23_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06619_ _02267_ _02273_ _02274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_118_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09338_ _03588_ _04529_ _04530_ _00486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_51_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09269_ _04463_ _04442_ _04464_ _04465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output81_I net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10113_ _00372_ clknet_leaf_11_wb_clk_i cpu.timer_top\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05247__I _00916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_76_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_76_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10044_ _00303_ clknet_leaf_52_wb_clk_i cpu.orig_flags\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_59_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08558__I _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06125__A1 cpu.timer_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09378__A1 _03057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05157__I cpu.base_address\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06970_ _02548_ _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input5_I io_in[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05921_ _01583_ _01377_ _01381_ _01584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09550__A1 cpu.PORTB_DDR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08640_ _02419_ _03851_ _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05852_ _01515_ _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xrebuffer15 _00576_ net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_89_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08571_ _03816_ _03827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_88_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05783_ _00897_ _01447_ _01448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07522_ _03000_ _03003_ _03004_ _00196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06116__A1 cpu.uart.dout\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07453_ cpu.timer_div\[0\] _02936_ _02933_ cpu.timer_div\[1\] _02937_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_64_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06404_ _01968_ _02059_ _02060_ _02061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09123_ _04298_ _04323_ _04324_ _00477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07384_ _02871_ _02878_ _01931_ _02879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_118_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06335_ _00744_ _01955_ _01991_ _01992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06266_ _01906_ _01922_ _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_89_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09054_ _04149_ _04258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08005_ cpu.uart.receive_div_counter\[15\] _03389_ _03392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05217_ _00887_ _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07547__I _02455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06197_ _00810_ _01801_ _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05148_ cpu.PORTA_DDR\[7\] net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_110_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09956_ _00215_ clknet_leaf_41_wb_clk_i cpu.spi.data_in_buff\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05079_ cpu.regs\[0\]\[4\] _00768_ _00769_ cpu.regs\[3\]\[4\] _00770_ _00771_ _00772_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_90_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08907_ _00671_ _00681_ _04115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09887_ _00146_ clknet_leaf_87_wb_clk_i cpu.regs\[7\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09541__A1 _03801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08838_ _04041_ _04044_ _04047_ _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_99_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08769_ _03936_ _03988_ _03989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06107__A1 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07607__A1 _03043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08062__B _03430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput51 net51 io_oeb[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput40 net40 io_oeb[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput62 net62 io_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput73 net73 io_out[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput84 net84 sram_addr[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput95 net95 sram_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_37_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10027_ _00286_ clknet_leaf_31_wb_clk_i cpu.uart.receive_div_counter\[9\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09532__A1 _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_90_Left_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08099__A1 _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06120_ cpu.timer_div\[6\] _01397_ _01221_ _01780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06051_ cpu.timer_capture\[5\] _01402_ _01227_ _01712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05002_ cpu.regs\[0\]\[0\] cpu.multiplier.a\[0\] _00696_ cpu.regs\[3\]\[0\] _00697_
+ _00698_ _00699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_41_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_113_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_99_Right_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09810_ _00073_ clknet_leaf_116_wb_clk_i cpu.toggle_top\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09582__I _04710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06953_ _02552_ _02566_ _02568_ _00063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09741_ _02237_ _04854_ _02600_ _04855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05904_ _01543_ _01566_ _01567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08326__A2 _02433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09672_ _04794_ _04797_ _03837_ _04798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06884_ _02509_ _02499_ _02510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_68_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08623_ _01525_ _03867_ _03873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05835_ cpu.timer_capture\[2\] _01223_ _01234_ _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08554_ _00617_ _03813_ _03814_ _00418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05766_ _01304_ _01431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05560__A2 _01225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07505_ cpu.timer\[10\] _02989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05697_ _01360_ _01361_ _01190_ _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08485_ _03760_ _03763_ _03765_ _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07436_ cpu.spi.dout\[5\] _02916_ _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07367_ _02098_ _02101_ _02863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_45_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08661__I _03829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09106_ _04305_ _04306_ _04307_ _04308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06318_ _00861_ net125 _00868_ _00866_ _01974_ _01975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_32_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09037_ _02570_ _04239_ _04240_ _04241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_60_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07298_ cpu.regs\[5\]\[2\] _02815_ _02816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06249_ _01003_ _01906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_4_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06576__A1 _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09939_ _00198_ clknet_leaf_18_wb_clk_i cpu.spi.data_out_buff\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output44_I net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08057__B _03430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07056__A2 cpu.uart.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08571__I _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer6 _02036_ net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_91_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_91_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06091__I _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08556__A2 _02609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06567__A1 _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_20_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_20_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09505__A1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05435__I _01034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_30_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05620_ _00838_ _01286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07650__I _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_47_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05551_ cpu.spi.dout\[0\] _01177_ _01182_ _01216_ _01217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05482_ _01147_ _01148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07295__A2 _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05170__I _00006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08270_ _03588_ _03596_ _03597_ _00351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08492__A1 cpu.timer_capture\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07221_ _02764_ _02765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07047__A2 _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07152_ _01679_ cpu.regs\[12\]\[4\] _02713_ _02724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06103_ net57 _00596_ _01358_ _01127_ _01763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_07083_ _02679_ _02669_ _02680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06034_ cpu.uart.divisor\[5\] _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_2_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08547__A2 _01115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07985_ cpu.uart.receive_div_counter\[11\] _03376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06936_ _02551_ _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09724_ _04043_ _00985_ _01970_ _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09655_ _02308_ _04551_ _04757_ _04782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06867_ _01694_ _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05818_ _01480_ _01481_ _01186_ _01482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08606_ _03857_ _03858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08180__B1 cpu.toggle_top\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06798_ cpu.uart.divisor\[0\] _02437_ _02391_ _02438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08656__I _03899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06730__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09586_ cpu.PORTA_DDR\[5\] _04719_ _04720_ _04722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08537_ _02459_ _03801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05749_ _01409_ _01412_ _01413_ _01414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08468_ _03741_ _03751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07419_ _01901_ _02910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_80_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05013__C _00003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08399_ _02509_ _03693_ _03694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08786__A2 _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10292_ _00550_ clknet_leaf_59_wb_clk_i net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_114_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05080__S0 _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09726__A1 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07770_ _03145_ _03201_ _00645_ _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_04982_ _00680_ _00681_ _00643_ _00682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_75_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06721_ _02372_ _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05763__A2 _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06960__A1 _02569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09440_ cpu.ROM_spi_dat_out\[4\] _04598_ _04603_ _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06652_ cpu.startup_cycle\[6\] _02305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_91_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08476__I _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09371_ _04549_ _04554_ _04559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05603_ _01257_ _01262_ _01265_ _01268_ _01269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06583_ _02189_ _02239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05534_ net59 _01198_ _01199_ _01200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08322_ cpu.timer_div_counter\[6\] _03630_ _03632_ _00368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08253_ _03370_ _03585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05465_ _01085_ _01088_ _01129_ _01131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07204_ _02757_ _00125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05396_ _01048_ _00597_ _01062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_61_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08184_ _03522_ _03532_ cpu.toggle_top\[0\] _03528_ _03533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06228__B1 cpu.spi.divisor\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07135_ _01148_ _01154_ _02544_ _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_07066_ _02637_ _02647_ _02665_ _02666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_76_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06017_ _01678_ _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_100_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07968_ _03359_ _03356_ _03362_ _03310_ _00284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09707_ _04827_ _00558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06919_ _02536_ _02533_ _02537_ _02531_ _00060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07899_ _03055_ _03310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_87_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09638_ _02326_ _04765_ _02329_ _02340_ _04766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__05803__I _01467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09569_ _01395_ _01071_ _04663_ _04710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_38_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07893__C _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10275_ _00533_ clknet_leaf_49_wb_clk_i cpu.PORTB_DDR\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05993__A2 _01304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09613__C _02439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06170__A2 _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08447__A1 cpu.timer_capture\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05250_ _00912_ _00918_ _00886_ _00920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05681__A1 _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05181_ _00841_ _00846_ _00850_ _00852_ _00853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_4_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08940_ _00608_ _01161_ _04147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08871_ _01303_ _00935_ _04079_ _04080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_07822_ _03094_ _03247_ _03242_ _00253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_71_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06933__A1 _02203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07753_ _03134_ _03189_ _03192_ _03113_ _00239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_04965_ _00664_ _00612_ _00665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06704_ cpu.ROM_addr_buff\[3\] _02355_ _02356_ cpu.ROM_addr_buff\[7\] _02327_ _02357_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_07684_ cpu.uart.div_counter\[5\] _03133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_04896_ _00589_ _00598_ _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09423_ _03829_ _04603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06635_ _01927_ _02288_ _02289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09354_ cpu.startup_cycle\[0\] _04543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06161__A2 _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06566_ _02207_ _02208_ _02222_ _02223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_08305_ _02390_ _03621_ _03622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09285_ _04478_ _04479_ _04480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05517_ cpu.uart.divisor\[0\] _01183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_90_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06497_ _02128_ _02152_ _02153_ _02154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08236_ _03563_ _03574_ _00340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05448_ _01113_ _01114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08167_ _03514_ cpu.toggle_top\[5\] cpu.toggle_top\[4\] _03515_ _03516_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05379_ _01023_ _01032_ _01035_ _01044_ _01045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_07118_ _01353_ _02699_ _02701_ _00095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08098_ cpu.orig_PC\[9\] _03454_ _03457_ _03462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05424__A1 _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07049_ _02648_ _02649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_10060_ _00319_ clknet_leaf_70_wb_clk_i cpu.orig_PC\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10258_ _00516_ clknet_leaf_45_wb_clk_i net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__08904__A2 _01151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10189_ _00447_ clknet_leaf_69_wb_clk_i cpu.ROM_addr_buff\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_89_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06143__A2 _01691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06420_ _00814_ _02041_ _02076_ _02077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_29_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07340__A1 _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06351_ _01989_ _02005_ _02007_ _02008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_112_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09070_ _04072_ _04273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05302_ cpu.regs\[4\]\[5\] cpu.regs\[5\]\[5\] cpu.regs\[6\]\[5\] cpu.regs\[7\]\[5\]
+ _00968_ _00969_ _00970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_16_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06282_ _01938_ _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08021_ _01076_ _03402_ _03405_ _00294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05233_ _00888_ net118 _00903_ _00904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05164_ _00835_ _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_116_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09972_ _00231_ clknet_leaf_34_wb_clk_i cpu.spi.counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05095_ cpu.regs\[0\]\[5\] _00783_ _00784_ cpu.regs\[3\]\[5\] _00785_ _00786_ _00787_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_40_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08923_ _04130_ _00471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_110_Left_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08854_ _04056_ _04060_ _04063_ _04055_ _04064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08785_ _03999_ _03970_ _04000_ _03993_ _00463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07805_ _02390_ _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05997_ _00780_ _01659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_04948_ _00647_ _00648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07736_ _03177_ _03178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08659__A1 _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_04879_ net71 _00581_ _00582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07667_ _02649_ _03115_ cpu.uart.div_counter\[8\] _02642_ _03116_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_09406_ _02312_ _04585_ _04586_ _04570_ _04587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_07598_ _03065_ _03062_ _03066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_23_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06618_ _02268_ _02270_ _02272_ _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09337_ _02338_ _01916_ _04480_ _04530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06549_ cpu.PC\[11\] _02206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_51_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09268_ _02204_ _01537_ _04464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08219_ _03562_ _03563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09199_ _00913_ _04256_ _04397_ _04262_ _04398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_15_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09387__A2 _04571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08332__C _02542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output74_I net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10112_ _00371_ clknet_leaf_3_wb_clk_i cpu.timer_top\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10043_ _00302_ clknet_leaf_52_wb_clk_i cpu.orig_flags\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_59_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05263__I _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05008__S0 _00703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_45_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_45_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08574__I _03607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09075__A1 cpu.PC\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05884__A1 net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06061__A1 cpu.toggle_top\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05920_ cpu.uart.divisor\[3\] _01583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_05851_ _01272_ _01514_ _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xrebuffer16 net129 net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_89_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08570_ _03816_ _03826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_83_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06269__I _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07521_ cpu.spi.data_out_buff\[7\] _02911_ _03003_ _03004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05782_ _00847_ _00851_ _01284_ _01447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05173__I _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09302__A2 cpu.ROM_addr_buff\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07452_ cpu.timer_div_counter\[0\] _02936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05175__I0 cpu.regs\[12\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__04945__C _00645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09066__A1 _02186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05875__A1 _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06403_ _01951_ _01691_ _02059_ _02033_ _02060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07383_ _02852_ _02877_ _02878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09122_ _00693_ _04324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06334_ _01943_ _01990_ _00744_ _01991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_45_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06265_ _01907_ _01921_ _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09053_ _04150_ _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08004_ _03390_ _03391_ _03242_ _00291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06196_ _00810_ _01801_ _01855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05216_ _00848_ _00887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05147_ cpu.PORTB_DDR\[7\] net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_40_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06052__A1 _01710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09955_ _00214_ clknet_leaf_41_wb_clk_i cpu.spi.data_in_buff\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05078_ _00753_ _00771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_90_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08906_ _04110_ _04112_ _04113_ _04114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09886_ _00145_ clknet_leaf_88_wb_clk_i cpu.regs\[7\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08837_ _01169_ _04045_ _04046_ _04047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07552__A1 _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08768_ _03969_ _03988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07719_ _03009_ cpu.spi.counter\[1\] _03165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08699_ _03916_ _03933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_0_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_0_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08804__A1 _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06043__A1 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput52 net52 io_oeb[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput41 net41 io_oeb[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput74 net74 io_out[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput63 net63 io_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput85 net85 sram_addr[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_8_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput96 net96 sram_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06798__B _02391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10026_ _00285_ clknet_leaf_31_wb_clk_i cpu.uart.receive_div_counter\[8\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05229__S0 _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_20_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06817__I _01694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09048__A1 _02214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06050_ cpu.timer_div\[5\] _01398_ _01222_ _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05001_ _00001_ _00698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_113_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09740_ _01973_ _01985_ _04854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08479__I _03739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06952_ _00768_ _02567_ _02568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
.ends

