VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tholin_avalonsemi_tbb1143
  CLASS BLOCK ;
  FOREIGN tholin_avalonsemi_tbb1143 ;
  ORIGIN 0.000 0.000 ;
  SIZE 230.000 BY 230.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 13.440 230.000 14.000 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 47.040 230.000 47.600 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 63.840 230.000 64.400 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 80.640 230.000 81.200 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 97.440 230.000 98.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 114.240 230.000 114.800 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 131.040 230.000 131.600 ;
    END
  END io_in[5]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 147.840 230.000 148.400 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 164.640 230.000 165.200 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 181.440 230.000 182.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 198.240 230.000 198.800 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 215.040 230.000 215.600 ;
    END
  END io_out[4]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 30.240 230.000 30.800 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 211.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 211.980 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 211.980 ;
    END
  END vss
  OBS
      LAYER Pwell ;
        RECT 6.290 209.920 223.310 212.110 ;
      LAYER Nwell ;
        RECT 6.290 205.725 223.310 209.920 ;
        RECT 6.290 205.600 162.785 205.725 ;
      LAYER Pwell ;
        RECT 6.290 202.080 223.310 205.600 ;
      LAYER Nwell ;
        RECT 6.290 201.955 138.145 202.080 ;
        RECT 6.290 197.885 223.310 201.955 ;
        RECT 6.290 197.760 149.905 197.885 ;
      LAYER Pwell ;
        RECT 6.290 194.240 223.310 197.760 ;
      LAYER Nwell ;
        RECT 6.290 194.115 139.825 194.240 ;
        RECT 6.290 190.045 223.310 194.115 ;
        RECT 6.290 189.920 168.990 190.045 ;
      LAYER Pwell ;
        RECT 6.290 186.400 223.310 189.920 ;
      LAYER Nwell ;
        RECT 6.290 182.215 223.310 186.400 ;
        RECT 6.290 182.205 86.320 182.215 ;
        RECT 6.290 182.080 45.960 182.205 ;
      LAYER Pwell ;
        RECT 6.290 178.560 223.310 182.080 ;
      LAYER Nwell ;
        RECT 6.290 178.435 105.105 178.560 ;
        RECT 6.290 174.365 223.310 178.435 ;
        RECT 6.290 174.240 46.865 174.365 ;
      LAYER Pwell ;
        RECT 6.290 170.720 223.310 174.240 ;
      LAYER Nwell ;
        RECT 6.290 170.595 71.295 170.720 ;
        RECT 6.290 170.585 95.840 170.595 ;
        RECT 6.290 166.525 223.310 170.585 ;
        RECT 6.290 166.400 42.385 166.525 ;
      LAYER Pwell ;
        RECT 6.290 162.880 223.310 166.400 ;
      LAYER Nwell ;
        RECT 6.290 162.755 39.800 162.880 ;
        RECT 6.290 162.745 63.920 162.755 ;
        RECT 6.290 158.695 223.310 162.745 ;
        RECT 6.290 158.685 125.520 158.695 ;
        RECT 6.290 158.560 40.145 158.685 ;
      LAYER Pwell ;
        RECT 6.290 155.040 223.310 158.560 ;
      LAYER Nwell ;
        RECT 6.290 154.905 63.360 155.040 ;
        RECT 6.290 150.855 223.310 154.905 ;
        RECT 6.290 150.845 126.080 150.855 ;
        RECT 6.290 150.730 77.285 150.845 ;
        RECT 6.290 150.720 70.720 150.730 ;
      LAYER Pwell ;
        RECT 6.290 147.200 223.310 150.720 ;
      LAYER Nwell ;
        RECT 6.290 147.075 39.800 147.200 ;
        RECT 6.290 143.015 223.310 147.075 ;
        RECT 6.290 143.005 134.480 143.015 ;
        RECT 6.290 142.880 41.825 143.005 ;
      LAYER Pwell ;
        RECT 6.290 139.360 223.310 142.880 ;
      LAYER Nwell ;
        RECT 6.290 139.235 66.960 139.360 ;
        RECT 6.290 135.175 223.310 139.235 ;
        RECT 6.290 135.165 130.000 135.175 ;
        RECT 6.290 135.050 89.605 135.165 ;
        RECT 6.290 135.040 83.040 135.050 ;
      LAYER Pwell ;
        RECT 6.290 131.520 223.310 135.040 ;
      LAYER Nwell ;
        RECT 6.290 131.510 52.800 131.520 ;
        RECT 6.290 131.395 59.365 131.510 ;
        RECT 6.290 127.325 223.310 131.395 ;
        RECT 6.290 127.200 48.480 127.325 ;
      LAYER Pwell ;
        RECT 6.290 123.680 223.310 127.200 ;
      LAYER Nwell ;
        RECT 6.290 123.555 53.520 123.680 ;
        RECT 6.290 123.545 100.880 123.555 ;
        RECT 6.290 119.485 223.310 123.545 ;
        RECT 6.290 119.360 78.160 119.485 ;
      LAYER Pwell ;
        RECT 6.290 115.840 223.310 119.360 ;
      LAYER Nwell ;
        RECT 6.290 115.830 56.160 115.840 ;
        RECT 6.290 115.715 62.725 115.830 ;
        RECT 6.290 111.645 223.310 115.715 ;
        RECT 6.290 111.530 43.125 111.645 ;
        RECT 6.290 111.520 36.560 111.530 ;
      LAYER Pwell ;
        RECT 6.290 108.000 223.310 111.520 ;
      LAYER Nwell ;
        RECT 6.290 107.990 21.440 108.000 ;
        RECT 6.290 107.875 28.005 107.990 ;
        RECT 6.290 103.805 223.310 107.875 ;
        RECT 6.290 103.680 44.000 103.805 ;
      LAYER Pwell ;
        RECT 6.290 100.160 223.310 103.680 ;
      LAYER Nwell ;
        RECT 6.290 100.150 12.480 100.160 ;
        RECT 6.290 100.035 19.045 100.150 ;
        RECT 6.290 100.025 189.360 100.035 ;
        RECT 6.290 95.965 223.310 100.025 ;
        RECT 6.290 95.840 80.120 95.965 ;
      LAYER Pwell ;
        RECT 6.290 92.320 223.310 95.840 ;
      LAYER Nwell ;
        RECT 6.290 92.195 9.840 92.320 ;
        RECT 6.290 88.125 223.310 92.195 ;
        RECT 6.290 88.000 30.560 88.125 ;
      LAYER Pwell ;
        RECT 6.290 84.480 223.310 88.000 ;
      LAYER Nwell ;
        RECT 6.290 84.345 32.845 84.480 ;
        RECT 6.290 80.285 223.310 84.345 ;
        RECT 6.290 80.160 127.140 80.285 ;
      LAYER Pwell ;
        RECT 6.290 76.640 223.310 80.160 ;
      LAYER Nwell ;
        RECT 6.290 76.515 51.905 76.640 ;
        RECT 6.290 72.445 223.310 76.515 ;
        RECT 6.290 72.320 49.105 72.445 ;
      LAYER Pwell ;
        RECT 6.290 68.800 223.310 72.320 ;
      LAYER Nwell ;
        RECT 6.290 68.675 58.625 68.800 ;
        RECT 6.290 68.665 189.360 68.675 ;
        RECT 6.290 64.605 223.310 68.665 ;
        RECT 6.290 64.480 78.785 64.605 ;
      LAYER Pwell ;
        RECT 6.290 60.960 223.310 64.480 ;
      LAYER Nwell ;
        RECT 6.290 60.835 73.745 60.960 ;
        RECT 6.290 56.765 223.310 60.835 ;
        RECT 6.290 56.640 90.200 56.765 ;
      LAYER Pwell ;
        RECT 6.290 53.120 223.310 56.640 ;
      LAYER Nwell ;
        RECT 6.290 52.995 101.400 53.120 ;
        RECT 6.290 48.925 223.310 52.995 ;
        RECT 6.290 48.800 50.785 48.925 ;
      LAYER Pwell ;
        RECT 6.290 45.280 223.310 48.800 ;
      LAYER Nwell ;
        RECT 6.290 45.155 57.160 45.280 ;
        RECT 6.290 41.085 223.310 45.155 ;
        RECT 6.290 40.960 83.365 41.085 ;
      LAYER Pwell ;
        RECT 6.290 37.440 223.310 40.960 ;
      LAYER Nwell ;
        RECT 6.290 37.430 55.600 37.440 ;
        RECT 6.290 37.315 62.165 37.430 ;
        RECT 6.290 33.255 223.310 37.315 ;
        RECT 6.290 33.120 52.720 33.255 ;
      LAYER Pwell ;
        RECT 6.290 29.600 223.310 33.120 ;
      LAYER Nwell ;
        RECT 6.290 29.590 69.040 29.600 ;
        RECT 6.290 29.475 75.605 29.590 ;
        RECT 6.290 25.405 223.310 29.475 ;
        RECT 6.290 25.280 59.790 25.405 ;
      LAYER Pwell ;
        RECT 6.290 21.760 223.310 25.280 ;
      LAYER Nwell ;
        RECT 6.290 21.750 62.320 21.760 ;
        RECT 6.290 21.635 68.885 21.750 ;
        RECT 6.290 17.565 223.310 21.635 ;
        RECT 6.290 17.440 72.950 17.565 ;
      LAYER Pwell ;
        RECT 6.290 15.250 223.310 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 222.880 211.980 ;
      LAYER Metal2 ;
        RECT 7.980 13.530 223.300 215.510 ;
      LAYER Metal3 ;
        RECT 10.170 214.740 225.700 215.460 ;
        RECT 10.170 199.100 226.660 214.740 ;
        RECT 10.170 197.940 225.700 199.100 ;
        RECT 10.170 182.300 226.660 197.940 ;
        RECT 10.170 181.140 225.700 182.300 ;
        RECT 10.170 165.500 226.660 181.140 ;
        RECT 10.170 164.340 225.700 165.500 ;
        RECT 10.170 148.700 226.660 164.340 ;
        RECT 10.170 147.540 225.700 148.700 ;
        RECT 10.170 131.900 226.660 147.540 ;
        RECT 10.170 130.740 225.700 131.900 ;
        RECT 10.170 115.100 226.660 130.740 ;
        RECT 10.170 113.940 225.700 115.100 ;
        RECT 10.170 98.300 226.660 113.940 ;
        RECT 10.170 97.140 225.700 98.300 ;
        RECT 10.170 81.500 226.660 97.140 ;
        RECT 10.170 80.340 225.700 81.500 ;
        RECT 10.170 64.700 226.660 80.340 ;
        RECT 10.170 63.540 225.700 64.700 ;
        RECT 10.170 47.900 226.660 63.540 ;
        RECT 10.170 46.740 225.700 47.900 ;
        RECT 10.170 31.100 226.660 46.740 ;
        RECT 10.170 29.940 225.700 31.100 ;
        RECT 10.170 14.300 226.660 29.940 ;
        RECT 10.170 13.580 225.700 14.300 ;
      LAYER Metal4 ;
        RECT 94.220 30.330 98.740 210.470 ;
        RECT 100.940 30.330 175.540 210.470 ;
        RECT 177.740 30.330 181.860 210.470 ;
  END
END tholin_avalonsemi_tbb1143
END LIBRARY

