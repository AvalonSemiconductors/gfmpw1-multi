VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO diceroll
  CLASS BLOCK ;
  FOREIGN diceroll ;
  ORIGIN 0.000 0.000 ;
  SIZE 230.000 BY 230.000 ;
  PIN io_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 226.000 47.600 230.000 ;
    END
  END io_in
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 226.000 66.640 230.000 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 85.120 226.000 85.680 230.000 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 226.000 104.720 230.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 123.200 226.000 123.760 230.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 142.240 226.000 142.800 230.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 226.000 161.840 230.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 180.320 226.000 180.880 230.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 199.360 226.000 199.920 230.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 226.000 218.960 230.000 ;
    END
  END io_out[8]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 28.000 226.000 28.560 230.000 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 211.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 211.980 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 211.980 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 8.960 226.000 9.520 230.000 ;
    END
  END wb_clk_i
  OBS
      LAYER Pwell ;
        RECT 6.290 209.920 223.310 212.110 ;
      LAYER Nwell ;
        RECT 6.290 205.600 223.310 209.920 ;
      LAYER Pwell ;
        RECT 6.290 202.080 223.310 205.600 ;
      LAYER Nwell ;
        RECT 6.290 201.955 18.865 202.080 ;
        RECT 6.290 197.885 223.310 201.955 ;
        RECT 6.290 197.760 91.105 197.885 ;
      LAYER Pwell ;
        RECT 6.290 194.240 223.310 197.760 ;
      LAYER Nwell ;
        RECT 6.290 194.115 13.265 194.240 ;
        RECT 6.290 190.045 223.310 194.115 ;
        RECT 6.290 189.920 51.500 190.045 ;
      LAYER Pwell ;
        RECT 6.290 186.400 223.310 189.920 ;
      LAYER Nwell ;
        RECT 6.290 186.275 104.545 186.400 ;
        RECT 6.290 182.080 223.310 186.275 ;
      LAYER Pwell ;
        RECT 6.290 178.560 223.310 182.080 ;
      LAYER Nwell ;
        RECT 6.290 178.435 13.265 178.560 ;
        RECT 6.290 174.365 223.310 178.435 ;
        RECT 6.290 174.240 154.945 174.365 ;
      LAYER Pwell ;
        RECT 6.290 170.720 223.310 174.240 ;
      LAYER Nwell ;
        RECT 6.290 170.595 25.025 170.720 ;
        RECT 6.290 166.400 223.310 170.595 ;
      LAYER Pwell ;
        RECT 6.290 162.880 223.310 166.400 ;
      LAYER Nwell ;
        RECT 6.290 162.755 103.985 162.880 ;
        RECT 6.290 158.685 223.310 162.755 ;
        RECT 6.290 158.560 14.945 158.685 ;
      LAYER Pwell ;
        RECT 6.290 155.040 223.310 158.560 ;
      LAYER Nwell ;
        RECT 6.290 154.915 34.545 155.040 ;
        RECT 6.290 150.845 223.310 154.915 ;
        RECT 6.290 150.720 57.160 150.845 ;
      LAYER Pwell ;
        RECT 6.290 147.200 223.310 150.720 ;
      LAYER Nwell ;
        RECT 6.290 147.075 13.265 147.200 ;
        RECT 6.290 142.880 223.310 147.075 ;
      LAYER Pwell ;
        RECT 6.290 139.360 223.310 142.880 ;
      LAYER Nwell ;
        RECT 6.290 139.235 108.120 139.360 ;
        RECT 6.290 135.165 223.310 139.235 ;
        RECT 6.290 135.040 209.265 135.165 ;
      LAYER Pwell ;
        RECT 6.290 131.520 223.310 135.040 ;
      LAYER Nwell ;
        RECT 6.290 127.325 223.310 131.520 ;
        RECT 6.290 127.200 197.830 127.325 ;
      LAYER Pwell ;
        RECT 6.290 123.680 223.310 127.200 ;
      LAYER Nwell ;
        RECT 6.290 123.555 181.265 123.680 ;
        RECT 6.290 119.485 223.310 123.555 ;
        RECT 6.290 119.360 91.755 119.485 ;
      LAYER Pwell ;
        RECT 6.290 115.840 223.310 119.360 ;
      LAYER Nwell ;
        RECT 6.290 115.715 65.910 115.840 ;
        RECT 6.290 111.645 223.310 115.715 ;
        RECT 6.290 111.520 13.265 111.645 ;
      LAYER Pwell ;
        RECT 6.290 108.000 223.310 111.520 ;
      LAYER Nwell ;
        RECT 6.290 107.875 70.150 108.000 ;
        RECT 6.290 103.680 223.310 107.875 ;
      LAYER Pwell ;
        RECT 6.290 100.160 223.310 103.680 ;
      LAYER Nwell ;
        RECT 6.290 100.035 16.065 100.160 ;
        RECT 6.290 95.965 223.310 100.035 ;
        RECT 6.290 95.840 118.545 95.965 ;
      LAYER Pwell ;
        RECT 6.290 92.320 223.310 95.840 ;
      LAYER Nwell ;
        RECT 6.290 92.195 103.080 92.320 ;
        RECT 6.290 88.125 223.310 92.195 ;
        RECT 6.290 88.000 208.705 88.125 ;
      LAYER Pwell ;
        RECT 6.290 84.480 223.310 88.000 ;
      LAYER Nwell ;
        RECT 6.290 84.355 22.225 84.480 ;
        RECT 6.290 80.285 223.310 84.355 ;
        RECT 6.290 80.160 13.265 80.285 ;
      LAYER Pwell ;
        RECT 6.290 76.640 223.310 80.160 ;
      LAYER Nwell ;
        RECT 6.290 76.515 138.920 76.640 ;
        RECT 6.290 72.320 223.310 76.515 ;
      LAYER Pwell ;
        RECT 6.290 68.800 223.310 72.320 ;
      LAYER Nwell ;
        RECT 6.290 68.675 209.265 68.800 ;
        RECT 6.290 64.480 223.310 68.675 ;
      LAYER Pwell ;
        RECT 6.290 60.960 223.310 64.480 ;
      LAYER Nwell ;
        RECT 6.290 60.835 21.105 60.960 ;
        RECT 6.290 56.765 223.310 60.835 ;
        RECT 6.290 56.640 13.265 56.765 ;
      LAYER Pwell ;
        RECT 6.290 53.120 223.310 56.640 ;
      LAYER Nwell ;
        RECT 6.290 52.995 152.145 53.120 ;
        RECT 6.290 48.925 223.310 52.995 ;
        RECT 6.290 48.800 132.545 48.925 ;
      LAYER Pwell ;
        RECT 6.290 45.280 223.310 48.800 ;
      LAYER Nwell ;
        RECT 6.290 45.155 179.025 45.280 ;
        RECT 6.290 41.085 223.310 45.155 ;
        RECT 6.290 40.960 37.560 41.085 ;
      LAYER Pwell ;
        RECT 6.290 37.440 223.310 40.960 ;
      LAYER Nwell ;
        RECT 6.290 33.245 223.310 37.440 ;
        RECT 6.290 33.120 57.720 33.245 ;
      LAYER Pwell ;
        RECT 6.290 29.600 223.310 33.120 ;
      LAYER Nwell ;
        RECT 6.290 29.475 130.305 29.600 ;
        RECT 6.290 25.405 223.310 29.475 ;
        RECT 6.290 25.280 82.705 25.405 ;
      LAYER Pwell ;
        RECT 6.290 21.760 223.310 25.280 ;
      LAYER Nwell ;
        RECT 6.290 21.635 71.505 21.760 ;
        RECT 6.290 17.440 223.310 21.635 ;
      LAYER Pwell ;
        RECT 6.290 15.250 223.310 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 222.880 211.980 ;
      LAYER Metal2 ;
        RECT 9.820 225.700 27.700 226.660 ;
        RECT 28.860 225.700 46.740 226.660 ;
        RECT 47.900 225.700 65.780 226.660 ;
        RECT 66.940 225.700 84.820 226.660 ;
        RECT 85.980 225.700 103.860 226.660 ;
        RECT 105.020 225.700 122.900 226.660 ;
        RECT 124.060 225.700 141.940 226.660 ;
        RECT 143.100 225.700 160.980 226.660 ;
        RECT 162.140 225.700 180.020 226.660 ;
        RECT 181.180 225.700 199.060 226.660 ;
        RECT 200.220 225.700 218.100 226.660 ;
        RECT 219.260 225.700 220.500 226.660 ;
        RECT 9.100 15.490 220.500 225.700 ;
      LAYER Metal3 ;
        RECT 9.610 15.540 220.550 211.820 ;
      LAYER Metal4 ;
        RECT 76.860 44.890 79.380 54.230 ;
  END
END diceroll
END LIBRARY

