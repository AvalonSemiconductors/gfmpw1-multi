VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO hellorld
  CLASS BLOCK ;
  FOREIGN hellorld ;
  ORIGIN 0.000 0.000 ;
  SIZE 130.000 BY 130.000 ;
  PIN custom_settings[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 126.000 8.960 130.000 9.520 ;
    END
  END custom_settings[0]
  PIN custom_settings[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 126.000 109.760 130.000 110.320 ;
    END
  END custom_settings[10]
  PIN custom_settings[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 126.000 119.840 130.000 120.400 ;
    END
  END custom_settings[11]
  PIN custom_settings[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 126.000 19.040 130.000 19.600 ;
    END
  END custom_settings[1]
  PIN custom_settings[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 126.000 29.120 130.000 29.680 ;
    END
  END custom_settings[2]
  PIN custom_settings[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 126.000 39.200 130.000 39.760 ;
    END
  END custom_settings[3]
  PIN custom_settings[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 126.000 49.280 130.000 49.840 ;
    END
  END custom_settings[4]
  PIN custom_settings[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 126.000 59.360 130.000 59.920 ;
    END
  END custom_settings[5]
  PIN custom_settings[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 126.000 69.440 130.000 70.000 ;
    END
  END custom_settings[6]
  PIN custom_settings[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 126.000 79.520 130.000 80.080 ;
    END
  END custom_settings[7]
  PIN custom_settings[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 126.000 89.600 130.000 90.160 ;
    END
  END custom_settings[8]
  PIN custom_settings[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 126.000 99.680 130.000 100.240 ;
    END
  END custom_settings[9]
  PIN io_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 106.400 126.000 106.960 130.000 ;
    END
  END io_out
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 126.000 64.400 130.000 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 20.480 15.380 22.080 113.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 49.600 15.380 51.200 113.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 78.720 15.380 80.320 113.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 107.840 15.380 109.440 113.980 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 35.040 15.380 36.640 113.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 64.160 15.380 65.760 113.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 93.280 15.380 94.880 113.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.400 15.380 124.000 113.980 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.352000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 21.280 126.000 21.840 130.000 ;
    END
  END wb_clk_i
  OBS
      LAYER Nwell ;
        RECT 6.290 111.530 123.630 114.110 ;
      LAYER Pwell ;
        RECT 6.290 107.990 123.630 111.530 ;
      LAYER Nwell ;
        RECT 6.290 103.690 123.630 107.990 ;
      LAYER Pwell ;
        RECT 6.290 100.150 123.630 103.690 ;
      LAYER Nwell ;
        RECT 6.290 95.850 123.630 100.150 ;
      LAYER Pwell ;
        RECT 6.290 92.310 123.630 95.850 ;
      LAYER Nwell ;
        RECT 6.290 88.010 123.630 92.310 ;
      LAYER Pwell ;
        RECT 6.290 84.470 123.630 88.010 ;
      LAYER Nwell ;
        RECT 6.290 80.170 123.630 84.470 ;
      LAYER Pwell ;
        RECT 6.290 76.630 123.630 80.170 ;
      LAYER Nwell ;
        RECT 6.290 72.330 123.630 76.630 ;
      LAYER Pwell ;
        RECT 6.290 68.790 123.630 72.330 ;
      LAYER Nwell ;
        RECT 6.290 64.490 123.630 68.790 ;
      LAYER Pwell ;
        RECT 6.290 60.950 123.630 64.490 ;
      LAYER Nwell ;
        RECT 6.290 56.650 123.630 60.950 ;
      LAYER Pwell ;
        RECT 6.290 53.110 123.630 56.650 ;
      LAYER Nwell ;
        RECT 6.290 48.810 123.630 53.110 ;
      LAYER Pwell ;
        RECT 6.290 45.270 123.630 48.810 ;
      LAYER Nwell ;
        RECT 6.290 40.970 123.630 45.270 ;
      LAYER Pwell ;
        RECT 6.290 37.430 123.630 40.970 ;
      LAYER Nwell ;
        RECT 6.290 33.130 123.630 37.430 ;
      LAYER Pwell ;
        RECT 6.290 29.590 123.630 33.130 ;
      LAYER Nwell ;
        RECT 6.290 25.290 123.630 29.590 ;
      LAYER Pwell ;
        RECT 6.290 21.750 123.630 25.290 ;
      LAYER Nwell ;
        RECT 6.290 17.450 123.630 21.750 ;
      LAYER Pwell ;
        RECT 6.290 15.250 123.630 17.450 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 124.000 114.650 ;
      LAYER Metal2 ;
        RECT 7.980 125.700 20.980 126.000 ;
        RECT 22.140 125.700 63.540 126.000 ;
        RECT 64.700 125.700 106.100 126.000 ;
        RECT 107.260 125.700 125.300 126.000 ;
        RECT 7.980 9.050 125.300 125.700 ;
      LAYER Metal3 ;
        RECT 7.930 119.540 125.700 120.260 ;
        RECT 7.930 110.620 126.000 119.540 ;
        RECT 7.930 109.460 125.700 110.620 ;
        RECT 7.930 100.540 126.000 109.460 ;
        RECT 7.930 99.380 125.700 100.540 ;
        RECT 7.930 90.460 126.000 99.380 ;
        RECT 7.930 89.300 125.700 90.460 ;
        RECT 7.930 80.380 126.000 89.300 ;
        RECT 7.930 79.220 125.700 80.380 ;
        RECT 7.930 70.300 126.000 79.220 ;
        RECT 7.930 69.140 125.700 70.300 ;
        RECT 7.930 60.220 126.000 69.140 ;
        RECT 7.930 59.060 125.700 60.220 ;
        RECT 7.930 50.140 126.000 59.060 ;
        RECT 7.930 48.980 125.700 50.140 ;
        RECT 7.930 40.060 126.000 48.980 ;
        RECT 7.930 38.900 125.700 40.060 ;
        RECT 7.930 29.980 126.000 38.900 ;
        RECT 7.930 28.820 125.700 29.980 ;
        RECT 7.930 19.900 126.000 28.820 ;
        RECT 7.930 18.740 125.700 19.900 ;
        RECT 7.930 9.820 126.000 18.740 ;
        RECT 7.930 9.100 125.700 9.820 ;
      LAYER Metal4 ;
        RECT 33.740 52.170 34.740 101.830 ;
        RECT 36.940 52.170 49.300 101.830 ;
        RECT 51.500 52.170 63.860 101.830 ;
        RECT 66.060 52.170 78.420 101.830 ;
        RECT 80.620 52.170 92.980 101.830 ;
        RECT 95.180 52.170 107.540 101.830 ;
        RECT 109.740 52.170 113.540 101.830 ;
  END
END hellorld
END LIBRARY

